--------------------------------------------------------------------------------
-- Company:        ENSIMAG
-- Engineer:       Hans Julien, Perraud Frédéric
-- 
-- Create Date:    08:11:44 03/12/2015 
-- Design Name: 
-- Module Name:    Rom with a complete image
-- Project Name:   pedestre detection HLS
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
--------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;

entity MEM_ROM is
  port ( clk :     in std_logic;
         address : in std_logic_vector(16 downto 0);
         data :    out std_logic_vector(7 downto 0) );
end entity MEM_ROM;

architecture behavioral of MEM_ROM is
  type mem is array ( 0 to 320*240 - 1) of std_logic_vector(7 downto 0);
  constant my_Rom : mem := (

0	 => std_logic_vector(to_unsigned(10,8) ,
1	 => std_logic_vector(to_unsigned(112,8) ,
2	 => std_logic_vector(to_unsigned(118,8) ,
3	 => std_logic_vector(to_unsigned(116,8) ,
4	 => std_logic_vector(to_unsigned(114,8) ,
5	 => std_logic_vector(to_unsigned(108,8) ,
6	 => std_logic_vector(to_unsigned(109,8) ,
7	 => std_logic_vector(to_unsigned(108,8) ,
8	 => std_logic_vector(to_unsigned(107,8) ,
9	 => std_logic_vector(to_unsigned(105,8) ,
10	 => std_logic_vector(to_unsigned(107,8) ,
11	 => std_logic_vector(to_unsigned(104,8) ,
12	 => std_logic_vector(to_unsigned(104,8) ,
13	 => std_logic_vector(to_unsigned(111,8) ,
14	 => std_logic_vector(to_unsigned(107,8) ,
15	 => std_logic_vector(to_unsigned(107,8) ,
16	 => std_logic_vector(to_unsigned(104,8) ,
17	 => std_logic_vector(to_unsigned(99,8) ,
18	 => std_logic_vector(to_unsigned(101,8) ,
19	 => std_logic_vector(to_unsigned(96,8) ,
20	 => std_logic_vector(to_unsigned(93,8) ,
21	 => std_logic_vector(to_unsigned(90,8) ,
22	 => std_logic_vector(to_unsigned(95,8) ,
23	 => std_logic_vector(to_unsigned(96,8) ,
24	 => std_logic_vector(to_unsigned(93,8) ,
25	 => std_logic_vector(to_unsigned(104,8) ,
26	 => std_logic_vector(to_unsigned(105,8) ,
27	 => std_logic_vector(to_unsigned(105,8) ,
28	 => std_logic_vector(to_unsigned(108,8) ,
29	 => std_logic_vector(to_unsigned(103,8) ,
30	 => std_logic_vector(to_unsigned(108,8) ,
31	 => std_logic_vector(to_unsigned(111,8) ,
32	 => std_logic_vector(to_unsigned(109,8) ,
33	 => std_logic_vector(to_unsigned(109,8) ,
34	 => std_logic_vector(to_unsigned(114,8) ,
35	 => std_logic_vector(to_unsigned(111,8) ,
36	 => std_logic_vector(to_unsigned(109,8) ,
37	 => std_logic_vector(to_unsigned(114,8) ,
38	 => std_logic_vector(to_unsigned(115,8) ,
39	 => std_logic_vector(to_unsigned(115,8) ,
40	 => std_logic_vector(to_unsigned(118,8) ,
41	 => std_logic_vector(to_unsigned(116,8) ,
42	 => std_logic_vector(to_unsigned(119,8) ,
43	 => std_logic_vector(to_unsigned(116,8) ,
44	 => std_logic_vector(to_unsigned(114,8) ,
45	 => std_logic_vector(to_unsigned(115,8) ,
46	 => std_logic_vector(to_unsigned(116,8) ,
47	 => std_logic_vector(to_unsigned(115,8) ,
48	 => std_logic_vector(to_unsigned(119,8) ,
49	 => std_logic_vector(to_unsigned(118,8) ,
50	 => std_logic_vector(to_unsigned(116,8) ,
51	 => std_logic_vector(to_unsigned(116,8) ,
52	 => std_logic_vector(to_unsigned(115,8) ,
53	 => std_logic_vector(to_unsigned(111,8) ,
54	 => std_logic_vector(to_unsigned(115,8) ,
55	 => std_logic_vector(to_unsigned(118,8) ,
56	 => std_logic_vector(to_unsigned(115,8) ,
57	 => std_logic_vector(to_unsigned(116,8) ,
58	 => std_logic_vector(to_unsigned(118,8) ,
59	 => std_logic_vector(to_unsigned(112,8) ,
60	 => std_logic_vector(to_unsigned(104,8) ,
61	 => std_logic_vector(to_unsigned(104,8) ,
62	 => std_logic_vector(to_unsigned(111,8) ,
63	 => std_logic_vector(to_unsigned(118,8) ,
64	 => std_logic_vector(to_unsigned(116,8) ,
65	 => std_logic_vector(to_unsigned(114,8) ,
66	 => std_logic_vector(to_unsigned(116,8) ,
67	 => std_logic_vector(to_unsigned(119,8) ,
68	 => std_logic_vector(to_unsigned(118,8) ,
69	 => std_logic_vector(to_unsigned(115,8) ,
70	 => std_logic_vector(to_unsigned(114,8) ,
71	 => std_logic_vector(to_unsigned(112,8) ,
72	 => std_logic_vector(to_unsigned(115,8) ,
73	 => std_logic_vector(to_unsigned(118,8) ,
74	 => std_logic_vector(to_unsigned(114,8) ,
75	 => std_logic_vector(to_unsigned(112,8) ,
76	 => std_logic_vector(to_unsigned(109,8) ,
77	 => std_logic_vector(to_unsigned(115,8) ,
78	 => std_logic_vector(to_unsigned(114,8) ,
79	 => std_logic_vector(to_unsigned(107,8) ,
80	 => std_logic_vector(to_unsigned(108,8) ,
81	 => std_logic_vector(to_unsigned(112,8) ,
82	 => std_logic_vector(to_unsigned(107,8) ,
83	 => std_logic_vector(to_unsigned(115,8) ,
84	 => std_logic_vector(to_unsigned(115,8) ,
85	 => std_logic_vector(to_unsigned(114,8) ,
86	 => std_logic_vector(to_unsigned(115,8) ,
87	 => std_logic_vector(to_unsigned(109,8) ,
88	 => std_logic_vector(to_unsigned(112,8) ,
89	 => std_logic_vector(to_unsigned(109,8) ,
90	 => std_logic_vector(to_unsigned(109,8) ,
91	 => std_logic_vector(to_unsigned(109,8) ,
92	 => std_logic_vector(to_unsigned(109,8) ,
93	 => std_logic_vector(to_unsigned(108,8) ,
94	 => std_logic_vector(to_unsigned(105,8) ,
95	 => std_logic_vector(to_unsigned(100,8) ,
96	 => std_logic_vector(to_unsigned(100,8) ,
97	 => std_logic_vector(to_unsigned(107,8) ,
98	 => std_logic_vector(to_unsigned(103,8) ,
99	 => std_logic_vector(to_unsigned(105,8) ,
100	 => std_logic_vector(to_unsigned(104,8) ,
101	 => std_logic_vector(to_unsigned(107,8) ,
102	 => std_logic_vector(to_unsigned(111,8) ,
103	 => std_logic_vector(to_unsigned(107,8) ,
104	 => std_logic_vector(to_unsigned(105,8) ,
105	 => std_logic_vector(to_unsigned(109,8) ,
106	 => std_logic_vector(to_unsigned(107,8) ,
107	 => std_logic_vector(to_unsigned(103,8) ,
108	 => std_logic_vector(to_unsigned(111,8) ,
109	 => std_logic_vector(to_unsigned(115,8) ,
110	 => std_logic_vector(to_unsigned(112,8) ,
111	 => std_logic_vector(to_unsigned(107,8) ,
112	 => std_logic_vector(to_unsigned(108,8) ,
113	 => std_logic_vector(to_unsigned(114,8) ,
114	 => std_logic_vector(to_unsigned(114,8) ,
115	 => std_logic_vector(to_unsigned(115,8) ,
116	 => std_logic_vector(to_unsigned(111,8) ,
117	 => std_logic_vector(to_unsigned(104,8) ,
118	 => std_logic_vector(to_unsigned(103,8) ,
119	 => std_logic_vector(to_unsigned(107,8) ,
120	 => std_logic_vector(to_unsigned(105,8) ,
121	 => std_logic_vector(to_unsigned(101,8) ,
122	 => std_logic_vector(to_unsigned(99,8) ,
123	 => std_logic_vector(to_unsigned(99,8) ,
124	 => std_logic_vector(to_unsigned(100,8) ,
125	 => std_logic_vector(to_unsigned(104,8) ,
126	 => std_logic_vector(to_unsigned(103,8) ,
127	 => std_logic_vector(to_unsigned(101,8) ,
128	 => std_logic_vector(to_unsigned(103,8) ,
129	 => std_logic_vector(to_unsigned(103,8) ,
130	 => std_logic_vector(to_unsigned(101,8) ,
131	 => std_logic_vector(to_unsigned(103,8) ,
132	 => std_logic_vector(to_unsigned(105,8) ,
133	 => std_logic_vector(to_unsigned(103,8) ,
134	 => std_logic_vector(to_unsigned(101,8) ,
135	 => std_logic_vector(to_unsigned(99,8) ,
136	 => std_logic_vector(to_unsigned(97,8) ,
137	 => std_logic_vector(to_unsigned(99,8) ,
138	 => std_logic_vector(to_unsigned(100,8) ,
139	 => std_logic_vector(to_unsigned(99,8) ,
140	 => std_logic_vector(to_unsigned(104,8) ,
141	 => std_logic_vector(to_unsigned(104,8) ,
142	 => std_logic_vector(to_unsigned(104,8) ,
143	 => std_logic_vector(to_unsigned(101,8) ,
144	 => std_logic_vector(to_unsigned(101,8) ,
145	 => std_logic_vector(to_unsigned(101,8) ,
146	 => std_logic_vector(to_unsigned(101,8) ,
147	 => std_logic_vector(to_unsigned(101,8) ,
148	 => std_logic_vector(to_unsigned(104,8) ,
149	 => std_logic_vector(to_unsigned(104,8) ,
150	 => std_logic_vector(to_unsigned(108,8) ,
151	 => std_logic_vector(to_unsigned(100,8) ,
152	 => std_logic_vector(to_unsigned(97,8) ,
153	 => std_logic_vector(to_unsigned(97,8) ,
154	 => std_logic_vector(to_unsigned(93,8) ,
155	 => std_logic_vector(to_unsigned(97,8) ,
156	 => std_logic_vector(to_unsigned(90,8) ,
157	 => std_logic_vector(to_unsigned(90,8) ,
158	 => std_logic_vector(to_unsigned(92,8) ,
159	 => std_logic_vector(to_unsigned(93,8) ,
160	 => std_logic_vector(to_unsigned(91,8) ,
161	 => std_logic_vector(to_unsigned(92,8) ,
162	 => std_logic_vector(to_unsigned(95,8) ,
163	 => std_logic_vector(to_unsigned(92,8) ,
164	 => std_logic_vector(to_unsigned(92,8) ,
165	 => std_logic_vector(to_unsigned(93,8) ,
166	 => std_logic_vector(to_unsigned(92,8) ,
167	 => std_logic_vector(to_unsigned(90,8) ,
168	 => std_logic_vector(to_unsigned(90,8) ,
169	 => std_logic_vector(to_unsigned(96,8) ,
170	 => std_logic_vector(to_unsigned(95,8) ,
171	 => std_logic_vector(to_unsigned(95,8) ,
172	 => std_logic_vector(to_unsigned(95,8) ,
173	 => std_logic_vector(to_unsigned(90,8) ,
174	 => std_logic_vector(to_unsigned(91,8) ,
175	 => std_logic_vector(to_unsigned(92,8) ,
176	 => std_logic_vector(to_unsigned(85,8) ,
177	 => std_logic_vector(to_unsigned(82,8) ,
178	 => std_logic_vector(to_unsigned(84,8) ,
179	 => std_logic_vector(to_unsigned(87,8) ,
180	 => std_logic_vector(to_unsigned(91,8) ,
181	 => std_logic_vector(to_unsigned(88,8) ,
182	 => std_logic_vector(to_unsigned(86,8) ,
183	 => std_logic_vector(to_unsigned(90,8) ,
184	 => std_logic_vector(to_unsigned(92,8) ,
185	 => std_logic_vector(to_unsigned(90,8) ,
186	 => std_logic_vector(to_unsigned(90,8) ,
187	 => std_logic_vector(to_unsigned(91,8) ,
188	 => std_logic_vector(to_unsigned(90,8) ,
189	 => std_logic_vector(to_unsigned(92,8) ,
190	 => std_logic_vector(to_unsigned(92,8) ,
191	 => std_logic_vector(to_unsigned(91,8) ,
192	 => std_logic_vector(to_unsigned(88,8) ,
193	 => std_logic_vector(to_unsigned(88,8) ,
194	 => std_logic_vector(to_unsigned(88,8) ,
195	 => std_logic_vector(to_unsigned(90,8) ,
196	 => std_logic_vector(to_unsigned(87,8) ,
197	 => std_logic_vector(to_unsigned(84,8) ,
198	 => std_logic_vector(to_unsigned(90,8) ,
199	 => std_logic_vector(to_unsigned(91,8) ,
200	 => std_logic_vector(to_unsigned(88,8) ,
201	 => std_logic_vector(to_unsigned(92,8) ,
202	 => std_logic_vector(to_unsigned(96,8) ,
203	 => std_logic_vector(to_unsigned(91,8) ,
204	 => std_logic_vector(to_unsigned(92,8) ,
205	 => std_logic_vector(to_unsigned(97,8) ,
206	 => std_logic_vector(to_unsigned(99,8) ,
207	 => std_logic_vector(to_unsigned(99,8) ,
208	 => std_logic_vector(to_unsigned(99,8) ,
209	 => std_logic_vector(to_unsigned(97,8) ,
210	 => std_logic_vector(to_unsigned(99,8) ,
211	 => std_logic_vector(to_unsigned(99,8) ,
212	 => std_logic_vector(to_unsigned(95,8) ,
213	 => std_logic_vector(to_unsigned(99,8) ,
214	 => std_logic_vector(to_unsigned(100,8) ,
215	 => std_logic_vector(to_unsigned(93,8) ,
216	 => std_logic_vector(to_unsigned(96,8) ,
217	 => std_logic_vector(to_unsigned(96,8) ,
218	 => std_logic_vector(to_unsigned(91,8) ,
219	 => std_logic_vector(to_unsigned(97,8) ,
220	 => std_logic_vector(to_unsigned(95,8) ,
221	 => std_logic_vector(to_unsigned(95,8) ,
222	 => std_logic_vector(to_unsigned(93,8) ,
223	 => std_logic_vector(to_unsigned(91,8) ,
224	 => std_logic_vector(to_unsigned(90,8) ,
225	 => std_logic_vector(to_unsigned(95,8) ,
226	 => std_logic_vector(to_unsigned(95,8) ,
227	 => std_logic_vector(to_unsigned(97,8) ,
228	 => std_logic_vector(to_unsigned(101,8) ,
229	 => std_logic_vector(to_unsigned(96,8) ,
230	 => std_logic_vector(to_unsigned(99,8) ,
231	 => std_logic_vector(to_unsigned(100,8) ,
232	 => std_logic_vector(to_unsigned(103,8) ,
233	 => std_logic_vector(to_unsigned(103,8) ,
234	 => std_logic_vector(to_unsigned(101,8) ,
235	 => std_logic_vector(to_unsigned(19,8) ,
236	 => std_logic_vector(to_unsigned(0,8) ,
237	 => std_logic_vector(to_unsigned(0,8) ,
238	 => std_logic_vector(to_unsigned(10,8) ,
239	 => std_logic_vector(to_unsigned(100,8) ,
240	 => std_logic_vector(to_unsigned(95,8) ,
241	 => std_logic_vector(to_unsigned(88,8) ,
242	 => std_logic_vector(to_unsigned(88,8) ,
243	 => std_logic_vector(to_unsigned(95,8) ,
244	 => std_logic_vector(to_unsigned(99,8) ,
245	 => std_logic_vector(to_unsigned(100,8) ,
246	 => std_logic_vector(to_unsigned(105,8) ,
247	 => std_logic_vector(to_unsigned(103,8) ,
248	 => std_logic_vector(to_unsigned(108,8) ,
249	 => std_logic_vector(to_unsigned(114,8) ,
250	 => std_logic_vector(to_unsigned(115,8) ,
251	 => std_logic_vector(to_unsigned(114,8) ,
252	 => std_logic_vector(to_unsigned(107,8) ,
253	 => std_logic_vector(to_unsigned(107,8) ,
254	 => std_logic_vector(to_unsigned(112,8) ,
255	 => std_logic_vector(to_unsigned(119,8) ,
256	 => std_logic_vector(to_unsigned(118,8) ,
257	 => std_logic_vector(to_unsigned(109,8) ,
258	 => std_logic_vector(to_unsigned(111,8) ,
259	 => std_logic_vector(to_unsigned(112,8) ,
260	 => std_logic_vector(to_unsigned(114,8) ,
261	 => std_logic_vector(to_unsigned(115,8) ,
262	 => std_logic_vector(to_unsigned(114,8) ,
263	 => std_logic_vector(to_unsigned(118,8) ,
264	 => std_logic_vector(to_unsigned(116,8) ,
265	 => std_logic_vector(to_unsigned(119,8) ,
266	 => std_logic_vector(to_unsigned(118,8) ,
267	 => std_logic_vector(to_unsigned(112,8) ,
268	 => std_logic_vector(to_unsigned(115,8) ,
269	 => std_logic_vector(to_unsigned(116,8) ,
270	 => std_logic_vector(to_unsigned(118,8) ,
271	 => std_logic_vector(to_unsigned(125,8) ,
272	 => std_logic_vector(to_unsigned(125,8) ,
273	 => std_logic_vector(to_unsigned(127,8) ,
274	 => std_logic_vector(to_unsigned(131,8) ,
275	 => std_logic_vector(to_unsigned(130,8) ,
276	 => std_logic_vector(to_unsigned(134,8) ,
277	 => std_logic_vector(to_unsigned(141,8) ,
278	 => std_logic_vector(to_unsigned(138,8) ,
279	 => std_logic_vector(to_unsigned(138,8) ,
280	 => std_logic_vector(to_unsigned(138,8) ,
281	 => std_logic_vector(to_unsigned(144,8) ,
282	 => std_logic_vector(to_unsigned(147,8) ,
283	 => std_logic_vector(to_unsigned(151,8) ,
284	 => std_logic_vector(to_unsigned(149,8) ,
285	 => std_logic_vector(to_unsigned(147,8) ,
286	 => std_logic_vector(to_unsigned(147,8) ,
287	 => std_logic_vector(to_unsigned(149,8) ,
288	 => std_logic_vector(to_unsigned(152,8) ,
289	 => std_logic_vector(to_unsigned(157,8) ,
290	 => std_logic_vector(to_unsigned(157,8) ,
291	 => std_logic_vector(to_unsigned(156,8) ,
292	 => std_logic_vector(to_unsigned(156,8) ,
293	 => std_logic_vector(to_unsigned(157,8) ,
294	 => std_logic_vector(to_unsigned(157,8) ,
295	 => std_logic_vector(to_unsigned(161,8) ,
296	 => std_logic_vector(to_unsigned(161,8) ,
297	 => std_logic_vector(to_unsigned(157,8) ,
298	 => std_logic_vector(to_unsigned(159,8) ,
299	 => std_logic_vector(to_unsigned(161,8) ,
300	 => std_logic_vector(to_unsigned(161,8) ,
301	 => std_logic_vector(to_unsigned(157,8) ,
302	 => std_logic_vector(to_unsigned(156,8) ,
303	 => std_logic_vector(to_unsigned(161,8) ,
304	 => std_logic_vector(to_unsigned(161,8) ,
305	 => std_logic_vector(to_unsigned(161,8) ,
306	 => std_logic_vector(to_unsigned(164,8) ,
307	 => std_logic_vector(to_unsigned(163,8) ,
308	 => std_logic_vector(to_unsigned(163,8) ,
309	 => std_logic_vector(to_unsigned(166,8) ,
310	 => std_logic_vector(to_unsigned(164,8) ,
311	 => std_logic_vector(to_unsigned(163,8) ,
312	 => std_logic_vector(to_unsigned(161,8) ,
313	 => std_logic_vector(to_unsigned(163,8) ,
314	 => std_logic_vector(to_unsigned(163,8) ,
315	 => std_logic_vector(to_unsigned(161,8) ,
316	 => std_logic_vector(to_unsigned(161,8) ,
317	 => std_logic_vector(to_unsigned(163,8) ,
318	 => std_logic_vector(to_unsigned(166,8) ,
319	 => std_logic_vector(to_unsigned(164,8) ,
320	 => std_logic_vector(to_unsigned(161,8) ,
321	 => std_logic_vector(to_unsigned(111,8) ,
322	 => std_logic_vector(to_unsigned(107,8) ,
323	 => std_logic_vector(to_unsigned(109,8) ,
324	 => std_logic_vector(to_unsigned(114,8) ,
325	 => std_logic_vector(to_unsigned(109,8) ,
326	 => std_logic_vector(to_unsigned(107,8) ,
327	 => std_logic_vector(to_unsigned(104,8) ,
328	 => std_logic_vector(to_unsigned(105,8) ,
329	 => std_logic_vector(to_unsigned(105,8) ,
330	 => std_logic_vector(to_unsigned(105,8) ,
331	 => std_logic_vector(to_unsigned(104,8) ,
332	 => std_logic_vector(to_unsigned(105,8) ,
333	 => std_logic_vector(to_unsigned(108,8) ,
334	 => std_logic_vector(to_unsigned(99,8) ,
335	 => std_logic_vector(to_unsigned(97,8) ,
336	 => std_logic_vector(to_unsigned(93,8) ,
337	 => std_logic_vector(to_unsigned(88,8) ,
338	 => std_logic_vector(to_unsigned(95,8) ,
339	 => std_logic_vector(to_unsigned(96,8) ,
340	 => std_logic_vector(to_unsigned(92,8) ,
341	 => std_logic_vector(to_unsigned(88,8) ,
342	 => std_logic_vector(to_unsigned(91,8) ,
343	 => std_logic_vector(to_unsigned(92,8) ,
344	 => std_logic_vector(to_unsigned(100,8) ,
345	 => std_logic_vector(to_unsigned(108,8) ,
346	 => std_logic_vector(to_unsigned(101,8) ,
347	 => std_logic_vector(to_unsigned(107,8) ,
348	 => std_logic_vector(to_unsigned(107,8) ,
349	 => std_logic_vector(to_unsigned(107,8) ,
350	 => std_logic_vector(to_unsigned(107,8) ,
351	 => std_logic_vector(to_unsigned(107,8) ,
352	 => std_logic_vector(to_unsigned(104,8) ,
353	 => std_logic_vector(to_unsigned(104,8) ,
354	 => std_logic_vector(to_unsigned(109,8) ,
355	 => std_logic_vector(to_unsigned(111,8) ,
356	 => std_logic_vector(to_unsigned(109,8) ,
357	 => std_logic_vector(to_unsigned(109,8) ,
358	 => std_logic_vector(to_unsigned(108,8) ,
359	 => std_logic_vector(to_unsigned(116,8) ,
360	 => std_logic_vector(to_unsigned(119,8) ,
361	 => std_logic_vector(to_unsigned(114,8) ,
362	 => std_logic_vector(to_unsigned(114,8) ,
363	 => std_logic_vector(to_unsigned(112,8) ,
364	 => std_logic_vector(to_unsigned(112,8) ,
365	 => std_logic_vector(to_unsigned(115,8) ,
366	 => std_logic_vector(to_unsigned(115,8) ,
367	 => std_logic_vector(to_unsigned(114,8) ,
368	 => std_logic_vector(to_unsigned(115,8) ,
369	 => std_logic_vector(to_unsigned(116,8) ,
370	 => std_logic_vector(to_unsigned(115,8) ,
371	 => std_logic_vector(to_unsigned(118,8) ,
372	 => std_logic_vector(to_unsigned(114,8) ,
373	 => std_logic_vector(to_unsigned(105,8) ,
374	 => std_logic_vector(to_unsigned(114,8) ,
375	 => std_logic_vector(to_unsigned(116,8) ,
376	 => std_logic_vector(to_unsigned(112,8) ,
377	 => std_logic_vector(to_unsigned(115,8) ,
378	 => std_logic_vector(to_unsigned(119,8) ,
379	 => std_logic_vector(to_unsigned(112,8) ,
380	 => std_logic_vector(to_unsigned(100,8) ,
381	 => std_logic_vector(to_unsigned(99,8) ,
382	 => std_logic_vector(to_unsigned(109,8) ,
383	 => std_logic_vector(to_unsigned(116,8) ,
384	 => std_logic_vector(to_unsigned(115,8) ,
385	 => std_logic_vector(to_unsigned(119,8) ,
386	 => std_logic_vector(to_unsigned(119,8) ,
387	 => std_logic_vector(to_unsigned(115,8) ,
388	 => std_logic_vector(to_unsigned(114,8) ,
389	 => std_logic_vector(to_unsigned(116,8) ,
390	 => std_logic_vector(to_unsigned(116,8) ,
391	 => std_logic_vector(to_unsigned(114,8) ,
392	 => std_logic_vector(to_unsigned(116,8) ,
393	 => std_logic_vector(to_unsigned(114,8) ,
394	 => std_logic_vector(to_unsigned(115,8) ,
395	 => std_logic_vector(to_unsigned(114,8) ,
396	 => std_logic_vector(to_unsigned(111,8) ,
397	 => std_logic_vector(to_unsigned(115,8) ,
398	 => std_logic_vector(to_unsigned(112,8) ,
399	 => std_logic_vector(to_unsigned(107,8) ,
400	 => std_logic_vector(to_unsigned(109,8) ,
401	 => std_logic_vector(to_unsigned(114,8) ,
402	 => std_logic_vector(to_unsigned(111,8) ,
403	 => std_logic_vector(to_unsigned(115,8) ,
404	 => std_logic_vector(to_unsigned(112,8) ,
405	 => std_logic_vector(to_unsigned(115,8) ,
406	 => std_logic_vector(to_unsigned(119,8) ,
407	 => std_logic_vector(to_unsigned(109,8) ,
408	 => std_logic_vector(to_unsigned(111,8) ,
409	 => std_logic_vector(to_unsigned(111,8) ,
410	 => std_logic_vector(to_unsigned(108,8) ,
411	 => std_logic_vector(to_unsigned(111,8) ,
412	 => std_logic_vector(to_unsigned(108,8) ,
413	 => std_logic_vector(to_unsigned(105,8) ,
414	 => std_logic_vector(to_unsigned(101,8) ,
415	 => std_logic_vector(to_unsigned(101,8) ,
416	 => std_logic_vector(to_unsigned(105,8) ,
417	 => std_logic_vector(to_unsigned(108,8) ,
418	 => std_logic_vector(to_unsigned(103,8) ,
419	 => std_logic_vector(to_unsigned(105,8) ,
420	 => std_logic_vector(to_unsigned(107,8) ,
421	 => std_logic_vector(to_unsigned(108,8) ,
422	 => std_logic_vector(to_unsigned(109,8) ,
423	 => std_logic_vector(to_unsigned(108,8) ,
424	 => std_logic_vector(to_unsigned(107,8) ,
425	 => std_logic_vector(to_unsigned(108,8) ,
426	 => std_logic_vector(to_unsigned(108,8) ,
427	 => std_logic_vector(to_unsigned(104,8) ,
428	 => std_logic_vector(to_unsigned(111,8) ,
429	 => std_logic_vector(to_unsigned(114,8) ,
430	 => std_logic_vector(to_unsigned(108,8) ,
431	 => std_logic_vector(to_unsigned(104,8) ,
432	 => std_logic_vector(to_unsigned(107,8) ,
433	 => std_logic_vector(to_unsigned(108,8) ,
434	 => std_logic_vector(to_unsigned(107,8) ,
435	 => std_logic_vector(to_unsigned(114,8) ,
436	 => std_logic_vector(to_unsigned(114,8) ,
437	 => std_logic_vector(to_unsigned(105,8) ,
438	 => std_logic_vector(to_unsigned(101,8) ,
439	 => std_logic_vector(to_unsigned(103,8) ,
440	 => std_logic_vector(to_unsigned(107,8) ,
441	 => std_logic_vector(to_unsigned(107,8) ,
442	 => std_logic_vector(to_unsigned(103,8) ,
443	 => std_logic_vector(to_unsigned(100,8) ,
444	 => std_logic_vector(to_unsigned(103,8) ,
445	 => std_logic_vector(to_unsigned(100,8) ,
446	 => std_logic_vector(to_unsigned(97,8) ,
447	 => std_logic_vector(to_unsigned(100,8) ,
448	 => std_logic_vector(to_unsigned(101,8) ,
449	 => std_logic_vector(to_unsigned(97,8) ,
450	 => std_logic_vector(to_unsigned(97,8) ,
451	 => std_logic_vector(to_unsigned(99,8) ,
452	 => std_logic_vector(to_unsigned(97,8) ,
453	 => std_logic_vector(to_unsigned(100,8) ,
454	 => std_logic_vector(to_unsigned(101,8) ,
455	 => std_logic_vector(to_unsigned(101,8) ,
456	 => std_logic_vector(to_unsigned(103,8) ,
457	 => std_logic_vector(to_unsigned(101,8) ,
458	 => std_logic_vector(to_unsigned(100,8) ,
459	 => std_logic_vector(to_unsigned(99,8) ,
460	 => std_logic_vector(to_unsigned(97,8) ,
461	 => std_logic_vector(to_unsigned(100,8) ,
462	 => std_logic_vector(to_unsigned(103,8) ,
463	 => std_logic_vector(to_unsigned(101,8) ,
464	 => std_logic_vector(to_unsigned(104,8) ,
465	 => std_logic_vector(to_unsigned(103,8) ,
466	 => std_logic_vector(to_unsigned(104,8) ,
467	 => std_logic_vector(to_unsigned(105,8) ,
468	 => std_logic_vector(to_unsigned(107,8) ,
469	 => std_logic_vector(to_unsigned(103,8) ,
470	 => std_logic_vector(to_unsigned(107,8) ,
471	 => std_logic_vector(to_unsigned(97,8) ,
472	 => std_logic_vector(to_unsigned(96,8) ,
473	 => std_logic_vector(to_unsigned(99,8) ,
474	 => std_logic_vector(to_unsigned(95,8) ,
475	 => std_logic_vector(to_unsigned(96,8) ,
476	 => std_logic_vector(to_unsigned(93,8) ,
477	 => std_logic_vector(to_unsigned(91,8) ,
478	 => std_logic_vector(to_unsigned(88,8) ,
479	 => std_logic_vector(to_unsigned(92,8) ,
480	 => std_logic_vector(to_unsigned(91,8) ,
481	 => std_logic_vector(to_unsigned(87,8) ,
482	 => std_logic_vector(to_unsigned(93,8) ,
483	 => std_logic_vector(to_unsigned(95,8) ,
484	 => std_logic_vector(to_unsigned(93,8) ,
485	 => std_logic_vector(to_unsigned(92,8) ,
486	 => std_logic_vector(to_unsigned(90,8) ,
487	 => std_logic_vector(to_unsigned(87,8) ,
488	 => std_logic_vector(to_unsigned(88,8) ,
489	 => std_logic_vector(to_unsigned(90,8) ,
490	 => std_logic_vector(to_unsigned(88,8) ,
491	 => std_logic_vector(to_unsigned(92,8) ,
492	 => std_logic_vector(to_unsigned(96,8) ,
493	 => std_logic_vector(to_unsigned(93,8) ,
494	 => std_logic_vector(to_unsigned(90,8) ,
495	 => std_logic_vector(to_unsigned(88,8) ,
496	 => std_logic_vector(to_unsigned(91,8) ,
497	 => std_logic_vector(to_unsigned(90,8) ,
498	 => std_logic_vector(to_unsigned(87,8) ,
499	 => std_logic_vector(to_unsigned(91,8) ,
500	 => std_logic_vector(to_unsigned(86,8) ,
501	 => std_logic_vector(to_unsigned(84,8) ,
502	 => std_logic_vector(to_unsigned(85,8) ,
503	 => std_logic_vector(to_unsigned(88,8) ,
504	 => std_logic_vector(to_unsigned(92,8) ,
505	 => std_logic_vector(to_unsigned(90,8) ,
506	 => std_logic_vector(to_unsigned(90,8) ,
507	 => std_logic_vector(to_unsigned(88,8) ,
508	 => std_logic_vector(to_unsigned(88,8) ,
509	 => std_logic_vector(to_unsigned(91,8) ,
510	 => std_logic_vector(to_unsigned(90,8) ,
511	 => std_logic_vector(to_unsigned(87,8) ,
512	 => std_logic_vector(to_unsigned(85,8) ,
513	 => std_logic_vector(to_unsigned(85,8) ,
514	 => std_logic_vector(to_unsigned(90,8) ,
515	 => std_logic_vector(to_unsigned(91,8) ,
516	 => std_logic_vector(to_unsigned(88,8) ,
517	 => std_logic_vector(to_unsigned(88,8) ,
518	 => std_logic_vector(to_unsigned(86,8) ,
519	 => std_logic_vector(to_unsigned(90,8) ,
520	 => std_logic_vector(to_unsigned(90,8) ,
521	 => std_logic_vector(to_unsigned(88,8) ,
522	 => std_logic_vector(to_unsigned(91,8) ,
523	 => std_logic_vector(to_unsigned(87,8) ,
524	 => std_logic_vector(to_unsigned(85,8) ,
525	 => std_logic_vector(to_unsigned(90,8) ,
526	 => std_logic_vector(to_unsigned(91,8) ,
527	 => std_logic_vector(to_unsigned(92,8) ,
528	 => std_logic_vector(to_unsigned(90,8) ,
529	 => std_logic_vector(to_unsigned(91,8) ,
530	 => std_logic_vector(to_unsigned(96,8) ,
531	 => std_logic_vector(to_unsigned(97,8) ,
532	 => std_logic_vector(to_unsigned(96,8) ,
533	 => std_logic_vector(to_unsigned(96,8) ,
534	 => std_logic_vector(to_unsigned(95,8) ,
535	 => std_logic_vector(to_unsigned(90,8) ,
536	 => std_logic_vector(to_unsigned(91,8) ,
537	 => std_logic_vector(to_unsigned(90,8) ,
538	 => std_logic_vector(to_unsigned(87,8) ,
539	 => std_logic_vector(to_unsigned(91,8) ,
540	 => std_logic_vector(to_unsigned(91,8) ,
541	 => std_logic_vector(to_unsigned(93,8) ,
542	 => std_logic_vector(to_unsigned(90,8) ,
543	 => std_logic_vector(to_unsigned(88,8) ,
544	 => std_logic_vector(to_unsigned(93,8) ,
545	 => std_logic_vector(to_unsigned(99,8) ,
546	 => std_logic_vector(to_unsigned(96,8) ,
547	 => std_logic_vector(to_unsigned(97,8) ,
548	 => std_logic_vector(to_unsigned(93,8) ,
549	 => std_logic_vector(to_unsigned(95,8) ,
550	 => std_logic_vector(to_unsigned(95,8) ,
551	 => std_logic_vector(to_unsigned(95,8) ,
552	 => std_logic_vector(to_unsigned(97,8) ,
553	 => std_logic_vector(to_unsigned(95,8) ,
554	 => std_logic_vector(to_unsigned(96,8) ,
555	 => std_logic_vector(to_unsigned(21,8) ,
556	 => std_logic_vector(to_unsigned(0,8) ,
557	 => std_logic_vector(to_unsigned(0,8) ,
558	 => std_logic_vector(to_unsigned(4,8) ,
559	 => std_logic_vector(to_unsigned(81,8) ,
560	 => std_logic_vector(to_unsigned(97,8) ,
561	 => std_logic_vector(to_unsigned(88,8) ,
562	 => std_logic_vector(to_unsigned(91,8) ,
563	 => std_logic_vector(to_unsigned(93,8) ,
564	 => std_logic_vector(to_unsigned(93,8) ,
565	 => std_logic_vector(to_unsigned(92,8) ,
566	 => std_logic_vector(to_unsigned(95,8) ,
567	 => std_logic_vector(to_unsigned(101,8) ,
568	 => std_logic_vector(to_unsigned(108,8) ,
569	 => std_logic_vector(to_unsigned(112,8) ,
570	 => std_logic_vector(to_unsigned(111,8) ,
571	 => std_logic_vector(to_unsigned(105,8) ,
572	 => std_logic_vector(to_unsigned(100,8) ,
573	 => std_logic_vector(to_unsigned(109,8) ,
574	 => std_logic_vector(to_unsigned(112,8) ,
575	 => std_logic_vector(to_unsigned(111,8) ,
576	 => std_logic_vector(to_unsigned(111,8) ,
577	 => std_logic_vector(to_unsigned(111,8) ,
578	 => std_logic_vector(to_unsigned(116,8) ,
579	 => std_logic_vector(to_unsigned(114,8) ,
580	 => std_logic_vector(to_unsigned(111,8) ,
581	 => std_logic_vector(to_unsigned(112,8) ,
582	 => std_logic_vector(to_unsigned(112,8) ,
583	 => std_logic_vector(to_unsigned(116,8) ,
584	 => std_logic_vector(to_unsigned(114,8) ,
585	 => std_logic_vector(to_unsigned(111,8) ,
586	 => std_logic_vector(to_unsigned(108,8) ,
587	 => std_logic_vector(to_unsigned(108,8) ,
588	 => std_logic_vector(to_unsigned(112,8) ,
589	 => std_logic_vector(to_unsigned(115,8) ,
590	 => std_logic_vector(to_unsigned(118,8) ,
591	 => std_logic_vector(to_unsigned(119,8) ,
592	 => std_logic_vector(to_unsigned(118,8) ,
593	 => std_logic_vector(to_unsigned(122,8) ,
594	 => std_logic_vector(to_unsigned(127,8) ,
595	 => std_logic_vector(to_unsigned(130,8) ,
596	 => std_logic_vector(to_unsigned(133,8) ,
597	 => std_logic_vector(to_unsigned(136,8) ,
598	 => std_logic_vector(to_unsigned(136,8) ,
599	 => std_logic_vector(to_unsigned(139,8) ,
600	 => std_logic_vector(to_unsigned(139,8) ,
601	 => std_logic_vector(to_unsigned(144,8) ,
602	 => std_logic_vector(to_unsigned(144,8) ,
603	 => std_logic_vector(to_unsigned(149,8) ,
604	 => std_logic_vector(to_unsigned(154,8) ,
605	 => std_logic_vector(to_unsigned(154,8) ,
606	 => std_logic_vector(to_unsigned(152,8) ,
607	 => std_logic_vector(to_unsigned(149,8) ,
608	 => std_logic_vector(to_unsigned(147,8) ,
609	 => std_logic_vector(to_unsigned(152,8) ,
610	 => std_logic_vector(to_unsigned(154,8) ,
611	 => std_logic_vector(to_unsigned(154,8) ,
612	 => std_logic_vector(to_unsigned(154,8) ,
613	 => std_logic_vector(to_unsigned(156,8) ,
614	 => std_logic_vector(to_unsigned(157,8) ,
615	 => std_logic_vector(to_unsigned(159,8) ,
616	 => std_logic_vector(to_unsigned(159,8) ,
617	 => std_logic_vector(to_unsigned(157,8) ,
618	 => std_logic_vector(to_unsigned(159,8) ,
619	 => std_logic_vector(to_unsigned(161,8) ,
620	 => std_logic_vector(to_unsigned(161,8) ,
621	 => std_logic_vector(to_unsigned(156,8) ,
622	 => std_logic_vector(to_unsigned(156,8) ,
623	 => std_logic_vector(to_unsigned(163,8) ,
624	 => std_logic_vector(to_unsigned(161,8) ,
625	 => std_logic_vector(to_unsigned(159,8) ,
626	 => std_logic_vector(to_unsigned(161,8) ,
627	 => std_logic_vector(to_unsigned(159,8) ,
628	 => std_logic_vector(to_unsigned(161,8) ,
629	 => std_logic_vector(to_unsigned(164,8) ,
630	 => std_logic_vector(to_unsigned(164,8) ,
631	 => std_logic_vector(to_unsigned(166,8) ,
632	 => std_logic_vector(to_unsigned(163,8) ,
633	 => std_logic_vector(to_unsigned(161,8) ,
634	 => std_logic_vector(to_unsigned(164,8) ,
635	 => std_logic_vector(to_unsigned(166,8) ,
636	 => std_logic_vector(to_unsigned(164,8) ,
637	 => std_logic_vector(to_unsigned(159,8) ,
638	 => std_logic_vector(to_unsigned(159,8) ,
639	 => std_logic_vector(to_unsigned(163,8) ,
640	 => std_logic_vector(to_unsigned(163,8) ,
641	 => std_logic_vector(to_unsigned(108,8) ,
642	 => std_logic_vector(to_unsigned(107,8) ,
643	 => std_logic_vector(to_unsigned(107,8) ,
644	 => std_logic_vector(to_unsigned(105,8) ,
645	 => std_logic_vector(to_unsigned(101,8) ,
646	 => std_logic_vector(to_unsigned(105,8) ,
647	 => std_logic_vector(to_unsigned(109,8) ,
648	 => std_logic_vector(to_unsigned(105,8) ,
649	 => std_logic_vector(to_unsigned(101,8) ,
650	 => std_logic_vector(to_unsigned(97,8) ,
651	 => std_logic_vector(to_unsigned(99,8) ,
652	 => std_logic_vector(to_unsigned(104,8) ,
653	 => std_logic_vector(to_unsigned(105,8) ,
654	 => std_logic_vector(to_unsigned(95,8) ,
655	 => std_logic_vector(to_unsigned(93,8) ,
656	 => std_logic_vector(to_unsigned(93,8) ,
657	 => std_logic_vector(to_unsigned(92,8) ,
658	 => std_logic_vector(to_unsigned(92,8) ,
659	 => std_logic_vector(to_unsigned(90,8) ,
660	 => std_logic_vector(to_unsigned(90,8) ,
661	 => std_logic_vector(to_unsigned(90,8) ,
662	 => std_logic_vector(to_unsigned(92,8) ,
663	 => std_logic_vector(to_unsigned(96,8) ,
664	 => std_logic_vector(to_unsigned(104,8) ,
665	 => std_logic_vector(to_unsigned(105,8) ,
666	 => std_logic_vector(to_unsigned(104,8) ,
667	 => std_logic_vector(to_unsigned(111,8) ,
668	 => std_logic_vector(to_unsigned(108,8) ,
669	 => std_logic_vector(to_unsigned(105,8) ,
670	 => std_logic_vector(to_unsigned(100,8) ,
671	 => std_logic_vector(to_unsigned(105,8) ,
672	 => std_logic_vector(to_unsigned(104,8) ,
673	 => std_logic_vector(to_unsigned(101,8) ,
674	 => std_logic_vector(to_unsigned(105,8) ,
675	 => std_logic_vector(to_unsigned(107,8) ,
676	 => std_logic_vector(to_unsigned(105,8) ,
677	 => std_logic_vector(to_unsigned(104,8) ,
678	 => std_logic_vector(to_unsigned(100,8) ,
679	 => std_logic_vector(to_unsigned(105,8) ,
680	 => std_logic_vector(to_unsigned(111,8) ,
681	 => std_logic_vector(to_unsigned(108,8) ,
682	 => std_logic_vector(to_unsigned(112,8) ,
683	 => std_logic_vector(to_unsigned(112,8) ,
684	 => std_logic_vector(to_unsigned(109,8) ,
685	 => std_logic_vector(to_unsigned(111,8) ,
686	 => std_logic_vector(to_unsigned(112,8) ,
687	 => std_logic_vector(to_unsigned(111,8) ,
688	 => std_logic_vector(to_unsigned(108,8) ,
689	 => std_logic_vector(to_unsigned(112,8) ,
690	 => std_logic_vector(to_unsigned(119,8) ,
691	 => std_logic_vector(to_unsigned(115,8) ,
692	 => std_logic_vector(to_unsigned(108,8) ,
693	 => std_logic_vector(to_unsigned(111,8) ,
694	 => std_logic_vector(to_unsigned(116,8) ,
695	 => std_logic_vector(to_unsigned(108,8) ,
696	 => std_logic_vector(to_unsigned(108,8) ,
697	 => std_logic_vector(to_unsigned(116,8) ,
698	 => std_logic_vector(to_unsigned(112,8) ,
699	 => std_logic_vector(to_unsigned(107,8) ,
700	 => std_logic_vector(to_unsigned(100,8) ,
701	 => std_logic_vector(to_unsigned(101,8) ,
702	 => std_logic_vector(to_unsigned(108,8) ,
703	 => std_logic_vector(to_unsigned(109,8) ,
704	 => std_logic_vector(to_unsigned(111,8) ,
705	 => std_logic_vector(to_unsigned(118,8) ,
706	 => std_logic_vector(to_unsigned(119,8) ,
707	 => std_logic_vector(to_unsigned(112,8) ,
708	 => std_logic_vector(to_unsigned(114,8) ,
709	 => std_logic_vector(to_unsigned(118,8) ,
710	 => std_logic_vector(to_unsigned(118,8) ,
711	 => std_logic_vector(to_unsigned(118,8) ,
712	 => std_logic_vector(to_unsigned(119,8) ,
713	 => std_logic_vector(to_unsigned(116,8) ,
714	 => std_logic_vector(to_unsigned(118,8) ,
715	 => std_logic_vector(to_unsigned(111,8) ,
716	 => std_logic_vector(to_unsigned(108,8) ,
717	 => std_logic_vector(to_unsigned(112,8) ,
718	 => std_logic_vector(to_unsigned(114,8) ,
719	 => std_logic_vector(to_unsigned(114,8) ,
720	 => std_logic_vector(to_unsigned(112,8) ,
721	 => std_logic_vector(to_unsigned(114,8) ,
722	 => std_logic_vector(to_unsigned(109,8) ,
723	 => std_logic_vector(to_unsigned(111,8) ,
724	 => std_logic_vector(to_unsigned(108,8) ,
725	 => std_logic_vector(to_unsigned(111,8) ,
726	 => std_logic_vector(to_unsigned(119,8) ,
727	 => std_logic_vector(to_unsigned(114,8) ,
728	 => std_logic_vector(to_unsigned(109,8) ,
729	 => std_logic_vector(to_unsigned(111,8) ,
730	 => std_logic_vector(to_unsigned(115,8) ,
731	 => std_logic_vector(to_unsigned(114,8) ,
732	 => std_logic_vector(to_unsigned(107,8) ,
733	 => std_logic_vector(to_unsigned(104,8) ,
734	 => std_logic_vector(to_unsigned(107,8) ,
735	 => std_logic_vector(to_unsigned(105,8) ,
736	 => std_logic_vector(to_unsigned(104,8) ,
737	 => std_logic_vector(to_unsigned(104,8) ,
738	 => std_logic_vector(to_unsigned(103,8) ,
739	 => std_logic_vector(to_unsigned(104,8) ,
740	 => std_logic_vector(to_unsigned(101,8) ,
741	 => std_logic_vector(to_unsigned(104,8) ,
742	 => std_logic_vector(to_unsigned(105,8) ,
743	 => std_logic_vector(to_unsigned(108,8) ,
744	 => std_logic_vector(to_unsigned(105,8) ,
745	 => std_logic_vector(to_unsigned(105,8) ,
746	 => std_logic_vector(to_unsigned(109,8) ,
747	 => std_logic_vector(to_unsigned(114,8) ,
748	 => std_logic_vector(to_unsigned(116,8) ,
749	 => std_logic_vector(to_unsigned(114,8) ,
750	 => std_logic_vector(to_unsigned(108,8) ,
751	 => std_logic_vector(to_unsigned(105,8) ,
752	 => std_logic_vector(to_unsigned(112,8) ,
753	 => std_logic_vector(to_unsigned(107,8) ,
754	 => std_logic_vector(to_unsigned(104,8) ,
755	 => std_logic_vector(to_unsigned(111,8) ,
756	 => std_logic_vector(to_unsigned(109,8) ,
757	 => std_logic_vector(to_unsigned(105,8) ,
758	 => std_logic_vector(to_unsigned(103,8) ,
759	 => std_logic_vector(to_unsigned(104,8) ,
760	 => std_logic_vector(to_unsigned(105,8) ,
761	 => std_logic_vector(to_unsigned(105,8) ,
762	 => std_logic_vector(to_unsigned(99,8) ,
763	 => std_logic_vector(to_unsigned(101,8) ,
764	 => std_logic_vector(to_unsigned(105,8) ,
765	 => std_logic_vector(to_unsigned(103,8) ,
766	 => std_logic_vector(to_unsigned(100,8) ,
767	 => std_logic_vector(to_unsigned(100,8) ,
768	 => std_logic_vector(to_unsigned(101,8) ,
769	 => std_logic_vector(to_unsigned(100,8) ,
770	 => std_logic_vector(to_unsigned(97,8) ,
771	 => std_logic_vector(to_unsigned(95,8) ,
772	 => std_logic_vector(to_unsigned(96,8) ,
773	 => std_logic_vector(to_unsigned(97,8) ,
774	 => std_logic_vector(to_unsigned(97,8) ,
775	 => std_logic_vector(to_unsigned(97,8) ,
776	 => std_logic_vector(to_unsigned(99,8) ,
777	 => std_logic_vector(to_unsigned(100,8) ,
778	 => std_logic_vector(to_unsigned(101,8) ,
779	 => std_logic_vector(to_unsigned(99,8) ,
780	 => std_logic_vector(to_unsigned(95,8) ,
781	 => std_logic_vector(to_unsigned(100,8) ,
782	 => std_logic_vector(to_unsigned(103,8) ,
783	 => std_logic_vector(to_unsigned(99,8) ,
784	 => std_logic_vector(to_unsigned(101,8) ,
785	 => std_logic_vector(to_unsigned(100,8) ,
786	 => std_logic_vector(to_unsigned(103,8) ,
787	 => std_logic_vector(to_unsigned(109,8) ,
788	 => std_logic_vector(to_unsigned(107,8) ,
789	 => std_logic_vector(to_unsigned(100,8) ,
790	 => std_logic_vector(to_unsigned(103,8) ,
791	 => std_logic_vector(to_unsigned(101,8) ,
792	 => std_logic_vector(to_unsigned(97,8) ,
793	 => std_logic_vector(to_unsigned(99,8) ,
794	 => std_logic_vector(to_unsigned(95,8) ,
795	 => std_logic_vector(to_unsigned(91,8) ,
796	 => std_logic_vector(to_unsigned(93,8) ,
797	 => std_logic_vector(to_unsigned(88,8) ,
798	 => std_logic_vector(to_unsigned(86,8) ,
799	 => std_logic_vector(to_unsigned(90,8) ,
800	 => std_logic_vector(to_unsigned(87,8) ,
801	 => std_logic_vector(to_unsigned(87,8) ,
802	 => std_logic_vector(to_unsigned(92,8) ,
803	 => std_logic_vector(to_unsigned(92,8) ,
804	 => std_logic_vector(to_unsigned(90,8) ,
805	 => std_logic_vector(to_unsigned(88,8) ,
806	 => std_logic_vector(to_unsigned(86,8) ,
807	 => std_logic_vector(to_unsigned(84,8) ,
808	 => std_logic_vector(to_unsigned(84,8) ,
809	 => std_logic_vector(to_unsigned(84,8) ,
810	 => std_logic_vector(to_unsigned(86,8) ,
811	 => std_logic_vector(to_unsigned(90,8) ,
812	 => std_logic_vector(to_unsigned(95,8) ,
813	 => std_logic_vector(to_unsigned(92,8) ,
814	 => std_logic_vector(to_unsigned(88,8) ,
815	 => std_logic_vector(to_unsigned(86,8) ,
816	 => std_logic_vector(to_unsigned(88,8) ,
817	 => std_logic_vector(to_unsigned(90,8) ,
818	 => std_logic_vector(to_unsigned(85,8) ,
819	 => std_logic_vector(to_unsigned(91,8) ,
820	 => std_logic_vector(to_unsigned(88,8) ,
821	 => std_logic_vector(to_unsigned(86,8) ,
822	 => std_logic_vector(to_unsigned(84,8) ,
823	 => std_logic_vector(to_unsigned(84,8) ,
824	 => std_logic_vector(to_unsigned(87,8) ,
825	 => std_logic_vector(to_unsigned(88,8) ,
826	 => std_logic_vector(to_unsigned(91,8) ,
827	 => std_logic_vector(to_unsigned(86,8) ,
828	 => std_logic_vector(to_unsigned(85,8) ,
829	 => std_logic_vector(to_unsigned(87,8) ,
830	 => std_logic_vector(to_unsigned(87,8) ,
831	 => std_logic_vector(to_unsigned(85,8) ,
832	 => std_logic_vector(to_unsigned(82,8) ,
833	 => std_logic_vector(to_unsigned(85,8) ,
834	 => std_logic_vector(to_unsigned(88,8) ,
835	 => std_logic_vector(to_unsigned(87,8) ,
836	 => std_logic_vector(to_unsigned(87,8) ,
837	 => std_logic_vector(to_unsigned(87,8) ,
838	 => std_logic_vector(to_unsigned(85,8) ,
839	 => std_logic_vector(to_unsigned(90,8) ,
840	 => std_logic_vector(to_unsigned(93,8) ,
841	 => std_logic_vector(to_unsigned(93,8) ,
842	 => std_logic_vector(to_unsigned(91,8) ,
843	 => std_logic_vector(to_unsigned(86,8) ,
844	 => std_logic_vector(to_unsigned(80,8) ,
845	 => std_logic_vector(to_unsigned(85,8) ,
846	 => std_logic_vector(to_unsigned(90,8) ,
847	 => std_logic_vector(to_unsigned(85,8) ,
848	 => std_logic_vector(to_unsigned(85,8) ,
849	 => std_logic_vector(to_unsigned(86,8) ,
850	 => std_logic_vector(to_unsigned(86,8) ,
851	 => std_logic_vector(to_unsigned(88,8) ,
852	 => std_logic_vector(to_unsigned(95,8) ,
853	 => std_logic_vector(to_unsigned(93,8) ,
854	 => std_logic_vector(to_unsigned(90,8) ,
855	 => std_logic_vector(to_unsigned(87,8) ,
856	 => std_logic_vector(to_unsigned(88,8) ,
857	 => std_logic_vector(to_unsigned(87,8) ,
858	 => std_logic_vector(to_unsigned(87,8) ,
859	 => std_logic_vector(to_unsigned(90,8) ,
860	 => std_logic_vector(to_unsigned(88,8) ,
861	 => std_logic_vector(to_unsigned(91,8) ,
862	 => std_logic_vector(to_unsigned(92,8) ,
863	 => std_logic_vector(to_unsigned(87,8) ,
864	 => std_logic_vector(to_unsigned(92,8) ,
865	 => std_logic_vector(to_unsigned(99,8) ,
866	 => std_logic_vector(to_unsigned(93,8) ,
867	 => std_logic_vector(to_unsigned(92,8) ,
868	 => std_logic_vector(to_unsigned(86,8) ,
869	 => std_logic_vector(to_unsigned(92,8) ,
870	 => std_logic_vector(to_unsigned(97,8) ,
871	 => std_logic_vector(to_unsigned(99,8) ,
872	 => std_logic_vector(to_unsigned(95,8) ,
873	 => std_logic_vector(to_unsigned(88,8) ,
874	 => std_logic_vector(to_unsigned(101,8) ,
875	 => std_logic_vector(to_unsigned(40,8) ,
876	 => std_logic_vector(to_unsigned(1,8) ,
877	 => std_logic_vector(to_unsigned(0,8) ,
878	 => std_logic_vector(to_unsigned(1,8) ,
879	 => std_logic_vector(to_unsigned(54,8) ,
880	 => std_logic_vector(to_unsigned(105,8) ,
881	 => std_logic_vector(to_unsigned(87,8) ,
882	 => std_logic_vector(to_unsigned(92,8) ,
883	 => std_logic_vector(to_unsigned(90,8) ,
884	 => std_logic_vector(to_unsigned(90,8) ,
885	 => std_logic_vector(to_unsigned(92,8) ,
886	 => std_logic_vector(to_unsigned(93,8) ,
887	 => std_logic_vector(to_unsigned(99,8) ,
888	 => std_logic_vector(to_unsigned(101,8) ,
889	 => std_logic_vector(to_unsigned(103,8) ,
890	 => std_logic_vector(to_unsigned(107,8) ,
891	 => std_logic_vector(to_unsigned(111,8) ,
892	 => std_logic_vector(to_unsigned(109,8) ,
893	 => std_logic_vector(to_unsigned(114,8) ,
894	 => std_logic_vector(to_unsigned(107,8) ,
895	 => std_logic_vector(to_unsigned(104,8) ,
896	 => std_logic_vector(to_unsigned(108,8) ,
897	 => std_logic_vector(to_unsigned(111,8) ,
898	 => std_logic_vector(to_unsigned(115,8) ,
899	 => std_logic_vector(to_unsigned(109,8) ,
900	 => std_logic_vector(to_unsigned(105,8) ,
901	 => std_logic_vector(to_unsigned(109,8) ,
902	 => std_logic_vector(to_unsigned(111,8) ,
903	 => std_logic_vector(to_unsigned(112,8) ,
904	 => std_logic_vector(to_unsigned(115,8) ,
905	 => std_logic_vector(to_unsigned(109,8) ,
906	 => std_logic_vector(to_unsigned(107,8) ,
907	 => std_logic_vector(to_unsigned(111,8) ,
908	 => std_logic_vector(to_unsigned(112,8) ,
909	 => std_logic_vector(to_unsigned(115,8) ,
910	 => std_logic_vector(to_unsigned(118,8) ,
911	 => std_logic_vector(to_unsigned(119,8) ,
912	 => std_logic_vector(to_unsigned(118,8) ,
913	 => std_logic_vector(to_unsigned(118,8) ,
914	 => std_logic_vector(to_unsigned(124,8) ,
915	 => std_logic_vector(to_unsigned(128,8) ,
916	 => std_logic_vector(to_unsigned(134,8) ,
917	 => std_logic_vector(to_unsigned(136,8) ,
918	 => std_logic_vector(to_unsigned(141,8) ,
919	 => std_logic_vector(to_unsigned(149,8) ,
920	 => std_logic_vector(to_unsigned(142,8) ,
921	 => std_logic_vector(to_unsigned(141,8) ,
922	 => std_logic_vector(to_unsigned(142,8) ,
923	 => std_logic_vector(to_unsigned(144,8) ,
924	 => std_logic_vector(to_unsigned(152,8) ,
925	 => std_logic_vector(to_unsigned(157,8) ,
926	 => std_logic_vector(to_unsigned(152,8) ,
927	 => std_logic_vector(to_unsigned(147,8) ,
928	 => std_logic_vector(to_unsigned(147,8) ,
929	 => std_logic_vector(to_unsigned(151,8) ,
930	 => std_logic_vector(to_unsigned(149,8) ,
931	 => std_logic_vector(to_unsigned(149,8) ,
932	 => std_logic_vector(to_unsigned(149,8) ,
933	 => std_logic_vector(to_unsigned(151,8) ,
934	 => std_logic_vector(to_unsigned(154,8) ,
935	 => std_logic_vector(to_unsigned(159,8) ,
936	 => std_logic_vector(to_unsigned(159,8) ,
937	 => std_logic_vector(to_unsigned(157,8) ,
938	 => std_logic_vector(to_unsigned(159,8) ,
939	 => std_logic_vector(to_unsigned(161,8) ,
940	 => std_logic_vector(to_unsigned(163,8) ,
941	 => std_logic_vector(to_unsigned(161,8) ,
942	 => std_logic_vector(to_unsigned(159,8) ,
943	 => std_logic_vector(to_unsigned(161,8) ,
944	 => std_logic_vector(to_unsigned(163,8) ,
945	 => std_logic_vector(to_unsigned(163,8) ,
946	 => std_logic_vector(to_unsigned(163,8) ,
947	 => std_logic_vector(to_unsigned(163,8) ,
948	 => std_logic_vector(to_unsigned(164,8) ,
949	 => std_logic_vector(to_unsigned(164,8) ,
950	 => std_logic_vector(to_unsigned(163,8) ,
951	 => std_logic_vector(to_unsigned(163,8) ,
952	 => std_logic_vector(to_unsigned(161,8) ,
953	 => std_logic_vector(to_unsigned(161,8) ,
954	 => std_logic_vector(to_unsigned(164,8) ,
955	 => std_logic_vector(to_unsigned(164,8) ,
956	 => std_logic_vector(to_unsigned(164,8) ,
957	 => std_logic_vector(to_unsigned(163,8) ,
958	 => std_logic_vector(to_unsigned(163,8) ,
959	 => std_logic_vector(to_unsigned(164,8) ,
960	 => std_logic_vector(to_unsigned(163,8) ,
961	 => std_logic_vector(to_unsigned(100,8) ,
962	 => std_logic_vector(to_unsigned(104,8) ,
963	 => std_logic_vector(to_unsigned(104,8) ,
964	 => std_logic_vector(to_unsigned(99,8) ,
965	 => std_logic_vector(to_unsigned(101,8) ,
966	 => std_logic_vector(to_unsigned(107,8) ,
967	 => std_logic_vector(to_unsigned(108,8) ,
968	 => std_logic_vector(to_unsigned(107,8) ,
969	 => std_logic_vector(to_unsigned(103,8) ,
970	 => std_logic_vector(to_unsigned(101,8) ,
971	 => std_logic_vector(to_unsigned(101,8) ,
972	 => std_logic_vector(to_unsigned(97,8) ,
973	 => std_logic_vector(to_unsigned(99,8) ,
974	 => std_logic_vector(to_unsigned(96,8) ,
975	 => std_logic_vector(to_unsigned(95,8) ,
976	 => std_logic_vector(to_unsigned(95,8) ,
977	 => std_logic_vector(to_unsigned(97,8) ,
978	 => std_logic_vector(to_unsigned(91,8) ,
979	 => std_logic_vector(to_unsigned(81,8) ,
980	 => std_logic_vector(to_unsigned(86,8) ,
981	 => std_logic_vector(to_unsigned(92,8) ,
982	 => std_logic_vector(to_unsigned(96,8) ,
983	 => std_logic_vector(to_unsigned(96,8) ,
984	 => std_logic_vector(to_unsigned(99,8) ,
985	 => std_logic_vector(to_unsigned(104,8) ,
986	 => std_logic_vector(to_unsigned(105,8) ,
987	 => std_logic_vector(to_unsigned(100,8) ,
988	 => std_logic_vector(to_unsigned(103,8) ,
989	 => std_logic_vector(to_unsigned(101,8) ,
990	 => std_logic_vector(to_unsigned(100,8) ,
991	 => std_logic_vector(to_unsigned(104,8) ,
992	 => std_logic_vector(to_unsigned(107,8) ,
993	 => std_logic_vector(to_unsigned(104,8) ,
994	 => std_logic_vector(to_unsigned(104,8) ,
995	 => std_logic_vector(to_unsigned(103,8) ,
996	 => std_logic_vector(to_unsigned(104,8) ,
997	 => std_logic_vector(to_unsigned(103,8) ,
998	 => std_logic_vector(to_unsigned(103,8) ,
999	 => std_logic_vector(to_unsigned(101,8) ,
1000	 => std_logic_vector(to_unsigned(103,8) ,
1001	 => std_logic_vector(to_unsigned(108,8) ,
1002	 => std_logic_vector(to_unsigned(108,8) ,
1003	 => std_logic_vector(to_unsigned(109,8) ,
1004	 => std_logic_vector(to_unsigned(111,8) ,
1005	 => std_logic_vector(to_unsigned(109,8) ,
1006	 => std_logic_vector(to_unsigned(105,8) ,
1007	 => std_logic_vector(to_unsigned(108,8) ,
1008	 => std_logic_vector(to_unsigned(109,8) ,
1009	 => std_logic_vector(to_unsigned(114,8) ,
1010	 => std_logic_vector(to_unsigned(118,8) ,
1011	 => std_logic_vector(to_unsigned(115,8) ,
1012	 => std_logic_vector(to_unsigned(111,8) ,
1013	 => std_logic_vector(to_unsigned(112,8) ,
1014	 => std_logic_vector(to_unsigned(109,8) ,
1015	 => std_logic_vector(to_unsigned(103,8) ,
1016	 => std_logic_vector(to_unsigned(116,8) ,
1017	 => std_logic_vector(to_unsigned(118,8) ,
1018	 => std_logic_vector(to_unsigned(109,8) ,
1019	 => std_logic_vector(to_unsigned(107,8) ,
1020	 => std_logic_vector(to_unsigned(105,8) ,
1021	 => std_logic_vector(to_unsigned(108,8) ,
1022	 => std_logic_vector(to_unsigned(109,8) ,
1023	 => std_logic_vector(to_unsigned(108,8) ,
1024	 => std_logic_vector(to_unsigned(111,8) ,
1025	 => std_logic_vector(to_unsigned(115,8) ,
1026	 => std_logic_vector(to_unsigned(116,8) ,
1027	 => std_logic_vector(to_unsigned(112,8) ,
1028	 => std_logic_vector(to_unsigned(112,8) ,
1029	 => std_logic_vector(to_unsigned(116,8) ,
1030	 => std_logic_vector(to_unsigned(116,8) ,
1031	 => std_logic_vector(to_unsigned(115,8) ,
1032	 => std_logic_vector(to_unsigned(116,8) ,
1033	 => std_logic_vector(to_unsigned(116,8) ,
1034	 => std_logic_vector(to_unsigned(118,8) ,
1035	 => std_logic_vector(to_unsigned(109,8) ,
1036	 => std_logic_vector(to_unsigned(109,8) ,
1037	 => std_logic_vector(to_unsigned(111,8) ,
1038	 => std_logic_vector(to_unsigned(112,8) ,
1039	 => std_logic_vector(to_unsigned(115,8) ,
1040	 => std_logic_vector(to_unsigned(111,8) ,
1041	 => std_logic_vector(to_unsigned(105,8) ,
1042	 => std_logic_vector(to_unsigned(104,8) ,
1043	 => std_logic_vector(to_unsigned(114,8) ,
1044	 => std_logic_vector(to_unsigned(111,8) ,
1045	 => std_logic_vector(to_unsigned(105,8) ,
1046	 => std_logic_vector(to_unsigned(112,8) ,
1047	 => std_logic_vector(to_unsigned(116,8) ,
1048	 => std_logic_vector(to_unsigned(114,8) ,
1049	 => std_logic_vector(to_unsigned(108,8) ,
1050	 => std_logic_vector(to_unsigned(109,8) ,
1051	 => std_logic_vector(to_unsigned(114,8) ,
1052	 => std_logic_vector(to_unsigned(111,8) ,
1053	 => std_logic_vector(to_unsigned(108,8) ,
1054	 => std_logic_vector(to_unsigned(105,8) ,
1055	 => std_logic_vector(to_unsigned(105,8) ,
1056	 => std_logic_vector(to_unsigned(99,8) ,
1057	 => std_logic_vector(to_unsigned(95,8) ,
1058	 => std_logic_vector(to_unsigned(97,8) ,
1059	 => std_logic_vector(to_unsigned(101,8) ,
1060	 => std_logic_vector(to_unsigned(100,8) ,
1061	 => std_logic_vector(to_unsigned(100,8) ,
1062	 => std_logic_vector(to_unsigned(103,8) ,
1063	 => std_logic_vector(to_unsigned(100,8) ,
1064	 => std_logic_vector(to_unsigned(100,8) ,
1065	 => std_logic_vector(to_unsigned(103,8) ,
1066	 => std_logic_vector(to_unsigned(104,8) ,
1067	 => std_logic_vector(to_unsigned(112,8) ,
1068	 => std_logic_vector(to_unsigned(114,8) ,
1069	 => std_logic_vector(to_unsigned(111,8) ,
1070	 => std_logic_vector(to_unsigned(108,8) ,
1071	 => std_logic_vector(to_unsigned(107,8) ,
1072	 => std_logic_vector(to_unsigned(111,8) ,
1073	 => std_logic_vector(to_unsigned(108,8) ,
1074	 => std_logic_vector(to_unsigned(107,8) ,
1075	 => std_logic_vector(to_unsigned(109,8) ,
1076	 => std_logic_vector(to_unsigned(107,8) ,
1077	 => std_logic_vector(to_unsigned(108,8) ,
1078	 => std_logic_vector(to_unsigned(105,8) ,
1079	 => std_logic_vector(to_unsigned(107,8) ,
1080	 => std_logic_vector(to_unsigned(107,8) ,
1081	 => std_logic_vector(to_unsigned(105,8) ,
1082	 => std_logic_vector(to_unsigned(100,8) ,
1083	 => std_logic_vector(to_unsigned(101,8) ,
1084	 => std_logic_vector(to_unsigned(104,8) ,
1085	 => std_logic_vector(to_unsigned(107,8) ,
1086	 => std_logic_vector(to_unsigned(105,8) ,
1087	 => std_logic_vector(to_unsigned(103,8) ,
1088	 => std_logic_vector(to_unsigned(100,8) ,
1089	 => std_logic_vector(to_unsigned(101,8) ,
1090	 => std_logic_vector(to_unsigned(100,8) ,
1091	 => std_logic_vector(to_unsigned(100,8) ,
1092	 => std_logic_vector(to_unsigned(97,8) ,
1093	 => std_logic_vector(to_unsigned(97,8) ,
1094	 => std_logic_vector(to_unsigned(101,8) ,
1095	 => std_logic_vector(to_unsigned(100,8) ,
1096	 => std_logic_vector(to_unsigned(95,8) ,
1097	 => std_logic_vector(to_unsigned(96,8) ,
1098	 => std_logic_vector(to_unsigned(99,8) ,
1099	 => std_logic_vector(to_unsigned(97,8) ,
1100	 => std_logic_vector(to_unsigned(93,8) ,
1101	 => std_logic_vector(to_unsigned(103,8) ,
1102	 => std_logic_vector(to_unsigned(104,8) ,
1103	 => std_logic_vector(to_unsigned(99,8) ,
1104	 => std_logic_vector(to_unsigned(100,8) ,
1105	 => std_logic_vector(to_unsigned(103,8) ,
1106	 => std_logic_vector(to_unsigned(99,8) ,
1107	 => std_logic_vector(to_unsigned(101,8) ,
1108	 => std_logic_vector(to_unsigned(105,8) ,
1109	 => std_logic_vector(to_unsigned(105,8) ,
1110	 => std_logic_vector(to_unsigned(104,8) ,
1111	 => std_logic_vector(to_unsigned(100,8) ,
1112	 => std_logic_vector(to_unsigned(97,8) ,
1113	 => std_logic_vector(to_unsigned(96,8) ,
1114	 => std_logic_vector(to_unsigned(95,8) ,
1115	 => std_logic_vector(to_unsigned(90,8) ,
1116	 => std_logic_vector(to_unsigned(95,8) ,
1117	 => std_logic_vector(to_unsigned(95,8) ,
1118	 => std_logic_vector(to_unsigned(91,8) ,
1119	 => std_logic_vector(to_unsigned(92,8) ,
1120	 => std_logic_vector(to_unsigned(88,8) ,
1121	 => std_logic_vector(to_unsigned(88,8) ,
1122	 => std_logic_vector(to_unsigned(93,8) ,
1123	 => std_logic_vector(to_unsigned(95,8) ,
1124	 => std_logic_vector(to_unsigned(88,8) ,
1125	 => std_logic_vector(to_unsigned(90,8) ,
1126	 => std_logic_vector(to_unsigned(91,8) ,
1127	 => std_logic_vector(to_unsigned(85,8) ,
1128	 => std_logic_vector(to_unsigned(84,8) ,
1129	 => std_logic_vector(to_unsigned(90,8) ,
1130	 => std_logic_vector(to_unsigned(95,8) ,
1131	 => std_logic_vector(to_unsigned(90,8) ,
1132	 => std_logic_vector(to_unsigned(86,8) ,
1133	 => std_logic_vector(to_unsigned(92,8) ,
1134	 => std_logic_vector(to_unsigned(95,8) ,
1135	 => std_logic_vector(to_unsigned(91,8) ,
1136	 => std_logic_vector(to_unsigned(87,8) ,
1137	 => std_logic_vector(to_unsigned(87,8) ,
1138	 => std_logic_vector(to_unsigned(84,8) ,
1139	 => std_logic_vector(to_unsigned(86,8) ,
1140	 => std_logic_vector(to_unsigned(92,8) ,
1141	 => std_logic_vector(to_unsigned(88,8) ,
1142	 => std_logic_vector(to_unsigned(86,8) ,
1143	 => std_logic_vector(to_unsigned(86,8) ,
1144	 => std_logic_vector(to_unsigned(88,8) ,
1145	 => std_logic_vector(to_unsigned(91,8) ,
1146	 => std_logic_vector(to_unsigned(90,8) ,
1147	 => std_logic_vector(to_unsigned(82,8) ,
1148	 => std_logic_vector(to_unsigned(81,8) ,
1149	 => std_logic_vector(to_unsigned(88,8) ,
1150	 => std_logic_vector(to_unsigned(87,8) ,
1151	 => std_logic_vector(to_unsigned(88,8) ,
1152	 => std_logic_vector(to_unsigned(80,8) ,
1153	 => std_logic_vector(to_unsigned(84,8) ,
1154	 => std_logic_vector(to_unsigned(86,8) ,
1155	 => std_logic_vector(to_unsigned(85,8) ,
1156	 => std_logic_vector(to_unsigned(86,8) ,
1157	 => std_logic_vector(to_unsigned(85,8) ,
1158	 => std_logic_vector(to_unsigned(92,8) ,
1159	 => std_logic_vector(to_unsigned(92,8) ,
1160	 => std_logic_vector(to_unsigned(90,8) ,
1161	 => std_logic_vector(to_unsigned(88,8) ,
1162	 => std_logic_vector(to_unsigned(90,8) ,
1163	 => std_logic_vector(to_unsigned(91,8) ,
1164	 => std_logic_vector(to_unsigned(87,8) ,
1165	 => std_logic_vector(to_unsigned(87,8) ,
1166	 => std_logic_vector(to_unsigned(87,8) ,
1167	 => std_logic_vector(to_unsigned(85,8) ,
1168	 => std_logic_vector(to_unsigned(90,8) ,
1169	 => std_logic_vector(to_unsigned(88,8) ,
1170	 => std_logic_vector(to_unsigned(84,8) ,
1171	 => std_logic_vector(to_unsigned(86,8) ,
1172	 => std_logic_vector(to_unsigned(95,8) ,
1173	 => std_logic_vector(to_unsigned(91,8) ,
1174	 => std_logic_vector(to_unsigned(90,8) ,
1175	 => std_logic_vector(to_unsigned(91,8) ,
1176	 => std_logic_vector(to_unsigned(95,8) ,
1177	 => std_logic_vector(to_unsigned(90,8) ,
1178	 => std_logic_vector(to_unsigned(92,8) ,
1179	 => std_logic_vector(to_unsigned(96,8) ,
1180	 => std_logic_vector(to_unsigned(92,8) ,
1181	 => std_logic_vector(to_unsigned(91,8) ,
1182	 => std_logic_vector(to_unsigned(92,8) ,
1183	 => std_logic_vector(to_unsigned(90,8) ,
1184	 => std_logic_vector(to_unsigned(93,8) ,
1185	 => std_logic_vector(to_unsigned(100,8) ,
1186	 => std_logic_vector(to_unsigned(96,8) ,
1187	 => std_logic_vector(to_unsigned(92,8) ,
1188	 => std_logic_vector(to_unsigned(96,8) ,
1189	 => std_logic_vector(to_unsigned(96,8) ,
1190	 => std_logic_vector(to_unsigned(99,8) ,
1191	 => std_logic_vector(to_unsigned(97,8) ,
1192	 => std_logic_vector(to_unsigned(91,8) ,
1193	 => std_logic_vector(to_unsigned(81,8) ,
1194	 => std_logic_vector(to_unsigned(87,8) ,
1195	 => std_logic_vector(to_unsigned(68,8) ,
1196	 => std_logic_vector(to_unsigned(4,8) ,
1197	 => std_logic_vector(to_unsigned(0,8) ,
1198	 => std_logic_vector(to_unsigned(0,8) ,
1199	 => std_logic_vector(to_unsigned(23,8) ,
1200	 => std_logic_vector(to_unsigned(100,8) ,
1201	 => std_logic_vector(to_unsigned(88,8) ,
1202	 => std_logic_vector(to_unsigned(92,8) ,
1203	 => std_logic_vector(to_unsigned(91,8) ,
1204	 => std_logic_vector(to_unsigned(84,8) ,
1205	 => std_logic_vector(to_unsigned(92,8) ,
1206	 => std_logic_vector(to_unsigned(105,8) ,
1207	 => std_logic_vector(to_unsigned(111,8) ,
1208	 => std_logic_vector(to_unsigned(104,8) ,
1209	 => std_logic_vector(to_unsigned(104,8) ,
1210	 => std_logic_vector(to_unsigned(108,8) ,
1211	 => std_logic_vector(to_unsigned(114,8) ,
1212	 => std_logic_vector(to_unsigned(115,8) ,
1213	 => std_logic_vector(to_unsigned(115,8) ,
1214	 => std_logic_vector(to_unsigned(111,8) ,
1215	 => std_logic_vector(to_unsigned(114,8) ,
1216	 => std_logic_vector(to_unsigned(116,8) ,
1217	 => std_logic_vector(to_unsigned(109,8) ,
1218	 => std_logic_vector(to_unsigned(109,8) ,
1219	 => std_logic_vector(to_unsigned(112,8) ,
1220	 => std_logic_vector(to_unsigned(112,8) ,
1221	 => std_logic_vector(to_unsigned(111,8) ,
1222	 => std_logic_vector(to_unsigned(109,8) ,
1223	 => std_logic_vector(to_unsigned(111,8) ,
1224	 => std_logic_vector(to_unsigned(116,8) ,
1225	 => std_logic_vector(to_unsigned(115,8) ,
1226	 => std_logic_vector(to_unsigned(114,8) ,
1227	 => std_logic_vector(to_unsigned(115,8) ,
1228	 => std_logic_vector(to_unsigned(112,8) ,
1229	 => std_logic_vector(to_unsigned(112,8) ,
1230	 => std_logic_vector(to_unsigned(114,8) ,
1231	 => std_logic_vector(to_unsigned(118,8) ,
1232	 => std_logic_vector(to_unsigned(116,8) ,
1233	 => std_logic_vector(to_unsigned(121,8) ,
1234	 => std_logic_vector(to_unsigned(125,8) ,
1235	 => std_logic_vector(to_unsigned(130,8) ,
1236	 => std_logic_vector(to_unsigned(133,8) ,
1237	 => std_logic_vector(to_unsigned(134,8) ,
1238	 => std_logic_vector(to_unsigned(138,8) ,
1239	 => std_logic_vector(to_unsigned(146,8) ,
1240	 => std_logic_vector(to_unsigned(139,8) ,
1241	 => std_logic_vector(to_unsigned(141,8) ,
1242	 => std_logic_vector(to_unsigned(146,8) ,
1243	 => std_logic_vector(to_unsigned(144,8) ,
1244	 => std_logic_vector(to_unsigned(147,8) ,
1245	 => std_logic_vector(to_unsigned(149,8) ,
1246	 => std_logic_vector(to_unsigned(146,8) ,
1247	 => std_logic_vector(to_unsigned(142,8) ,
1248	 => std_logic_vector(to_unsigned(149,8) ,
1249	 => std_logic_vector(to_unsigned(152,8) ,
1250	 => std_logic_vector(to_unsigned(151,8) ,
1251	 => std_logic_vector(to_unsigned(151,8) ,
1252	 => std_logic_vector(to_unsigned(151,8) ,
1253	 => std_logic_vector(to_unsigned(152,8) ,
1254	 => std_logic_vector(to_unsigned(156,8) ,
1255	 => std_logic_vector(to_unsigned(161,8) ,
1256	 => std_logic_vector(to_unsigned(159,8) ,
1257	 => std_logic_vector(to_unsigned(157,8) ,
1258	 => std_logic_vector(to_unsigned(157,8) ,
1259	 => std_logic_vector(to_unsigned(159,8) ,
1260	 => std_logic_vector(to_unsigned(159,8) ,
1261	 => std_logic_vector(to_unsigned(161,8) ,
1262	 => std_logic_vector(to_unsigned(159,8) ,
1263	 => std_logic_vector(to_unsigned(159,8) ,
1264	 => std_logic_vector(to_unsigned(161,8) ,
1265	 => std_logic_vector(to_unsigned(166,8) ,
1266	 => std_logic_vector(to_unsigned(166,8) ,
1267	 => std_logic_vector(to_unsigned(164,8) ,
1268	 => std_logic_vector(to_unsigned(166,8) ,
1269	 => std_logic_vector(to_unsigned(164,8) ,
1270	 => std_logic_vector(to_unsigned(161,8) ,
1271	 => std_logic_vector(to_unsigned(161,8) ,
1272	 => std_logic_vector(to_unsigned(159,8) ,
1273	 => std_logic_vector(to_unsigned(161,8) ,
1274	 => std_logic_vector(to_unsigned(163,8) ,
1275	 => std_logic_vector(to_unsigned(161,8) ,
1276	 => std_logic_vector(to_unsigned(163,8) ,
1277	 => std_logic_vector(to_unsigned(166,8) ,
1278	 => std_logic_vector(to_unsigned(166,8) ,
1279	 => std_logic_vector(to_unsigned(164,8) ,
1280	 => std_logic_vector(to_unsigned(164,8) ,
1281	 => std_logic_vector(to_unsigned(103,8) ,
1282	 => std_logic_vector(to_unsigned(104,8) ,
1283	 => std_logic_vector(to_unsigned(104,8) ,
1284	 => std_logic_vector(to_unsigned(103,8) ,
1285	 => std_logic_vector(to_unsigned(105,8) ,
1286	 => std_logic_vector(to_unsigned(103,8) ,
1287	 => std_logic_vector(to_unsigned(101,8) ,
1288	 => std_logic_vector(to_unsigned(104,8) ,
1289	 => std_logic_vector(to_unsigned(101,8) ,
1290	 => std_logic_vector(to_unsigned(100,8) ,
1291	 => std_logic_vector(to_unsigned(101,8) ,
1292	 => std_logic_vector(to_unsigned(95,8) ,
1293	 => std_logic_vector(to_unsigned(91,8) ,
1294	 => std_logic_vector(to_unsigned(95,8) ,
1295	 => std_logic_vector(to_unsigned(95,8) ,
1296	 => std_logic_vector(to_unsigned(88,8) ,
1297	 => std_logic_vector(to_unsigned(90,8) ,
1298	 => std_logic_vector(to_unsigned(88,8) ,
1299	 => std_logic_vector(to_unsigned(85,8) ,
1300	 => std_logic_vector(to_unsigned(86,8) ,
1301	 => std_logic_vector(to_unsigned(86,8) ,
1302	 => std_logic_vector(to_unsigned(90,8) ,
1303	 => std_logic_vector(to_unsigned(95,8) ,
1304	 => std_logic_vector(to_unsigned(92,8) ,
1305	 => std_logic_vector(to_unsigned(93,8) ,
1306	 => std_logic_vector(to_unsigned(91,8) ,
1307	 => std_logic_vector(to_unsigned(92,8) ,
1308	 => std_logic_vector(to_unsigned(103,8) ,
1309	 => std_logic_vector(to_unsigned(99,8) ,
1310	 => std_logic_vector(to_unsigned(99,8) ,
1311	 => std_logic_vector(to_unsigned(103,8) ,
1312	 => std_logic_vector(to_unsigned(105,8) ,
1313	 => std_logic_vector(to_unsigned(100,8) ,
1314	 => std_logic_vector(to_unsigned(99,8) ,
1315	 => std_logic_vector(to_unsigned(100,8) ,
1316	 => std_logic_vector(to_unsigned(104,8) ,
1317	 => std_logic_vector(to_unsigned(104,8) ,
1318	 => std_logic_vector(to_unsigned(100,8) ,
1319	 => std_logic_vector(to_unsigned(101,8) ,
1320	 => std_logic_vector(to_unsigned(103,8) ,
1321	 => std_logic_vector(to_unsigned(105,8) ,
1322	 => std_logic_vector(to_unsigned(99,8) ,
1323	 => std_logic_vector(to_unsigned(99,8) ,
1324	 => std_logic_vector(to_unsigned(103,8) ,
1325	 => std_logic_vector(to_unsigned(107,8) ,
1326	 => std_logic_vector(to_unsigned(107,8) ,
1327	 => std_logic_vector(to_unsigned(109,8) ,
1328	 => std_logic_vector(to_unsigned(109,8) ,
1329	 => std_logic_vector(to_unsigned(111,8) ,
1330	 => std_logic_vector(to_unsigned(115,8) ,
1331	 => std_logic_vector(to_unsigned(109,8) ,
1332	 => std_logic_vector(to_unsigned(112,8) ,
1333	 => std_logic_vector(to_unsigned(109,8) ,
1334	 => std_logic_vector(to_unsigned(109,8) ,
1335	 => std_logic_vector(to_unsigned(111,8) ,
1336	 => std_logic_vector(to_unsigned(118,8) ,
1337	 => std_logic_vector(to_unsigned(116,8) ,
1338	 => std_logic_vector(to_unsigned(115,8) ,
1339	 => std_logic_vector(to_unsigned(112,8) ,
1340	 => std_logic_vector(to_unsigned(108,8) ,
1341	 => std_logic_vector(to_unsigned(109,8) ,
1342	 => std_logic_vector(to_unsigned(111,8) ,
1343	 => std_logic_vector(to_unsigned(114,8) ,
1344	 => std_logic_vector(to_unsigned(116,8) ,
1345	 => std_logic_vector(to_unsigned(115,8) ,
1346	 => std_logic_vector(to_unsigned(115,8) ,
1347	 => std_logic_vector(to_unsigned(114,8) ,
1348	 => std_logic_vector(to_unsigned(111,8) ,
1349	 => std_logic_vector(to_unsigned(109,8) ,
1350	 => std_logic_vector(to_unsigned(115,8) ,
1351	 => std_logic_vector(to_unsigned(111,8) ,
1352	 => std_logic_vector(to_unsigned(109,8) ,
1353	 => std_logic_vector(to_unsigned(111,8) ,
1354	 => std_logic_vector(to_unsigned(116,8) ,
1355	 => std_logic_vector(to_unsigned(112,8) ,
1356	 => std_logic_vector(to_unsigned(109,8) ,
1357	 => std_logic_vector(to_unsigned(108,8) ,
1358	 => std_logic_vector(to_unsigned(107,8) ,
1359	 => std_logic_vector(to_unsigned(107,8) ,
1360	 => std_logic_vector(to_unsigned(105,8) ,
1361	 => std_logic_vector(to_unsigned(107,8) ,
1362	 => std_logic_vector(to_unsigned(112,8) ,
1363	 => std_logic_vector(to_unsigned(115,8) ,
1364	 => std_logic_vector(to_unsigned(111,8) ,
1365	 => std_logic_vector(to_unsigned(111,8) ,
1366	 => std_logic_vector(to_unsigned(112,8) ,
1367	 => std_logic_vector(to_unsigned(107,8) ,
1368	 => std_logic_vector(to_unsigned(112,8) ,
1369	 => std_logic_vector(to_unsigned(112,8) ,
1370	 => std_logic_vector(to_unsigned(111,8) ,
1371	 => std_logic_vector(to_unsigned(111,8) ,
1372	 => std_logic_vector(to_unsigned(108,8) ,
1373	 => std_logic_vector(to_unsigned(107,8) ,
1374	 => std_logic_vector(to_unsigned(104,8) ,
1375	 => std_logic_vector(to_unsigned(105,8) ,
1376	 => std_logic_vector(to_unsigned(103,8) ,
1377	 => std_logic_vector(to_unsigned(93,8) ,
1378	 => std_logic_vector(to_unsigned(93,8) ,
1379	 => std_logic_vector(to_unsigned(96,8) ,
1380	 => std_logic_vector(to_unsigned(100,8) ,
1381	 => std_logic_vector(to_unsigned(104,8) ,
1382	 => std_logic_vector(to_unsigned(101,8) ,
1383	 => std_logic_vector(to_unsigned(97,8) ,
1384	 => std_logic_vector(to_unsigned(99,8) ,
1385	 => std_logic_vector(to_unsigned(104,8) ,
1386	 => std_logic_vector(to_unsigned(104,8) ,
1387	 => std_logic_vector(to_unsigned(104,8) ,
1388	 => std_logic_vector(to_unsigned(104,8) ,
1389	 => std_logic_vector(to_unsigned(108,8) ,
1390	 => std_logic_vector(to_unsigned(108,8) ,
1391	 => std_logic_vector(to_unsigned(104,8) ,
1392	 => std_logic_vector(to_unsigned(105,8) ,
1393	 => std_logic_vector(to_unsigned(104,8) ,
1394	 => std_logic_vector(to_unsigned(107,8) ,
1395	 => std_logic_vector(to_unsigned(111,8) ,
1396	 => std_logic_vector(to_unsigned(105,8) ,
1397	 => std_logic_vector(to_unsigned(105,8) ,
1398	 => std_logic_vector(to_unsigned(107,8) ,
1399	 => std_logic_vector(to_unsigned(104,8) ,
1400	 => std_logic_vector(to_unsigned(104,8) ,
1401	 => std_logic_vector(to_unsigned(104,8) ,
1402	 => std_logic_vector(to_unsigned(100,8) ,
1403	 => std_logic_vector(to_unsigned(97,8) ,
1404	 => std_logic_vector(to_unsigned(99,8) ,
1405	 => std_logic_vector(to_unsigned(100,8) ,
1406	 => std_logic_vector(to_unsigned(99,8) ,
1407	 => std_logic_vector(to_unsigned(100,8) ,
1408	 => std_logic_vector(to_unsigned(97,8) ,
1409	 => std_logic_vector(to_unsigned(95,8) ,
1410	 => std_logic_vector(to_unsigned(96,8) ,
1411	 => std_logic_vector(to_unsigned(99,8) ,
1412	 => std_logic_vector(to_unsigned(96,8) ,
1413	 => std_logic_vector(to_unsigned(96,8) ,
1414	 => std_logic_vector(to_unsigned(104,8) ,
1415	 => std_logic_vector(to_unsigned(104,8) ,
1416	 => std_logic_vector(to_unsigned(99,8) ,
1417	 => std_logic_vector(to_unsigned(100,8) ,
1418	 => std_logic_vector(to_unsigned(103,8) ,
1419	 => std_logic_vector(to_unsigned(99,8) ,
1420	 => std_logic_vector(to_unsigned(100,8) ,
1421	 => std_logic_vector(to_unsigned(103,8) ,
1422	 => std_logic_vector(to_unsigned(101,8) ,
1423	 => std_logic_vector(to_unsigned(97,8) ,
1424	 => std_logic_vector(to_unsigned(97,8) ,
1425	 => std_logic_vector(to_unsigned(104,8) ,
1426	 => std_logic_vector(to_unsigned(100,8) ,
1427	 => std_logic_vector(to_unsigned(103,8) ,
1428	 => std_logic_vector(to_unsigned(107,8) ,
1429	 => std_logic_vector(to_unsigned(105,8) ,
1430	 => std_logic_vector(to_unsigned(101,8) ,
1431	 => std_logic_vector(to_unsigned(103,8) ,
1432	 => std_logic_vector(to_unsigned(101,8) ,
1433	 => std_logic_vector(to_unsigned(97,8) ,
1434	 => std_logic_vector(to_unsigned(92,8) ,
1435	 => std_logic_vector(to_unsigned(90,8) ,
1436	 => std_logic_vector(to_unsigned(96,8) ,
1437	 => std_logic_vector(to_unsigned(92,8) ,
1438	 => std_logic_vector(to_unsigned(86,8) ,
1439	 => std_logic_vector(to_unsigned(88,8) ,
1440	 => std_logic_vector(to_unsigned(86,8) ,
1441	 => std_logic_vector(to_unsigned(85,8) ,
1442	 => std_logic_vector(to_unsigned(91,8) ,
1443	 => std_logic_vector(to_unsigned(96,8) ,
1444	 => std_logic_vector(to_unsigned(90,8) ,
1445	 => std_logic_vector(to_unsigned(88,8) ,
1446	 => std_logic_vector(to_unsigned(91,8) ,
1447	 => std_logic_vector(to_unsigned(90,8) ,
1448	 => std_logic_vector(to_unsigned(90,8) ,
1449	 => std_logic_vector(to_unsigned(88,8) ,
1450	 => std_logic_vector(to_unsigned(93,8) ,
1451	 => std_logic_vector(to_unsigned(90,8) ,
1452	 => std_logic_vector(to_unsigned(86,8) ,
1453	 => std_logic_vector(to_unsigned(95,8) ,
1454	 => std_logic_vector(to_unsigned(90,8) ,
1455	 => std_logic_vector(to_unsigned(88,8) ,
1456	 => std_logic_vector(to_unsigned(86,8) ,
1457	 => std_logic_vector(to_unsigned(87,8) ,
1458	 => std_logic_vector(to_unsigned(88,8) ,
1459	 => std_logic_vector(to_unsigned(88,8) ,
1460	 => std_logic_vector(to_unsigned(90,8) ,
1461	 => std_logic_vector(to_unsigned(86,8) ,
1462	 => std_logic_vector(to_unsigned(85,8) ,
1463	 => std_logic_vector(to_unsigned(86,8) ,
1464	 => std_logic_vector(to_unsigned(88,8) ,
1465	 => std_logic_vector(to_unsigned(90,8) ,
1466	 => std_logic_vector(to_unsigned(86,8) ,
1467	 => std_logic_vector(to_unsigned(78,8) ,
1468	 => std_logic_vector(to_unsigned(82,8) ,
1469	 => std_logic_vector(to_unsigned(87,8) ,
1470	 => std_logic_vector(to_unsigned(84,8) ,
1471	 => std_logic_vector(to_unsigned(85,8) ,
1472	 => std_logic_vector(to_unsigned(80,8) ,
1473	 => std_logic_vector(to_unsigned(84,8) ,
1474	 => std_logic_vector(to_unsigned(86,8) ,
1475	 => std_logic_vector(to_unsigned(86,8) ,
1476	 => std_logic_vector(to_unsigned(85,8) ,
1477	 => std_logic_vector(to_unsigned(86,8) ,
1478	 => std_logic_vector(to_unsigned(92,8) ,
1479	 => std_logic_vector(to_unsigned(91,8) ,
1480	 => std_logic_vector(to_unsigned(86,8) ,
1481	 => std_logic_vector(to_unsigned(84,8) ,
1482	 => std_logic_vector(to_unsigned(85,8) ,
1483	 => std_logic_vector(to_unsigned(87,8) ,
1484	 => std_logic_vector(to_unsigned(86,8) ,
1485	 => std_logic_vector(to_unsigned(87,8) ,
1486	 => std_logic_vector(to_unsigned(88,8) ,
1487	 => std_logic_vector(to_unsigned(91,8) ,
1488	 => std_logic_vector(to_unsigned(87,8) ,
1489	 => std_logic_vector(to_unsigned(85,8) ,
1490	 => std_logic_vector(to_unsigned(86,8) ,
1491	 => std_logic_vector(to_unsigned(90,8) ,
1492	 => std_logic_vector(to_unsigned(93,8) ,
1493	 => std_logic_vector(to_unsigned(88,8) ,
1494	 => std_logic_vector(to_unsigned(90,8) ,
1495	 => std_logic_vector(to_unsigned(90,8) ,
1496	 => std_logic_vector(to_unsigned(91,8) ,
1497	 => std_logic_vector(to_unsigned(90,8) ,
1498	 => std_logic_vector(to_unsigned(88,8) ,
1499	 => std_logic_vector(to_unsigned(93,8) ,
1500	 => std_logic_vector(to_unsigned(91,8) ,
1501	 => std_logic_vector(to_unsigned(85,8) ,
1502	 => std_logic_vector(to_unsigned(88,8) ,
1503	 => std_logic_vector(to_unsigned(88,8) ,
1504	 => std_logic_vector(to_unsigned(95,8) ,
1505	 => std_logic_vector(to_unsigned(99,8) ,
1506	 => std_logic_vector(to_unsigned(91,8) ,
1507	 => std_logic_vector(to_unsigned(90,8) ,
1508	 => std_logic_vector(to_unsigned(95,8) ,
1509	 => std_logic_vector(to_unsigned(93,8) ,
1510	 => std_logic_vector(to_unsigned(95,8) ,
1511	 => std_logic_vector(to_unsigned(93,8) ,
1512	 => std_logic_vector(to_unsigned(86,8) ,
1513	 => std_logic_vector(to_unsigned(76,8) ,
1514	 => std_logic_vector(to_unsigned(80,8) ,
1515	 => std_logic_vector(to_unsigned(85,8) ,
1516	 => std_logic_vector(to_unsigned(13,8) ,
1517	 => std_logic_vector(to_unsigned(0,8) ,
1518	 => std_logic_vector(to_unsigned(0,8) ,
1519	 => std_logic_vector(to_unsigned(7,8) ,
1520	 => std_logic_vector(to_unsigned(87,8) ,
1521	 => std_logic_vector(to_unsigned(93,8) ,
1522	 => std_logic_vector(to_unsigned(88,8) ,
1523	 => std_logic_vector(to_unsigned(90,8) ,
1524	 => std_logic_vector(to_unsigned(92,8) ,
1525	 => std_logic_vector(to_unsigned(99,8) ,
1526	 => std_logic_vector(to_unsigned(108,8) ,
1527	 => std_logic_vector(to_unsigned(109,8) ,
1528	 => std_logic_vector(to_unsigned(108,8) ,
1529	 => std_logic_vector(to_unsigned(111,8) ,
1530	 => std_logic_vector(to_unsigned(112,8) ,
1531	 => std_logic_vector(to_unsigned(111,8) ,
1532	 => std_logic_vector(to_unsigned(112,8) ,
1533	 => std_logic_vector(to_unsigned(115,8) ,
1534	 => std_logic_vector(to_unsigned(114,8) ,
1535	 => std_logic_vector(to_unsigned(116,8) ,
1536	 => std_logic_vector(to_unsigned(112,8) ,
1537	 => std_logic_vector(to_unsigned(107,8) ,
1538	 => std_logic_vector(to_unsigned(108,8) ,
1539	 => std_logic_vector(to_unsigned(116,8) ,
1540	 => std_logic_vector(to_unsigned(119,8) ,
1541	 => std_logic_vector(to_unsigned(112,8) ,
1542	 => std_logic_vector(to_unsigned(107,8) ,
1543	 => std_logic_vector(to_unsigned(109,8) ,
1544	 => std_logic_vector(to_unsigned(115,8) ,
1545	 => std_logic_vector(to_unsigned(114,8) ,
1546	 => std_logic_vector(to_unsigned(111,8) ,
1547	 => std_logic_vector(to_unsigned(109,8) ,
1548	 => std_logic_vector(to_unsigned(108,8) ,
1549	 => std_logic_vector(to_unsigned(111,8) ,
1550	 => std_logic_vector(to_unsigned(114,8) ,
1551	 => std_logic_vector(to_unsigned(114,8) ,
1552	 => std_logic_vector(to_unsigned(114,8) ,
1553	 => std_logic_vector(to_unsigned(115,8) ,
1554	 => std_logic_vector(to_unsigned(122,8) ,
1555	 => std_logic_vector(to_unsigned(131,8) ,
1556	 => std_logic_vector(to_unsigned(138,8) ,
1557	 => std_logic_vector(to_unsigned(138,8) ,
1558	 => std_logic_vector(to_unsigned(133,8) ,
1559	 => std_logic_vector(to_unsigned(139,8) ,
1560	 => std_logic_vector(to_unsigned(139,8) ,
1561	 => std_logic_vector(to_unsigned(144,8) ,
1562	 => std_logic_vector(to_unsigned(147,8) ,
1563	 => std_logic_vector(to_unsigned(144,8) ,
1564	 => std_logic_vector(to_unsigned(144,8) ,
1565	 => std_logic_vector(to_unsigned(144,8) ,
1566	 => std_logic_vector(to_unsigned(149,8) ,
1567	 => std_logic_vector(to_unsigned(146,8) ,
1568	 => std_logic_vector(to_unsigned(144,8) ,
1569	 => std_logic_vector(to_unsigned(144,8) ,
1570	 => std_logic_vector(to_unsigned(146,8) ,
1571	 => std_logic_vector(to_unsigned(147,8) ,
1572	 => std_logic_vector(to_unsigned(151,8) ,
1573	 => std_logic_vector(to_unsigned(151,8) ,
1574	 => std_logic_vector(to_unsigned(151,8) ,
1575	 => std_logic_vector(to_unsigned(154,8) ,
1576	 => std_logic_vector(to_unsigned(157,8) ,
1577	 => std_logic_vector(to_unsigned(159,8) ,
1578	 => std_logic_vector(to_unsigned(159,8) ,
1579	 => std_logic_vector(to_unsigned(161,8) ,
1580	 => std_logic_vector(to_unsigned(161,8) ,
1581	 => std_logic_vector(to_unsigned(161,8) ,
1582	 => std_logic_vector(to_unsigned(159,8) ,
1583	 => std_logic_vector(to_unsigned(157,8) ,
1584	 => std_logic_vector(to_unsigned(159,8) ,
1585	 => std_logic_vector(to_unsigned(159,8) ,
1586	 => std_logic_vector(to_unsigned(157,8) ,
1587	 => std_logic_vector(to_unsigned(161,8) ,
1588	 => std_logic_vector(to_unsigned(163,8) ,
1589	 => std_logic_vector(to_unsigned(161,8) ,
1590	 => std_logic_vector(to_unsigned(161,8) ,
1591	 => std_logic_vector(to_unsigned(161,8) ,
1592	 => std_logic_vector(to_unsigned(161,8) ,
1593	 => std_logic_vector(to_unsigned(157,8) ,
1594	 => std_logic_vector(to_unsigned(161,8) ,
1595	 => std_logic_vector(to_unsigned(164,8) ,
1596	 => std_logic_vector(to_unsigned(164,8) ,
1597	 => std_logic_vector(to_unsigned(163,8) ,
1598	 => std_logic_vector(to_unsigned(161,8) ,
1599	 => std_logic_vector(to_unsigned(161,8) ,
1600	 => std_logic_vector(to_unsigned(163,8) ,
1601	 => std_logic_vector(to_unsigned(101,8) ,
1602	 => std_logic_vector(to_unsigned(96,8) ,
1603	 => std_logic_vector(to_unsigned(100,8) ,
1604	 => std_logic_vector(to_unsigned(99,8) ,
1605	 => std_logic_vector(to_unsigned(96,8) ,
1606	 => std_logic_vector(to_unsigned(97,8) ,
1607	 => std_logic_vector(to_unsigned(97,8) ,
1608	 => std_logic_vector(to_unsigned(100,8) ,
1609	 => std_logic_vector(to_unsigned(97,8) ,
1610	 => std_logic_vector(to_unsigned(95,8) ,
1611	 => std_logic_vector(to_unsigned(95,8) ,
1612	 => std_logic_vector(to_unsigned(93,8) ,
1613	 => std_logic_vector(to_unsigned(92,8) ,
1614	 => std_logic_vector(to_unsigned(95,8) ,
1615	 => std_logic_vector(to_unsigned(95,8) ,
1616	 => std_logic_vector(to_unsigned(92,8) ,
1617	 => std_logic_vector(to_unsigned(92,8) ,
1618	 => std_logic_vector(to_unsigned(88,8) ,
1619	 => std_logic_vector(to_unsigned(87,8) ,
1620	 => std_logic_vector(to_unsigned(86,8) ,
1621	 => std_logic_vector(to_unsigned(84,8) ,
1622	 => std_logic_vector(to_unsigned(91,8) ,
1623	 => std_logic_vector(to_unsigned(96,8) ,
1624	 => std_logic_vector(to_unsigned(93,8) ,
1625	 => std_logic_vector(to_unsigned(88,8) ,
1626	 => std_logic_vector(to_unsigned(88,8) ,
1627	 => std_logic_vector(to_unsigned(101,8) ,
1628	 => std_logic_vector(to_unsigned(101,8) ,
1629	 => std_logic_vector(to_unsigned(97,8) ,
1630	 => std_logic_vector(to_unsigned(101,8) ,
1631	 => std_logic_vector(to_unsigned(104,8) ,
1632	 => std_logic_vector(to_unsigned(104,8) ,
1633	 => std_logic_vector(to_unsigned(99,8) ,
1634	 => std_logic_vector(to_unsigned(95,8) ,
1635	 => std_logic_vector(to_unsigned(95,8) ,
1636	 => std_logic_vector(to_unsigned(100,8) ,
1637	 => std_logic_vector(to_unsigned(101,8) ,
1638	 => std_logic_vector(to_unsigned(96,8) ,
1639	 => std_logic_vector(to_unsigned(103,8) ,
1640	 => std_logic_vector(to_unsigned(104,8) ,
1641	 => std_logic_vector(to_unsigned(104,8) ,
1642	 => std_logic_vector(to_unsigned(100,8) ,
1643	 => std_logic_vector(to_unsigned(101,8) ,
1644	 => std_logic_vector(to_unsigned(101,8) ,
1645	 => std_logic_vector(to_unsigned(104,8) ,
1646	 => std_logic_vector(to_unsigned(109,8) ,
1647	 => std_logic_vector(to_unsigned(114,8) ,
1648	 => std_logic_vector(to_unsigned(109,8) ,
1649	 => std_logic_vector(to_unsigned(111,8) ,
1650	 => std_logic_vector(to_unsigned(115,8) ,
1651	 => std_logic_vector(to_unsigned(111,8) ,
1652	 => std_logic_vector(to_unsigned(108,8) ,
1653	 => std_logic_vector(to_unsigned(109,8) ,
1654	 => std_logic_vector(to_unsigned(109,8) ,
1655	 => std_logic_vector(to_unsigned(105,8) ,
1656	 => std_logic_vector(to_unsigned(107,8) ,
1657	 => std_logic_vector(to_unsigned(115,8) ,
1658	 => std_logic_vector(to_unsigned(115,8) ,
1659	 => std_logic_vector(to_unsigned(112,8) ,
1660	 => std_logic_vector(to_unsigned(109,8) ,
1661	 => std_logic_vector(to_unsigned(109,8) ,
1662	 => std_logic_vector(to_unsigned(108,8) ,
1663	 => std_logic_vector(to_unsigned(111,8) ,
1664	 => std_logic_vector(to_unsigned(114,8) ,
1665	 => std_logic_vector(to_unsigned(116,8) ,
1666	 => std_logic_vector(to_unsigned(114,8) ,
1667	 => std_logic_vector(to_unsigned(112,8) ,
1668	 => std_logic_vector(to_unsigned(108,8) ,
1669	 => std_logic_vector(to_unsigned(103,8) ,
1670	 => std_logic_vector(to_unsigned(114,8) ,
1671	 => std_logic_vector(to_unsigned(114,8) ,
1672	 => std_logic_vector(to_unsigned(111,8) ,
1673	 => std_logic_vector(to_unsigned(111,8) ,
1674	 => std_logic_vector(to_unsigned(116,8) ,
1675	 => std_logic_vector(to_unsigned(112,8) ,
1676	 => std_logic_vector(to_unsigned(111,8) ,
1677	 => std_logic_vector(to_unsigned(112,8) ,
1678	 => std_logic_vector(to_unsigned(109,8) ,
1679	 => std_logic_vector(to_unsigned(104,8) ,
1680	 => std_logic_vector(to_unsigned(107,8) ,
1681	 => std_logic_vector(to_unsigned(111,8) ,
1682	 => std_logic_vector(to_unsigned(112,8) ,
1683	 => std_logic_vector(to_unsigned(111,8) ,
1684	 => std_logic_vector(to_unsigned(112,8) ,
1685	 => std_logic_vector(to_unsigned(115,8) ,
1686	 => std_logic_vector(to_unsigned(112,8) ,
1687	 => std_logic_vector(to_unsigned(108,8) ,
1688	 => std_logic_vector(to_unsigned(109,8) ,
1689	 => std_logic_vector(to_unsigned(108,8) ,
1690	 => std_logic_vector(to_unsigned(109,8) ,
1691	 => std_logic_vector(to_unsigned(112,8) ,
1692	 => std_logic_vector(to_unsigned(109,8) ,
1693	 => std_logic_vector(to_unsigned(104,8) ,
1694	 => std_logic_vector(to_unsigned(100,8) ,
1695	 => std_logic_vector(to_unsigned(103,8) ,
1696	 => std_logic_vector(to_unsigned(101,8) ,
1697	 => std_logic_vector(to_unsigned(93,8) ,
1698	 => std_logic_vector(to_unsigned(99,8) ,
1699	 => std_logic_vector(to_unsigned(95,8) ,
1700	 => std_logic_vector(to_unsigned(99,8) ,
1701	 => std_logic_vector(to_unsigned(104,8) ,
1702	 => std_logic_vector(to_unsigned(101,8) ,
1703	 => std_logic_vector(to_unsigned(103,8) ,
1704	 => std_logic_vector(to_unsigned(101,8) ,
1705	 => std_logic_vector(to_unsigned(104,8) ,
1706	 => std_logic_vector(to_unsigned(111,8) ,
1707	 => std_logic_vector(to_unsigned(107,8) ,
1708	 => std_logic_vector(to_unsigned(109,8) ,
1709	 => std_logic_vector(to_unsigned(112,8) ,
1710	 => std_logic_vector(to_unsigned(108,8) ,
1711	 => std_logic_vector(to_unsigned(105,8) ,
1712	 => std_logic_vector(to_unsigned(107,8) ,
1713	 => std_logic_vector(to_unsigned(109,8) ,
1714	 => std_logic_vector(to_unsigned(108,8) ,
1715	 => std_logic_vector(to_unsigned(111,8) ,
1716	 => std_logic_vector(to_unsigned(105,8) ,
1717	 => std_logic_vector(to_unsigned(107,8) ,
1718	 => std_logic_vector(to_unsigned(108,8) ,
1719	 => std_logic_vector(to_unsigned(103,8) ,
1720	 => std_logic_vector(to_unsigned(100,8) ,
1721	 => std_logic_vector(to_unsigned(104,8) ,
1722	 => std_logic_vector(to_unsigned(96,8) ,
1723	 => std_logic_vector(to_unsigned(99,8) ,
1724	 => std_logic_vector(to_unsigned(105,8) ,
1725	 => std_logic_vector(to_unsigned(103,8) ,
1726	 => std_logic_vector(to_unsigned(96,8) ,
1727	 => std_logic_vector(to_unsigned(96,8) ,
1728	 => std_logic_vector(to_unsigned(96,8) ,
1729	 => std_logic_vector(to_unsigned(97,8) ,
1730	 => std_logic_vector(to_unsigned(96,8) ,
1731	 => std_logic_vector(to_unsigned(96,8) ,
1732	 => std_logic_vector(to_unsigned(99,8) ,
1733	 => std_logic_vector(to_unsigned(99,8) ,
1734	 => std_logic_vector(to_unsigned(101,8) ,
1735	 => std_logic_vector(to_unsigned(99,8) ,
1736	 => std_logic_vector(to_unsigned(97,8) ,
1737	 => std_logic_vector(to_unsigned(100,8) ,
1738	 => std_logic_vector(to_unsigned(100,8) ,
1739	 => std_logic_vector(to_unsigned(99,8) ,
1740	 => std_logic_vector(to_unsigned(103,8) ,
1741	 => std_logic_vector(to_unsigned(101,8) ,
1742	 => std_logic_vector(to_unsigned(101,8) ,
1743	 => std_logic_vector(to_unsigned(103,8) ,
1744	 => std_logic_vector(to_unsigned(101,8) ,
1745	 => std_logic_vector(to_unsigned(104,8) ,
1746	 => std_logic_vector(to_unsigned(103,8) ,
1747	 => std_logic_vector(to_unsigned(109,8) ,
1748	 => std_logic_vector(to_unsigned(108,8) ,
1749	 => std_logic_vector(to_unsigned(104,8) ,
1750	 => std_logic_vector(to_unsigned(101,8) ,
1751	 => std_logic_vector(to_unsigned(101,8) ,
1752	 => std_logic_vector(to_unsigned(99,8) ,
1753	 => std_logic_vector(to_unsigned(95,8) ,
1754	 => std_logic_vector(to_unsigned(95,8) ,
1755	 => std_logic_vector(to_unsigned(90,8) ,
1756	 => std_logic_vector(to_unsigned(84,8) ,
1757	 => std_logic_vector(to_unsigned(82,8) ,
1758	 => std_logic_vector(to_unsigned(84,8) ,
1759	 => std_logic_vector(to_unsigned(86,8) ,
1760	 => std_logic_vector(to_unsigned(85,8) ,
1761	 => std_logic_vector(to_unsigned(87,8) ,
1762	 => std_logic_vector(to_unsigned(88,8) ,
1763	 => std_logic_vector(to_unsigned(86,8) ,
1764	 => std_logic_vector(to_unsigned(88,8) ,
1765	 => std_logic_vector(to_unsigned(85,8) ,
1766	 => std_logic_vector(to_unsigned(87,8) ,
1767	 => std_logic_vector(to_unsigned(91,8) ,
1768	 => std_logic_vector(to_unsigned(88,8) ,
1769	 => std_logic_vector(to_unsigned(84,8) ,
1770	 => std_logic_vector(to_unsigned(86,8) ,
1771	 => std_logic_vector(to_unsigned(85,8) ,
1772	 => std_logic_vector(to_unsigned(90,8) ,
1773	 => std_logic_vector(to_unsigned(93,8) ,
1774	 => std_logic_vector(to_unsigned(82,8) ,
1775	 => std_logic_vector(to_unsigned(87,8) ,
1776	 => std_logic_vector(to_unsigned(90,8) ,
1777	 => std_logic_vector(to_unsigned(85,8) ,
1778	 => std_logic_vector(to_unsigned(88,8) ,
1779	 => std_logic_vector(to_unsigned(90,8) ,
1780	 => std_logic_vector(to_unsigned(88,8) ,
1781	 => std_logic_vector(to_unsigned(87,8) ,
1782	 => std_logic_vector(to_unsigned(81,8) ,
1783	 => std_logic_vector(to_unsigned(82,8) ,
1784	 => std_logic_vector(to_unsigned(85,8) ,
1785	 => std_logic_vector(to_unsigned(84,8) ,
1786	 => std_logic_vector(to_unsigned(85,8) ,
1787	 => std_logic_vector(to_unsigned(87,8) ,
1788	 => std_logic_vector(to_unsigned(90,8) ,
1789	 => std_logic_vector(to_unsigned(84,8) ,
1790	 => std_logic_vector(to_unsigned(82,8) ,
1791	 => std_logic_vector(to_unsigned(81,8) ,
1792	 => std_logic_vector(to_unsigned(81,8) ,
1793	 => std_logic_vector(to_unsigned(90,8) ,
1794	 => std_logic_vector(to_unsigned(90,8) ,
1795	 => std_logic_vector(to_unsigned(84,8) ,
1796	 => std_logic_vector(to_unsigned(80,8) ,
1797	 => std_logic_vector(to_unsigned(84,8) ,
1798	 => std_logic_vector(to_unsigned(82,8) ,
1799	 => std_logic_vector(to_unsigned(86,8) ,
1800	 => std_logic_vector(to_unsigned(88,8) ,
1801	 => std_logic_vector(to_unsigned(85,8) ,
1802	 => std_logic_vector(to_unsigned(87,8) ,
1803	 => std_logic_vector(to_unsigned(86,8) ,
1804	 => std_logic_vector(to_unsigned(85,8) ,
1805	 => std_logic_vector(to_unsigned(86,8) ,
1806	 => std_logic_vector(to_unsigned(88,8) ,
1807	 => std_logic_vector(to_unsigned(88,8) ,
1808	 => std_logic_vector(to_unsigned(86,8) ,
1809	 => std_logic_vector(to_unsigned(84,8) ,
1810	 => std_logic_vector(to_unsigned(82,8) ,
1811	 => std_logic_vector(to_unsigned(84,8) ,
1812	 => std_logic_vector(to_unsigned(87,8) ,
1813	 => std_logic_vector(to_unsigned(87,8) ,
1814	 => std_logic_vector(to_unsigned(90,8) ,
1815	 => std_logic_vector(to_unsigned(86,8) ,
1816	 => std_logic_vector(to_unsigned(86,8) ,
1817	 => std_logic_vector(to_unsigned(87,8) ,
1818	 => std_logic_vector(to_unsigned(88,8) ,
1819	 => std_logic_vector(to_unsigned(88,8) ,
1820	 => std_logic_vector(to_unsigned(86,8) ,
1821	 => std_logic_vector(to_unsigned(87,8) ,
1822	 => std_logic_vector(to_unsigned(91,8) ,
1823	 => std_logic_vector(to_unsigned(88,8) ,
1824	 => std_logic_vector(to_unsigned(91,8) ,
1825	 => std_logic_vector(to_unsigned(92,8) ,
1826	 => std_logic_vector(to_unsigned(88,8) ,
1827	 => std_logic_vector(to_unsigned(91,8) ,
1828	 => std_logic_vector(to_unsigned(92,8) ,
1829	 => std_logic_vector(to_unsigned(96,8) ,
1830	 => std_logic_vector(to_unsigned(96,8) ,
1831	 => std_logic_vector(to_unsigned(90,8) ,
1832	 => std_logic_vector(to_unsigned(84,8) ,
1833	 => std_logic_vector(to_unsigned(82,8) ,
1834	 => std_logic_vector(to_unsigned(86,8) ,
1835	 => std_logic_vector(to_unsigned(92,8) ,
1836	 => std_logic_vector(to_unsigned(25,8) ,
1837	 => std_logic_vector(to_unsigned(0,8) ,
1838	 => std_logic_vector(to_unsigned(0,8) ,
1839	 => std_logic_vector(to_unsigned(2,8) ,
1840	 => std_logic_vector(to_unsigned(70,8) ,
1841	 => std_logic_vector(to_unsigned(99,8) ,
1842	 => std_logic_vector(to_unsigned(81,8) ,
1843	 => std_logic_vector(to_unsigned(91,8) ,
1844	 => std_logic_vector(to_unsigned(96,8) ,
1845	 => std_logic_vector(to_unsigned(93,8) ,
1846	 => std_logic_vector(to_unsigned(96,8) ,
1847	 => std_logic_vector(to_unsigned(101,8) ,
1848	 => std_logic_vector(to_unsigned(101,8) ,
1849	 => std_logic_vector(to_unsigned(101,8) ,
1850	 => std_logic_vector(to_unsigned(104,8) ,
1851	 => std_logic_vector(to_unsigned(105,8) ,
1852	 => std_logic_vector(to_unsigned(111,8) ,
1853	 => std_logic_vector(to_unsigned(115,8) ,
1854	 => std_logic_vector(to_unsigned(107,8) ,
1855	 => std_logic_vector(to_unsigned(107,8) ,
1856	 => std_logic_vector(to_unsigned(109,8) ,
1857	 => std_logic_vector(to_unsigned(108,8) ,
1858	 => std_logic_vector(to_unsigned(111,8) ,
1859	 => std_logic_vector(to_unsigned(111,8) ,
1860	 => std_logic_vector(to_unsigned(112,8) ,
1861	 => std_logic_vector(to_unsigned(111,8) ,
1862	 => std_logic_vector(to_unsigned(108,8) ,
1863	 => std_logic_vector(to_unsigned(112,8) ,
1864	 => std_logic_vector(to_unsigned(116,8) ,
1865	 => std_logic_vector(to_unsigned(112,8) ,
1866	 => std_logic_vector(to_unsigned(109,8) ,
1867	 => std_logic_vector(to_unsigned(105,8) ,
1868	 => std_logic_vector(to_unsigned(105,8) ,
1869	 => std_logic_vector(to_unsigned(114,8) ,
1870	 => std_logic_vector(to_unsigned(118,8) ,
1871	 => std_logic_vector(to_unsigned(116,8) ,
1872	 => std_logic_vector(to_unsigned(116,8) ,
1873	 => std_logic_vector(to_unsigned(116,8) ,
1874	 => std_logic_vector(to_unsigned(119,8) ,
1875	 => std_logic_vector(to_unsigned(127,8) ,
1876	 => std_logic_vector(to_unsigned(138,8) ,
1877	 => std_logic_vector(to_unsigned(139,8) ,
1878	 => std_logic_vector(to_unsigned(131,8) ,
1879	 => std_logic_vector(to_unsigned(136,8) ,
1880	 => std_logic_vector(to_unsigned(139,8) ,
1881	 => std_logic_vector(to_unsigned(144,8) ,
1882	 => std_logic_vector(to_unsigned(146,8) ,
1883	 => std_logic_vector(to_unsigned(144,8) ,
1884	 => std_logic_vector(to_unsigned(142,8) ,
1885	 => std_logic_vector(to_unsigned(144,8) ,
1886	 => std_logic_vector(to_unsigned(151,8) ,
1887	 => std_logic_vector(to_unsigned(149,8) ,
1888	 => std_logic_vector(to_unsigned(142,8) ,
1889	 => std_logic_vector(to_unsigned(141,8) ,
1890	 => std_logic_vector(to_unsigned(144,8) ,
1891	 => std_logic_vector(to_unsigned(146,8) ,
1892	 => std_logic_vector(to_unsigned(149,8) ,
1893	 => std_logic_vector(to_unsigned(149,8) ,
1894	 => std_logic_vector(to_unsigned(147,8) ,
1895	 => std_logic_vector(to_unsigned(151,8) ,
1896	 => std_logic_vector(to_unsigned(154,8) ,
1897	 => std_logic_vector(to_unsigned(156,8) ,
1898	 => std_logic_vector(to_unsigned(157,8) ,
1899	 => std_logic_vector(to_unsigned(159,8) ,
1900	 => std_logic_vector(to_unsigned(157,8) ,
1901	 => std_logic_vector(to_unsigned(161,8) ,
1902	 => std_logic_vector(to_unsigned(161,8) ,
1903	 => std_logic_vector(to_unsigned(161,8) ,
1904	 => std_logic_vector(to_unsigned(163,8) ,
1905	 => std_logic_vector(to_unsigned(159,8) ,
1906	 => std_logic_vector(to_unsigned(156,8) ,
1907	 => std_logic_vector(to_unsigned(157,8) ,
1908	 => std_logic_vector(to_unsigned(159,8) ,
1909	 => std_logic_vector(to_unsigned(159,8) ,
1910	 => std_logic_vector(to_unsigned(159,8) ,
1911	 => std_logic_vector(to_unsigned(161,8) ,
1912	 => std_logic_vector(to_unsigned(159,8) ,
1913	 => std_logic_vector(to_unsigned(156,8) ,
1914	 => std_logic_vector(to_unsigned(159,8) ,
1915	 => std_logic_vector(to_unsigned(163,8) ,
1916	 => std_logic_vector(to_unsigned(161,8) ,
1917	 => std_logic_vector(to_unsigned(161,8) ,
1918	 => std_logic_vector(to_unsigned(161,8) ,
1919	 => std_logic_vector(to_unsigned(163,8) ,
1920	 => std_logic_vector(to_unsigned(161,8) ,
1921	 => std_logic_vector(to_unsigned(100,8) ,
1922	 => std_logic_vector(to_unsigned(92,8) ,
1923	 => std_logic_vector(to_unsigned(101,8) ,
1924	 => std_logic_vector(to_unsigned(99,8) ,
1925	 => std_logic_vector(to_unsigned(91,8) ,
1926	 => std_logic_vector(to_unsigned(99,8) ,
1927	 => std_logic_vector(to_unsigned(100,8) ,
1928	 => std_logic_vector(to_unsigned(99,8) ,
1929	 => std_logic_vector(to_unsigned(96,8) ,
1930	 => std_logic_vector(to_unsigned(100,8) ,
1931	 => std_logic_vector(to_unsigned(93,8) ,
1932	 => std_logic_vector(to_unsigned(93,8) ,
1933	 => std_logic_vector(to_unsigned(97,8) ,
1934	 => std_logic_vector(to_unsigned(91,8) ,
1935	 => std_logic_vector(to_unsigned(91,8) ,
1936	 => std_logic_vector(to_unsigned(93,8) ,
1937	 => std_logic_vector(to_unsigned(93,8) ,
1938	 => std_logic_vector(to_unsigned(88,8) ,
1939	 => std_logic_vector(to_unsigned(86,8) ,
1940	 => std_logic_vector(to_unsigned(88,8) ,
1941	 => std_logic_vector(to_unsigned(86,8) ,
1942	 => std_logic_vector(to_unsigned(90,8) ,
1943	 => std_logic_vector(to_unsigned(90,8) ,
1944	 => std_logic_vector(to_unsigned(90,8) ,
1945	 => std_logic_vector(to_unsigned(88,8) ,
1946	 => std_logic_vector(to_unsigned(86,8) ,
1947	 => std_logic_vector(to_unsigned(95,8) ,
1948	 => std_logic_vector(to_unsigned(99,8) ,
1949	 => std_logic_vector(to_unsigned(100,8) ,
1950	 => std_logic_vector(to_unsigned(100,8) ,
1951	 => std_logic_vector(to_unsigned(100,8) ,
1952	 => std_logic_vector(to_unsigned(95,8) ,
1953	 => std_logic_vector(to_unsigned(99,8) ,
1954	 => std_logic_vector(to_unsigned(96,8) ,
1955	 => std_logic_vector(to_unsigned(86,8) ,
1956	 => std_logic_vector(to_unsigned(92,8) ,
1957	 => std_logic_vector(to_unsigned(95,8) ,
1958	 => std_logic_vector(to_unsigned(99,8) ,
1959	 => std_logic_vector(to_unsigned(105,8) ,
1960	 => std_logic_vector(to_unsigned(105,8) ,
1961	 => std_logic_vector(to_unsigned(104,8) ,
1962	 => std_logic_vector(to_unsigned(103,8) ,
1963	 => std_logic_vector(to_unsigned(101,8) ,
1964	 => std_logic_vector(to_unsigned(103,8) ,
1965	 => std_logic_vector(to_unsigned(107,8) ,
1966	 => std_logic_vector(to_unsigned(109,8) ,
1967	 => std_logic_vector(to_unsigned(109,8) ,
1968	 => std_logic_vector(to_unsigned(109,8) ,
1969	 => std_logic_vector(to_unsigned(109,8) ,
1970	 => std_logic_vector(to_unsigned(116,8) ,
1971	 => std_logic_vector(to_unsigned(111,8) ,
1972	 => std_logic_vector(to_unsigned(101,8) ,
1973	 => std_logic_vector(to_unsigned(108,8) ,
1974	 => std_logic_vector(to_unsigned(107,8) ,
1975	 => std_logic_vector(to_unsigned(96,8) ,
1976	 => std_logic_vector(to_unsigned(103,8) ,
1977	 => std_logic_vector(to_unsigned(109,8) ,
1978	 => std_logic_vector(to_unsigned(108,8) ,
1979	 => std_logic_vector(to_unsigned(109,8) ,
1980	 => std_logic_vector(to_unsigned(114,8) ,
1981	 => std_logic_vector(to_unsigned(109,8) ,
1982	 => std_logic_vector(to_unsigned(107,8) ,
1983	 => std_logic_vector(to_unsigned(105,8) ,
1984	 => std_logic_vector(to_unsigned(107,8) ,
1985	 => std_logic_vector(to_unsigned(111,8) ,
1986	 => std_logic_vector(to_unsigned(107,8) ,
1987	 => std_logic_vector(to_unsigned(107,8) ,
1988	 => std_logic_vector(to_unsigned(105,8) ,
1989	 => std_logic_vector(to_unsigned(105,8) ,
1990	 => std_logic_vector(to_unsigned(114,8) ,
1991	 => std_logic_vector(to_unsigned(115,8) ,
1992	 => std_logic_vector(to_unsigned(114,8) ,
1993	 => std_logic_vector(to_unsigned(115,8) ,
1994	 => std_logic_vector(to_unsigned(118,8) ,
1995	 => std_logic_vector(to_unsigned(114,8) ,
1996	 => std_logic_vector(to_unsigned(111,8) ,
1997	 => std_logic_vector(to_unsigned(114,8) ,
1998	 => std_logic_vector(to_unsigned(109,8) ,
1999	 => std_logic_vector(to_unsigned(105,8) ,
2000	 => std_logic_vector(to_unsigned(108,8) ,
2001	 => std_logic_vector(to_unsigned(104,8) ,
2002	 => std_logic_vector(to_unsigned(107,8) ,
2003	 => std_logic_vector(to_unsigned(108,8) ,
2004	 => std_logic_vector(to_unsigned(116,8) ,
2005	 => std_logic_vector(to_unsigned(108,8) ,
2006	 => std_logic_vector(to_unsigned(105,8) ,
2007	 => std_logic_vector(to_unsigned(108,8) ,
2008	 => std_logic_vector(to_unsigned(108,8) ,
2009	 => std_logic_vector(to_unsigned(104,8) ,
2010	 => std_logic_vector(to_unsigned(105,8) ,
2011	 => std_logic_vector(to_unsigned(107,8) ,
2012	 => std_logic_vector(to_unsigned(104,8) ,
2013	 => std_logic_vector(to_unsigned(109,8) ,
2014	 => std_logic_vector(to_unsigned(100,8) ,
2015	 => std_logic_vector(to_unsigned(96,8) ,
2016	 => std_logic_vector(to_unsigned(97,8) ,
2017	 => std_logic_vector(to_unsigned(96,8) ,
2018	 => std_logic_vector(to_unsigned(100,8) ,
2019	 => std_logic_vector(to_unsigned(99,8) ,
2020	 => std_logic_vector(to_unsigned(96,8) ,
2021	 => std_logic_vector(to_unsigned(96,8) ,
2022	 => std_logic_vector(to_unsigned(100,8) ,
2023	 => std_logic_vector(to_unsigned(100,8) ,
2024	 => std_logic_vector(to_unsigned(99,8) ,
2025	 => std_logic_vector(to_unsigned(100,8) ,
2026	 => std_logic_vector(to_unsigned(104,8) ,
2027	 => std_logic_vector(to_unsigned(105,8) ,
2028	 => std_logic_vector(to_unsigned(112,8) ,
2029	 => std_logic_vector(to_unsigned(111,8) ,
2030	 => std_logic_vector(to_unsigned(105,8) ,
2031	 => std_logic_vector(to_unsigned(105,8) ,
2032	 => std_logic_vector(to_unsigned(109,8) ,
2033	 => std_logic_vector(to_unsigned(111,8) ,
2034	 => std_logic_vector(to_unsigned(108,8) ,
2035	 => std_logic_vector(to_unsigned(104,8) ,
2036	 => std_logic_vector(to_unsigned(100,8) ,
2037	 => std_logic_vector(to_unsigned(105,8) ,
2038	 => std_logic_vector(to_unsigned(108,8) ,
2039	 => std_logic_vector(to_unsigned(101,8) ,
2040	 => std_logic_vector(to_unsigned(101,8) ,
2041	 => std_logic_vector(to_unsigned(101,8) ,
2042	 => std_logic_vector(to_unsigned(100,8) ,
2043	 => std_logic_vector(to_unsigned(100,8) ,
2044	 => std_logic_vector(to_unsigned(100,8) ,
2045	 => std_logic_vector(to_unsigned(97,8) ,
2046	 => std_logic_vector(to_unsigned(95,8) ,
2047	 => std_logic_vector(to_unsigned(99,8) ,
2048	 => std_logic_vector(to_unsigned(96,8) ,
2049	 => std_logic_vector(to_unsigned(93,8) ,
2050	 => std_logic_vector(to_unsigned(93,8) ,
2051	 => std_logic_vector(to_unsigned(93,8) ,
2052	 => std_logic_vector(to_unsigned(93,8) ,
2053	 => std_logic_vector(to_unsigned(96,8) ,
2054	 => std_logic_vector(to_unsigned(96,8) ,
2055	 => std_logic_vector(to_unsigned(92,8) ,
2056	 => std_logic_vector(to_unsigned(92,8) ,
2057	 => std_logic_vector(to_unsigned(96,8) ,
2058	 => std_logic_vector(to_unsigned(97,8) ,
2059	 => std_logic_vector(to_unsigned(95,8) ,
2060	 => std_logic_vector(to_unsigned(97,8) ,
2061	 => std_logic_vector(to_unsigned(97,8) ,
2062	 => std_logic_vector(to_unsigned(96,8) ,
2063	 => std_logic_vector(to_unsigned(100,8) ,
2064	 => std_logic_vector(to_unsigned(104,8) ,
2065	 => std_logic_vector(to_unsigned(107,8) ,
2066	 => std_logic_vector(to_unsigned(103,8) ,
2067	 => std_logic_vector(to_unsigned(103,8) ,
2068	 => std_logic_vector(to_unsigned(100,8) ,
2069	 => std_logic_vector(to_unsigned(103,8) ,
2070	 => std_logic_vector(to_unsigned(101,8) ,
2071	 => std_logic_vector(to_unsigned(96,8) ,
2072	 => std_logic_vector(to_unsigned(97,8) ,
2073	 => std_logic_vector(to_unsigned(97,8) ,
2074	 => std_logic_vector(to_unsigned(95,8) ,
2075	 => std_logic_vector(to_unsigned(90,8) ,
2076	 => std_logic_vector(to_unsigned(85,8) ,
2077	 => std_logic_vector(to_unsigned(81,8) ,
2078	 => std_logic_vector(to_unsigned(82,8) ,
2079	 => std_logic_vector(to_unsigned(86,8) ,
2080	 => std_logic_vector(to_unsigned(88,8) ,
2081	 => std_logic_vector(to_unsigned(84,8) ,
2082	 => std_logic_vector(to_unsigned(87,8) ,
2083	 => std_logic_vector(to_unsigned(84,8) ,
2084	 => std_logic_vector(to_unsigned(84,8) ,
2085	 => std_logic_vector(to_unsigned(84,8) ,
2086	 => std_logic_vector(to_unsigned(85,8) ,
2087	 => std_logic_vector(to_unsigned(87,8) ,
2088	 => std_logic_vector(to_unsigned(87,8) ,
2089	 => std_logic_vector(to_unsigned(87,8) ,
2090	 => std_logic_vector(to_unsigned(88,8) ,
2091	 => std_logic_vector(to_unsigned(82,8) ,
2092	 => std_logic_vector(to_unsigned(88,8) ,
2093	 => std_logic_vector(to_unsigned(90,8) ,
2094	 => std_logic_vector(to_unsigned(82,8) ,
2095	 => std_logic_vector(to_unsigned(86,8) ,
2096	 => std_logic_vector(to_unsigned(87,8) ,
2097	 => std_logic_vector(to_unsigned(87,8) ,
2098	 => std_logic_vector(to_unsigned(87,8) ,
2099	 => std_logic_vector(to_unsigned(88,8) ,
2100	 => std_logic_vector(to_unsigned(87,8) ,
2101	 => std_logic_vector(to_unsigned(85,8) ,
2102	 => std_logic_vector(to_unsigned(78,8) ,
2103	 => std_logic_vector(to_unsigned(78,8) ,
2104	 => std_logic_vector(to_unsigned(82,8) ,
2105	 => std_logic_vector(to_unsigned(77,8) ,
2106	 => std_logic_vector(to_unsigned(79,8) ,
2107	 => std_logic_vector(to_unsigned(82,8) ,
2108	 => std_logic_vector(to_unsigned(88,8) ,
2109	 => std_logic_vector(to_unsigned(82,8) ,
2110	 => std_logic_vector(to_unsigned(77,8) ,
2111	 => std_logic_vector(to_unsigned(79,8) ,
2112	 => std_logic_vector(to_unsigned(78,8) ,
2113	 => std_logic_vector(to_unsigned(85,8) ,
2114	 => std_logic_vector(to_unsigned(93,8) ,
2115	 => std_logic_vector(to_unsigned(84,8) ,
2116	 => std_logic_vector(to_unsigned(81,8) ,
2117	 => std_logic_vector(to_unsigned(86,8) ,
2118	 => std_logic_vector(to_unsigned(84,8) ,
2119	 => std_logic_vector(to_unsigned(85,8) ,
2120	 => std_logic_vector(to_unsigned(87,8) ,
2121	 => std_logic_vector(to_unsigned(86,8) ,
2122	 => std_logic_vector(to_unsigned(82,8) ,
2123	 => std_logic_vector(to_unsigned(84,8) ,
2124	 => std_logic_vector(to_unsigned(86,8) ,
2125	 => std_logic_vector(to_unsigned(87,8) ,
2126	 => std_logic_vector(to_unsigned(86,8) ,
2127	 => std_logic_vector(to_unsigned(84,8) ,
2128	 => std_logic_vector(to_unsigned(86,8) ,
2129	 => std_logic_vector(to_unsigned(84,8) ,
2130	 => std_logic_vector(to_unsigned(81,8) ,
2131	 => std_logic_vector(to_unsigned(84,8) ,
2132	 => std_logic_vector(to_unsigned(81,8) ,
2133	 => std_logic_vector(to_unsigned(85,8) ,
2134	 => std_logic_vector(to_unsigned(87,8) ,
2135	 => std_logic_vector(to_unsigned(85,8) ,
2136	 => std_logic_vector(to_unsigned(82,8) ,
2137	 => std_logic_vector(to_unsigned(86,8) ,
2138	 => std_logic_vector(to_unsigned(91,8) ,
2139	 => std_logic_vector(to_unsigned(87,8) ,
2140	 => std_logic_vector(to_unsigned(84,8) ,
2141	 => std_logic_vector(to_unsigned(87,8) ,
2142	 => std_logic_vector(to_unsigned(90,8) ,
2143	 => std_logic_vector(to_unsigned(88,8) ,
2144	 => std_logic_vector(to_unsigned(86,8) ,
2145	 => std_logic_vector(to_unsigned(86,8) ,
2146	 => std_logic_vector(to_unsigned(88,8) ,
2147	 => std_logic_vector(to_unsigned(92,8) ,
2148	 => std_logic_vector(to_unsigned(91,8) ,
2149	 => std_logic_vector(to_unsigned(90,8) ,
2150	 => std_logic_vector(to_unsigned(95,8) ,
2151	 => std_logic_vector(to_unsigned(88,8) ,
2152	 => std_logic_vector(to_unsigned(86,8) ,
2153	 => std_logic_vector(to_unsigned(92,8) ,
2154	 => std_logic_vector(to_unsigned(81,8) ,
2155	 => std_logic_vector(to_unsigned(85,8) ,
2156	 => std_logic_vector(to_unsigned(50,8) ,
2157	 => std_logic_vector(to_unsigned(2,8) ,
2158	 => std_logic_vector(to_unsigned(0,8) ,
2159	 => std_logic_vector(to_unsigned(1,8) ,
2160	 => std_logic_vector(to_unsigned(45,8) ,
2161	 => std_logic_vector(to_unsigned(101,8) ,
2162	 => std_logic_vector(to_unsigned(80,8) ,
2163	 => std_logic_vector(to_unsigned(97,8) ,
2164	 => std_logic_vector(to_unsigned(100,8) ,
2165	 => std_logic_vector(to_unsigned(92,8) ,
2166	 => std_logic_vector(to_unsigned(95,8) ,
2167	 => std_logic_vector(to_unsigned(97,8) ,
2168	 => std_logic_vector(to_unsigned(101,8) ,
2169	 => std_logic_vector(to_unsigned(99,8) ,
2170	 => std_logic_vector(to_unsigned(99,8) ,
2171	 => std_logic_vector(to_unsigned(107,8) ,
2172	 => std_logic_vector(to_unsigned(111,8) ,
2173	 => std_logic_vector(to_unsigned(114,8) ,
2174	 => std_logic_vector(to_unsigned(109,8) ,
2175	 => std_logic_vector(to_unsigned(107,8) ,
2176	 => std_logic_vector(to_unsigned(112,8) ,
2177	 => std_logic_vector(to_unsigned(109,8) ,
2178	 => std_logic_vector(to_unsigned(105,8) ,
2179	 => std_logic_vector(to_unsigned(108,8) ,
2180	 => std_logic_vector(to_unsigned(116,8) ,
2181	 => std_logic_vector(to_unsigned(115,8) ,
2182	 => std_logic_vector(to_unsigned(109,8) ,
2183	 => std_logic_vector(to_unsigned(114,8) ,
2184	 => std_logic_vector(to_unsigned(114,8) ,
2185	 => std_logic_vector(to_unsigned(111,8) ,
2186	 => std_logic_vector(to_unsigned(104,8) ,
2187	 => std_logic_vector(to_unsigned(104,8) ,
2188	 => std_logic_vector(to_unsigned(109,8) ,
2189	 => std_logic_vector(to_unsigned(115,8) ,
2190	 => std_logic_vector(to_unsigned(115,8) ,
2191	 => std_logic_vector(to_unsigned(116,8) ,
2192	 => std_logic_vector(to_unsigned(114,8) ,
2193	 => std_logic_vector(to_unsigned(118,8) ,
2194	 => std_logic_vector(to_unsigned(124,8) ,
2195	 => std_logic_vector(to_unsigned(130,8) ,
2196	 => std_logic_vector(to_unsigned(133,8) ,
2197	 => std_logic_vector(to_unsigned(131,8) ,
2198	 => std_logic_vector(to_unsigned(128,8) ,
2199	 => std_logic_vector(to_unsigned(136,8) ,
2200	 => std_logic_vector(to_unsigned(138,8) ,
2201	 => std_logic_vector(to_unsigned(138,8) ,
2202	 => std_logic_vector(to_unsigned(138,8) ,
2203	 => std_logic_vector(to_unsigned(144,8) ,
2204	 => std_logic_vector(to_unsigned(147,8) ,
2205	 => std_logic_vector(to_unsigned(146,8) ,
2206	 => std_logic_vector(to_unsigned(144,8) ,
2207	 => std_logic_vector(to_unsigned(147,8) ,
2208	 => std_logic_vector(to_unsigned(146,8) ,
2209	 => std_logic_vector(to_unsigned(146,8) ,
2210	 => std_logic_vector(to_unsigned(151,8) ,
2211	 => std_logic_vector(to_unsigned(151,8) ,
2212	 => std_logic_vector(to_unsigned(149,8) ,
2213	 => std_logic_vector(to_unsigned(149,8) ,
2214	 => std_logic_vector(to_unsigned(151,8) ,
2215	 => std_logic_vector(to_unsigned(156,8) ,
2216	 => std_logic_vector(to_unsigned(157,8) ,
2217	 => std_logic_vector(to_unsigned(156,8) ,
2218	 => std_logic_vector(to_unsigned(157,8) ,
2219	 => std_logic_vector(to_unsigned(156,8) ,
2220	 => std_logic_vector(to_unsigned(157,8) ,
2221	 => std_logic_vector(to_unsigned(159,8) ,
2222	 => std_logic_vector(to_unsigned(163,8) ,
2223	 => std_logic_vector(to_unsigned(161,8) ,
2224	 => std_logic_vector(to_unsigned(159,8) ,
2225	 => std_logic_vector(to_unsigned(159,8) ,
2226	 => std_logic_vector(to_unsigned(159,8) ,
2227	 => std_logic_vector(to_unsigned(159,8) ,
2228	 => std_logic_vector(to_unsigned(161,8) ,
2229	 => std_logic_vector(to_unsigned(159,8) ,
2230	 => std_logic_vector(to_unsigned(157,8) ,
2231	 => std_logic_vector(to_unsigned(156,8) ,
2232	 => std_logic_vector(to_unsigned(157,8) ,
2233	 => std_logic_vector(to_unsigned(157,8) ,
2234	 => std_logic_vector(to_unsigned(161,8) ,
2235	 => std_logic_vector(to_unsigned(157,8) ,
2236	 => std_logic_vector(to_unsigned(156,8) ,
2237	 => std_logic_vector(to_unsigned(163,8) ,
2238	 => std_logic_vector(to_unsigned(164,8) ,
2239	 => std_logic_vector(to_unsigned(164,8) ,
2240	 => std_logic_vector(to_unsigned(164,8) ,
2241	 => std_logic_vector(to_unsigned(101,8) ,
2242	 => std_logic_vector(to_unsigned(101,8) ,
2243	 => std_logic_vector(to_unsigned(103,8) ,
2244	 => std_logic_vector(to_unsigned(93,8) ,
2245	 => std_logic_vector(to_unsigned(91,8) ,
2246	 => std_logic_vector(to_unsigned(97,8) ,
2247	 => std_logic_vector(to_unsigned(96,8) ,
2248	 => std_logic_vector(to_unsigned(95,8) ,
2249	 => std_logic_vector(to_unsigned(90,8) ,
2250	 => std_logic_vector(to_unsigned(90,8) ,
2251	 => std_logic_vector(to_unsigned(90,8) ,
2252	 => std_logic_vector(to_unsigned(90,8) ,
2253	 => std_logic_vector(to_unsigned(95,8) ,
2254	 => std_logic_vector(to_unsigned(92,8) ,
2255	 => std_logic_vector(to_unsigned(92,8) ,
2256	 => std_logic_vector(to_unsigned(86,8) ,
2257	 => std_logic_vector(to_unsigned(87,8) ,
2258	 => std_logic_vector(to_unsigned(87,8) ,
2259	 => std_logic_vector(to_unsigned(90,8) ,
2260	 => std_logic_vector(to_unsigned(93,8) ,
2261	 => std_logic_vector(to_unsigned(91,8) ,
2262	 => std_logic_vector(to_unsigned(91,8) ,
2263	 => std_logic_vector(to_unsigned(88,8) ,
2264	 => std_logic_vector(to_unsigned(87,8) ,
2265	 => std_logic_vector(to_unsigned(88,8) ,
2266	 => std_logic_vector(to_unsigned(86,8) ,
2267	 => std_logic_vector(to_unsigned(90,8) ,
2268	 => std_logic_vector(to_unsigned(91,8) ,
2269	 => std_logic_vector(to_unsigned(91,8) ,
2270	 => std_logic_vector(to_unsigned(92,8) ,
2271	 => std_logic_vector(to_unsigned(96,8) ,
2272	 => std_logic_vector(to_unsigned(93,8) ,
2273	 => std_logic_vector(to_unsigned(93,8) ,
2274	 => std_logic_vector(to_unsigned(91,8) ,
2275	 => std_logic_vector(to_unsigned(90,8) ,
2276	 => std_logic_vector(to_unsigned(97,8) ,
2277	 => std_logic_vector(to_unsigned(97,8) ,
2278	 => std_logic_vector(to_unsigned(96,8) ,
2279	 => std_logic_vector(to_unsigned(100,8) ,
2280	 => std_logic_vector(to_unsigned(99,8) ,
2281	 => std_logic_vector(to_unsigned(97,8) ,
2282	 => std_logic_vector(to_unsigned(100,8) ,
2283	 => std_logic_vector(to_unsigned(99,8) ,
2284	 => std_logic_vector(to_unsigned(101,8) ,
2285	 => std_logic_vector(to_unsigned(103,8) ,
2286	 => std_logic_vector(to_unsigned(104,8) ,
2287	 => std_logic_vector(to_unsigned(103,8) ,
2288	 => std_logic_vector(to_unsigned(105,8) ,
2289	 => std_logic_vector(to_unsigned(105,8) ,
2290	 => std_logic_vector(to_unsigned(105,8) ,
2291	 => std_logic_vector(to_unsigned(99,8) ,
2292	 => std_logic_vector(to_unsigned(101,8) ,
2293	 => std_logic_vector(to_unsigned(103,8) ,
2294	 => std_logic_vector(to_unsigned(103,8) ,
2295	 => std_logic_vector(to_unsigned(107,8) ,
2296	 => std_logic_vector(to_unsigned(105,8) ,
2297	 => std_logic_vector(to_unsigned(103,8) ,
2298	 => std_logic_vector(to_unsigned(111,8) ,
2299	 => std_logic_vector(to_unsigned(111,8) ,
2300	 => std_logic_vector(to_unsigned(109,8) ,
2301	 => std_logic_vector(to_unsigned(105,8) ,
2302	 => std_logic_vector(to_unsigned(108,8) ,
2303	 => std_logic_vector(to_unsigned(108,8) ,
2304	 => std_logic_vector(to_unsigned(103,8) ,
2305	 => std_logic_vector(to_unsigned(103,8) ,
2306	 => std_logic_vector(to_unsigned(104,8) ,
2307	 => std_logic_vector(to_unsigned(107,8) ,
2308	 => std_logic_vector(to_unsigned(109,8) ,
2309	 => std_logic_vector(to_unsigned(109,8) ,
2310	 => std_logic_vector(to_unsigned(112,8) ,
2311	 => std_logic_vector(to_unsigned(114,8) ,
2312	 => std_logic_vector(to_unsigned(114,8) ,
2313	 => std_logic_vector(to_unsigned(112,8) ,
2314	 => std_logic_vector(to_unsigned(111,8) ,
2315	 => std_logic_vector(to_unsigned(109,8) ,
2316	 => std_logic_vector(to_unsigned(108,8) ,
2317	 => std_logic_vector(to_unsigned(111,8) ,
2318	 => std_logic_vector(to_unsigned(108,8) ,
2319	 => std_logic_vector(to_unsigned(109,8) ,
2320	 => std_logic_vector(to_unsigned(111,8) ,
2321	 => std_logic_vector(to_unsigned(104,8) ,
2322	 => std_logic_vector(to_unsigned(105,8) ,
2323	 => std_logic_vector(to_unsigned(108,8) ,
2324	 => std_logic_vector(to_unsigned(107,8) ,
2325	 => std_logic_vector(to_unsigned(109,8) ,
2326	 => std_logic_vector(to_unsigned(105,8) ,
2327	 => std_logic_vector(to_unsigned(104,8) ,
2328	 => std_logic_vector(to_unsigned(108,8) ,
2329	 => std_logic_vector(to_unsigned(103,8) ,
2330	 => std_logic_vector(to_unsigned(103,8) ,
2331	 => std_logic_vector(to_unsigned(103,8) ,
2332	 => std_logic_vector(to_unsigned(103,8) ,
2333	 => std_logic_vector(to_unsigned(101,8) ,
2334	 => std_logic_vector(to_unsigned(93,8) ,
2335	 => std_logic_vector(to_unsigned(95,8) ,
2336	 => std_logic_vector(to_unsigned(101,8) ,
2337	 => std_logic_vector(to_unsigned(100,8) ,
2338	 => std_logic_vector(to_unsigned(97,8) ,
2339	 => std_logic_vector(to_unsigned(95,8) ,
2340	 => std_logic_vector(to_unsigned(92,8) ,
2341	 => std_logic_vector(to_unsigned(91,8) ,
2342	 => std_logic_vector(to_unsigned(95,8) ,
2343	 => std_logic_vector(to_unsigned(97,8) ,
2344	 => std_logic_vector(to_unsigned(97,8) ,
2345	 => std_logic_vector(to_unsigned(99,8) ,
2346	 => std_logic_vector(to_unsigned(99,8) ,
2347	 => std_logic_vector(to_unsigned(104,8) ,
2348	 => std_logic_vector(to_unsigned(111,8) ,
2349	 => std_logic_vector(to_unsigned(112,8) ,
2350	 => std_logic_vector(to_unsigned(109,8) ,
2351	 => std_logic_vector(to_unsigned(105,8) ,
2352	 => std_logic_vector(to_unsigned(108,8) ,
2353	 => std_logic_vector(to_unsigned(107,8) ,
2354	 => std_logic_vector(to_unsigned(107,8) ,
2355	 => std_logic_vector(to_unsigned(105,8) ,
2356	 => std_logic_vector(to_unsigned(101,8) ,
2357	 => std_logic_vector(to_unsigned(104,8) ,
2358	 => std_logic_vector(to_unsigned(101,8) ,
2359	 => std_logic_vector(to_unsigned(100,8) ,
2360	 => std_logic_vector(to_unsigned(104,8) ,
2361	 => std_logic_vector(to_unsigned(105,8) ,
2362	 => std_logic_vector(to_unsigned(104,8) ,
2363	 => std_logic_vector(to_unsigned(100,8) ,
2364	 => std_logic_vector(to_unsigned(97,8) ,
2365	 => std_logic_vector(to_unsigned(96,8) ,
2366	 => std_logic_vector(to_unsigned(95,8) ,
2367	 => std_logic_vector(to_unsigned(95,8) ,
2368	 => std_logic_vector(to_unsigned(92,8) ,
2369	 => std_logic_vector(to_unsigned(92,8) ,
2370	 => std_logic_vector(to_unsigned(91,8) ,
2371	 => std_logic_vector(to_unsigned(92,8) ,
2372	 => std_logic_vector(to_unsigned(92,8) ,
2373	 => std_logic_vector(to_unsigned(91,8) ,
2374	 => std_logic_vector(to_unsigned(92,8) ,
2375	 => std_logic_vector(to_unsigned(90,8) ,
2376	 => std_logic_vector(to_unsigned(91,8) ,
2377	 => std_logic_vector(to_unsigned(95,8) ,
2378	 => std_logic_vector(to_unsigned(93,8) ,
2379	 => std_logic_vector(to_unsigned(96,8) ,
2380	 => std_logic_vector(to_unsigned(99,8) ,
2381	 => std_logic_vector(to_unsigned(96,8) ,
2382	 => std_logic_vector(to_unsigned(96,8) ,
2383	 => std_logic_vector(to_unsigned(99,8) ,
2384	 => std_logic_vector(to_unsigned(103,8) ,
2385	 => std_logic_vector(to_unsigned(105,8) ,
2386	 => std_logic_vector(to_unsigned(105,8) ,
2387	 => std_logic_vector(to_unsigned(101,8) ,
2388	 => std_logic_vector(to_unsigned(97,8) ,
2389	 => std_logic_vector(to_unsigned(97,8) ,
2390	 => std_logic_vector(to_unsigned(101,8) ,
2391	 => std_logic_vector(to_unsigned(103,8) ,
2392	 => std_logic_vector(to_unsigned(103,8) ,
2393	 => std_logic_vector(to_unsigned(93,8) ,
2394	 => std_logic_vector(to_unsigned(88,8) ,
2395	 => std_logic_vector(to_unsigned(88,8) ,
2396	 => std_logic_vector(to_unsigned(90,8) ,
2397	 => std_logic_vector(to_unsigned(87,8) ,
2398	 => std_logic_vector(to_unsigned(88,8) ,
2399	 => std_logic_vector(to_unsigned(91,8) ,
2400	 => std_logic_vector(to_unsigned(90,8) ,
2401	 => std_logic_vector(to_unsigned(85,8) ,
2402	 => std_logic_vector(to_unsigned(86,8) ,
2403	 => std_logic_vector(to_unsigned(87,8) ,
2404	 => std_logic_vector(to_unsigned(85,8) ,
2405	 => std_logic_vector(to_unsigned(86,8) ,
2406	 => std_logic_vector(to_unsigned(90,8) ,
2407	 => std_logic_vector(to_unsigned(90,8) ,
2408	 => std_logic_vector(to_unsigned(91,8) ,
2409	 => std_logic_vector(to_unsigned(90,8) ,
2410	 => std_logic_vector(to_unsigned(92,8) ,
2411	 => std_logic_vector(to_unsigned(87,8) ,
2412	 => std_logic_vector(to_unsigned(90,8) ,
2413	 => std_logic_vector(to_unsigned(90,8) ,
2414	 => std_logic_vector(to_unsigned(87,8) ,
2415	 => std_logic_vector(to_unsigned(85,8) ,
2416	 => std_logic_vector(to_unsigned(82,8) ,
2417	 => std_logic_vector(to_unsigned(88,8) ,
2418	 => std_logic_vector(to_unsigned(91,8) ,
2419	 => std_logic_vector(to_unsigned(92,8) ,
2420	 => std_logic_vector(to_unsigned(86,8) ,
2421	 => std_logic_vector(to_unsigned(79,8) ,
2422	 => std_logic_vector(to_unsigned(77,8) ,
2423	 => std_logic_vector(to_unsigned(77,8) ,
2424	 => std_logic_vector(to_unsigned(81,8) ,
2425	 => std_logic_vector(to_unsigned(80,8) ,
2426	 => std_logic_vector(to_unsigned(78,8) ,
2427	 => std_logic_vector(to_unsigned(77,8) ,
2428	 => std_logic_vector(to_unsigned(84,8) ,
2429	 => std_logic_vector(to_unsigned(85,8) ,
2430	 => std_logic_vector(to_unsigned(79,8) ,
2431	 => std_logic_vector(to_unsigned(78,8) ,
2432	 => std_logic_vector(to_unsigned(72,8) ,
2433	 => std_logic_vector(to_unsigned(80,8) ,
2434	 => std_logic_vector(to_unsigned(86,8) ,
2435	 => std_logic_vector(to_unsigned(85,8) ,
2436	 => std_logic_vector(to_unsigned(81,8) ,
2437	 => std_logic_vector(to_unsigned(81,8) ,
2438	 => std_logic_vector(to_unsigned(85,8) ,
2439	 => std_logic_vector(to_unsigned(82,8) ,
2440	 => std_logic_vector(to_unsigned(82,8) ,
2441	 => std_logic_vector(to_unsigned(86,8) ,
2442	 => std_logic_vector(to_unsigned(82,8) ,
2443	 => std_logic_vector(to_unsigned(80,8) ,
2444	 => std_logic_vector(to_unsigned(81,8) ,
2445	 => std_logic_vector(to_unsigned(85,8) ,
2446	 => std_logic_vector(to_unsigned(91,8) ,
2447	 => std_logic_vector(to_unsigned(84,8) ,
2448	 => std_logic_vector(to_unsigned(82,8) ,
2449	 => std_logic_vector(to_unsigned(84,8) ,
2450	 => std_logic_vector(to_unsigned(81,8) ,
2451	 => std_logic_vector(to_unsigned(77,8) ,
2452	 => std_logic_vector(to_unsigned(78,8) ,
2453	 => std_logic_vector(to_unsigned(84,8) ,
2454	 => std_logic_vector(to_unsigned(85,8) ,
2455	 => std_logic_vector(to_unsigned(80,8) ,
2456	 => std_logic_vector(to_unsigned(77,8) ,
2457	 => std_logic_vector(to_unsigned(82,8) ,
2458	 => std_logic_vector(to_unsigned(84,8) ,
2459	 => std_logic_vector(to_unsigned(85,8) ,
2460	 => std_logic_vector(to_unsigned(84,8) ,
2461	 => std_logic_vector(to_unsigned(86,8) ,
2462	 => std_logic_vector(to_unsigned(91,8) ,
2463	 => std_logic_vector(to_unsigned(86,8) ,
2464	 => std_logic_vector(to_unsigned(84,8) ,
2465	 => std_logic_vector(to_unsigned(84,8) ,
2466	 => std_logic_vector(to_unsigned(88,8) ,
2467	 => std_logic_vector(to_unsigned(90,8) ,
2468	 => std_logic_vector(to_unsigned(88,8) ,
2469	 => std_logic_vector(to_unsigned(85,8) ,
2470	 => std_logic_vector(to_unsigned(86,8) ,
2471	 => std_logic_vector(to_unsigned(87,8) ,
2472	 => std_logic_vector(to_unsigned(87,8) ,
2473	 => std_logic_vector(to_unsigned(92,8) ,
2474	 => std_logic_vector(to_unsigned(82,8) ,
2475	 => std_logic_vector(to_unsigned(85,8) ,
2476	 => std_logic_vector(to_unsigned(69,8) ,
2477	 => std_logic_vector(to_unsigned(4,8) ,
2478	 => std_logic_vector(to_unsigned(0,8) ,
2479	 => std_logic_vector(to_unsigned(0,8) ,
2480	 => std_logic_vector(to_unsigned(22,8) ,
2481	 => std_logic_vector(to_unsigned(95,8) ,
2482	 => std_logic_vector(to_unsigned(80,8) ,
2483	 => std_logic_vector(to_unsigned(87,8) ,
2484	 => std_logic_vector(to_unsigned(100,8) ,
2485	 => std_logic_vector(to_unsigned(97,8) ,
2486	 => std_logic_vector(to_unsigned(92,8) ,
2487	 => std_logic_vector(to_unsigned(91,8) ,
2488	 => std_logic_vector(to_unsigned(99,8) ,
2489	 => std_logic_vector(to_unsigned(103,8) ,
2490	 => std_logic_vector(to_unsigned(100,8) ,
2491	 => std_logic_vector(to_unsigned(103,8) ,
2492	 => std_logic_vector(to_unsigned(103,8) ,
2493	 => std_logic_vector(to_unsigned(105,8) ,
2494	 => std_logic_vector(to_unsigned(109,8) ,
2495	 => std_logic_vector(to_unsigned(107,8) ,
2496	 => std_logic_vector(to_unsigned(104,8) ,
2497	 => std_logic_vector(to_unsigned(107,8) ,
2498	 => std_logic_vector(to_unsigned(104,8) ,
2499	 => std_logic_vector(to_unsigned(103,8) ,
2500	 => std_logic_vector(to_unsigned(109,8) ,
2501	 => std_logic_vector(to_unsigned(107,8) ,
2502	 => std_logic_vector(to_unsigned(109,8) ,
2503	 => std_logic_vector(to_unsigned(109,8) ,
2504	 => std_logic_vector(to_unsigned(101,8) ,
2505	 => std_logic_vector(to_unsigned(104,8) ,
2506	 => std_logic_vector(to_unsigned(104,8) ,
2507	 => std_logic_vector(to_unsigned(105,8) ,
2508	 => std_logic_vector(to_unsigned(112,8) ,
2509	 => std_logic_vector(to_unsigned(112,8) ,
2510	 => std_logic_vector(to_unsigned(111,8) ,
2511	 => std_logic_vector(to_unsigned(111,8) ,
2512	 => std_logic_vector(to_unsigned(108,8) ,
2513	 => std_logic_vector(to_unsigned(119,8) ,
2514	 => std_logic_vector(to_unsigned(130,8) ,
2515	 => std_logic_vector(to_unsigned(131,8) ,
2516	 => std_logic_vector(to_unsigned(133,8) ,
2517	 => std_logic_vector(to_unsigned(128,8) ,
2518	 => std_logic_vector(to_unsigned(125,8) ,
2519	 => std_logic_vector(to_unsigned(131,8) ,
2520	 => std_logic_vector(to_unsigned(138,8) ,
2521	 => std_logic_vector(to_unsigned(141,8) ,
2522	 => std_logic_vector(to_unsigned(141,8) ,
2523	 => std_logic_vector(to_unsigned(146,8) ,
2524	 => std_logic_vector(to_unsigned(146,8) ,
2525	 => std_logic_vector(to_unsigned(147,8) ,
2526	 => std_logic_vector(to_unsigned(147,8) ,
2527	 => std_logic_vector(to_unsigned(146,8) ,
2528	 => std_logic_vector(to_unsigned(146,8) ,
2529	 => std_logic_vector(to_unsigned(141,8) ,
2530	 => std_logic_vector(to_unsigned(146,8) ,
2531	 => std_logic_vector(to_unsigned(147,8) ,
2532	 => std_logic_vector(to_unsigned(151,8) ,
2533	 => std_logic_vector(to_unsigned(154,8) ,
2534	 => std_logic_vector(to_unsigned(154,8) ,
2535	 => std_logic_vector(to_unsigned(157,8) ,
2536	 => std_logic_vector(to_unsigned(159,8) ,
2537	 => std_logic_vector(to_unsigned(159,8) ,
2538	 => std_logic_vector(to_unsigned(161,8) ,
2539	 => std_logic_vector(to_unsigned(157,8) ,
2540	 => std_logic_vector(to_unsigned(157,8) ,
2541	 => std_logic_vector(to_unsigned(157,8) ,
2542	 => std_logic_vector(to_unsigned(159,8) ,
2543	 => std_logic_vector(to_unsigned(159,8) ,
2544	 => std_logic_vector(to_unsigned(157,8) ,
2545	 => std_logic_vector(to_unsigned(159,8) ,
2546	 => std_logic_vector(to_unsigned(161,8) ,
2547	 => std_logic_vector(to_unsigned(157,8) ,
2548	 => std_logic_vector(to_unsigned(159,8) ,
2549	 => std_logic_vector(to_unsigned(157,8) ,
2550	 => std_logic_vector(to_unsigned(156,8) ,
2551	 => std_logic_vector(to_unsigned(156,8) ,
2552	 => std_logic_vector(to_unsigned(157,8) ,
2553	 => std_logic_vector(to_unsigned(157,8) ,
2554	 => std_logic_vector(to_unsigned(161,8) ,
2555	 => std_logic_vector(to_unsigned(159,8) ,
2556	 => std_logic_vector(to_unsigned(159,8) ,
2557	 => std_logic_vector(to_unsigned(164,8) ,
2558	 => std_logic_vector(to_unsigned(163,8) ,
2559	 => std_logic_vector(to_unsigned(159,8) ,
2560	 => std_logic_vector(to_unsigned(163,8) ,
2561	 => std_logic_vector(to_unsigned(104,8) ,
2562	 => std_logic_vector(to_unsigned(103,8) ,
2563	 => std_logic_vector(to_unsigned(97,8) ,
2564	 => std_logic_vector(to_unsigned(90,8) ,
2565	 => std_logic_vector(to_unsigned(90,8) ,
2566	 => std_logic_vector(to_unsigned(90,8) ,
2567	 => std_logic_vector(to_unsigned(91,8) ,
2568	 => std_logic_vector(to_unsigned(91,8) ,
2569	 => std_logic_vector(to_unsigned(86,8) ,
2570	 => std_logic_vector(to_unsigned(90,8) ,
2571	 => std_logic_vector(to_unsigned(93,8) ,
2572	 => std_logic_vector(to_unsigned(88,8) ,
2573	 => std_logic_vector(to_unsigned(90,8) ,
2574	 => std_logic_vector(to_unsigned(96,8) ,
2575	 => std_logic_vector(to_unsigned(100,8) ,
2576	 => std_logic_vector(to_unsigned(85,8) ,
2577	 => std_logic_vector(to_unsigned(82,8) ,
2578	 => std_logic_vector(to_unsigned(87,8) ,
2579	 => std_logic_vector(to_unsigned(88,8) ,
2580	 => std_logic_vector(to_unsigned(87,8) ,
2581	 => std_logic_vector(to_unsigned(87,8) ,
2582	 => std_logic_vector(to_unsigned(91,8) ,
2583	 => std_logic_vector(to_unsigned(90,8) ,
2584	 => std_logic_vector(to_unsigned(88,8) ,
2585	 => std_logic_vector(to_unsigned(90,8) ,
2586	 => std_logic_vector(to_unsigned(88,8) ,
2587	 => std_logic_vector(to_unsigned(87,8) ,
2588	 => std_logic_vector(to_unsigned(90,8) ,
2589	 => std_logic_vector(to_unsigned(92,8) ,
2590	 => std_logic_vector(to_unsigned(91,8) ,
2591	 => std_logic_vector(to_unsigned(91,8) ,
2592	 => std_logic_vector(to_unsigned(93,8) ,
2593	 => std_logic_vector(to_unsigned(86,8) ,
2594	 => std_logic_vector(to_unsigned(87,8) ,
2595	 => std_logic_vector(to_unsigned(96,8) ,
2596	 => std_logic_vector(to_unsigned(99,8) ,
2597	 => std_logic_vector(to_unsigned(96,8) ,
2598	 => std_logic_vector(to_unsigned(95,8) ,
2599	 => std_logic_vector(to_unsigned(100,8) ,
2600	 => std_logic_vector(to_unsigned(99,8) ,
2601	 => std_logic_vector(to_unsigned(97,8) ,
2602	 => std_logic_vector(to_unsigned(103,8) ,
2603	 => std_logic_vector(to_unsigned(103,8) ,
2604	 => std_logic_vector(to_unsigned(100,8) ,
2605	 => std_logic_vector(to_unsigned(101,8) ,
2606	 => std_logic_vector(to_unsigned(99,8) ,
2607	 => std_logic_vector(to_unsigned(97,8) ,
2608	 => std_logic_vector(to_unsigned(104,8) ,
2609	 => std_logic_vector(to_unsigned(103,8) ,
2610	 => std_logic_vector(to_unsigned(99,8) ,
2611	 => std_logic_vector(to_unsigned(100,8) ,
2612	 => std_logic_vector(to_unsigned(103,8) ,
2613	 => std_logic_vector(to_unsigned(103,8) ,
2614	 => std_logic_vector(to_unsigned(103,8) ,
2615	 => std_logic_vector(to_unsigned(114,8) ,
2616	 => std_logic_vector(to_unsigned(111,8) ,
2617	 => std_logic_vector(to_unsigned(111,8) ,
2618	 => std_logic_vector(to_unsigned(112,8) ,
2619	 => std_logic_vector(to_unsigned(109,8) ,
2620	 => std_logic_vector(to_unsigned(108,8) ,
2621	 => std_logic_vector(to_unsigned(104,8) ,
2622	 => std_logic_vector(to_unsigned(107,8) ,
2623	 => std_logic_vector(to_unsigned(109,8) ,
2624	 => std_logic_vector(to_unsigned(101,8) ,
2625	 => std_logic_vector(to_unsigned(101,8) ,
2626	 => std_logic_vector(to_unsigned(107,8) ,
2627	 => std_logic_vector(to_unsigned(111,8) ,
2628	 => std_logic_vector(to_unsigned(111,8) ,
2629	 => std_logic_vector(to_unsigned(108,8) ,
2630	 => std_logic_vector(to_unsigned(107,8) ,
2631	 => std_logic_vector(to_unsigned(112,8) ,
2632	 => std_logic_vector(to_unsigned(116,8) ,
2633	 => std_logic_vector(to_unsigned(111,8) ,
2634	 => std_logic_vector(to_unsigned(112,8) ,
2635	 => std_logic_vector(to_unsigned(109,8) ,
2636	 => std_logic_vector(to_unsigned(109,8) ,
2637	 => std_logic_vector(to_unsigned(114,8) ,
2638	 => std_logic_vector(to_unsigned(108,8) ,
2639	 => std_logic_vector(to_unsigned(112,8) ,
2640	 => std_logic_vector(to_unsigned(112,8) ,
2641	 => std_logic_vector(to_unsigned(107,8) ,
2642	 => std_logic_vector(to_unsigned(103,8) ,
2643	 => std_logic_vector(to_unsigned(105,8) ,
2644	 => std_logic_vector(to_unsigned(104,8) ,
2645	 => std_logic_vector(to_unsigned(109,8) ,
2646	 => std_logic_vector(to_unsigned(108,8) ,
2647	 => std_logic_vector(to_unsigned(104,8) ,
2648	 => std_logic_vector(to_unsigned(108,8) ,
2649	 => std_logic_vector(to_unsigned(100,8) ,
2650	 => std_logic_vector(to_unsigned(100,8) ,
2651	 => std_logic_vector(to_unsigned(109,8) ,
2652	 => std_logic_vector(to_unsigned(108,8) ,
2653	 => std_logic_vector(to_unsigned(97,8) ,
2654	 => std_logic_vector(to_unsigned(93,8) ,
2655	 => std_logic_vector(to_unsigned(97,8) ,
2656	 => std_logic_vector(to_unsigned(100,8) ,
2657	 => std_logic_vector(to_unsigned(99,8) ,
2658	 => std_logic_vector(to_unsigned(97,8) ,
2659	 => std_logic_vector(to_unsigned(95,8) ,
2660	 => std_logic_vector(to_unsigned(92,8) ,
2661	 => std_logic_vector(to_unsigned(95,8) ,
2662	 => std_logic_vector(to_unsigned(101,8) ,
2663	 => std_logic_vector(to_unsigned(97,8) ,
2664	 => std_logic_vector(to_unsigned(93,8) ,
2665	 => std_logic_vector(to_unsigned(99,8) ,
2666	 => std_logic_vector(to_unsigned(101,8) ,
2667	 => std_logic_vector(to_unsigned(101,8) ,
2668	 => std_logic_vector(to_unsigned(108,8) ,
2669	 => std_logic_vector(to_unsigned(115,8) ,
2670	 => std_logic_vector(to_unsigned(105,8) ,
2671	 => std_logic_vector(to_unsigned(97,8) ,
2672	 => std_logic_vector(to_unsigned(105,8) ,
2673	 => std_logic_vector(to_unsigned(107,8) ,
2674	 => std_logic_vector(to_unsigned(108,8) ,
2675	 => std_logic_vector(to_unsigned(109,8) ,
2676	 => std_logic_vector(to_unsigned(103,8) ,
2677	 => std_logic_vector(to_unsigned(101,8) ,
2678	 => std_logic_vector(to_unsigned(104,8) ,
2679	 => std_logic_vector(to_unsigned(104,8) ,
2680	 => std_logic_vector(to_unsigned(105,8) ,
2681	 => std_logic_vector(to_unsigned(109,8) ,
2682	 => std_logic_vector(to_unsigned(105,8) ,
2683	 => std_logic_vector(to_unsigned(97,8) ,
2684	 => std_logic_vector(to_unsigned(97,8) ,
2685	 => std_logic_vector(to_unsigned(101,8) ,
2686	 => std_logic_vector(to_unsigned(100,8) ,
2687	 => std_logic_vector(to_unsigned(95,8) ,
2688	 => std_logic_vector(to_unsigned(91,8) ,
2689	 => std_logic_vector(to_unsigned(88,8) ,
2690	 => std_logic_vector(to_unsigned(92,8) ,
2691	 => std_logic_vector(to_unsigned(95,8) ,
2692	 => std_logic_vector(to_unsigned(92,8) ,
2693	 => std_logic_vector(to_unsigned(92,8) ,
2694	 => std_logic_vector(to_unsigned(96,8) ,
2695	 => std_logic_vector(to_unsigned(96,8) ,
2696	 => std_logic_vector(to_unsigned(95,8) ,
2697	 => std_logic_vector(to_unsigned(92,8) ,
2698	 => std_logic_vector(to_unsigned(92,8) ,
2699	 => std_logic_vector(to_unsigned(97,8) ,
2700	 => std_logic_vector(to_unsigned(104,8) ,
2701	 => std_logic_vector(to_unsigned(104,8) ,
2702	 => std_logic_vector(to_unsigned(105,8) ,
2703	 => std_logic_vector(to_unsigned(105,8) ,
2704	 => std_logic_vector(to_unsigned(104,8) ,
2705	 => std_logic_vector(to_unsigned(103,8) ,
2706	 => std_logic_vector(to_unsigned(101,8) ,
2707	 => std_logic_vector(to_unsigned(105,8) ,
2708	 => std_logic_vector(to_unsigned(105,8) ,
2709	 => std_logic_vector(to_unsigned(101,8) ,
2710	 => std_logic_vector(to_unsigned(104,8) ,
2711	 => std_logic_vector(to_unsigned(105,8) ,
2712	 => std_logic_vector(to_unsigned(100,8) ,
2713	 => std_logic_vector(to_unsigned(90,8) ,
2714	 => std_logic_vector(to_unsigned(87,8) ,
2715	 => std_logic_vector(to_unsigned(88,8) ,
2716	 => std_logic_vector(to_unsigned(86,8) ,
2717	 => std_logic_vector(to_unsigned(86,8) ,
2718	 => std_logic_vector(to_unsigned(90,8) ,
2719	 => std_logic_vector(to_unsigned(90,8) ,
2720	 => std_logic_vector(to_unsigned(86,8) ,
2721	 => std_logic_vector(to_unsigned(86,8) ,
2722	 => std_logic_vector(to_unsigned(82,8) ,
2723	 => std_logic_vector(to_unsigned(84,8) ,
2724	 => std_logic_vector(to_unsigned(84,8) ,
2725	 => std_logic_vector(to_unsigned(79,8) ,
2726	 => std_logic_vector(to_unsigned(81,8) ,
2727	 => std_logic_vector(to_unsigned(85,8) ,
2728	 => std_logic_vector(to_unsigned(91,8) ,
2729	 => std_logic_vector(to_unsigned(91,8) ,
2730	 => std_logic_vector(to_unsigned(86,8) ,
2731	 => std_logic_vector(to_unsigned(88,8) ,
2732	 => std_logic_vector(to_unsigned(97,8) ,
2733	 => std_logic_vector(to_unsigned(92,8) ,
2734	 => std_logic_vector(to_unsigned(85,8) ,
2735	 => std_logic_vector(to_unsigned(86,8) ,
2736	 => std_logic_vector(to_unsigned(85,8) ,
2737	 => std_logic_vector(to_unsigned(87,8) ,
2738	 => std_logic_vector(to_unsigned(86,8) ,
2739	 => std_logic_vector(to_unsigned(87,8) ,
2740	 => std_logic_vector(to_unsigned(80,8) ,
2741	 => std_logic_vector(to_unsigned(74,8) ,
2742	 => std_logic_vector(to_unsigned(76,8) ,
2743	 => std_logic_vector(to_unsigned(77,8) ,
2744	 => std_logic_vector(to_unsigned(74,8) ,
2745	 => std_logic_vector(to_unsigned(72,8) ,
2746	 => std_logic_vector(to_unsigned(77,8) ,
2747	 => std_logic_vector(to_unsigned(80,8) ,
2748	 => std_logic_vector(to_unsigned(80,8) ,
2749	 => std_logic_vector(to_unsigned(82,8) ,
2750	 => std_logic_vector(to_unsigned(79,8) ,
2751	 => std_logic_vector(to_unsigned(76,8) ,
2752	 => std_logic_vector(to_unsigned(70,8) ,
2753	 => std_logic_vector(to_unsigned(79,8) ,
2754	 => std_logic_vector(to_unsigned(78,8) ,
2755	 => std_logic_vector(to_unsigned(78,8) ,
2756	 => std_logic_vector(to_unsigned(84,8) ,
2757	 => std_logic_vector(to_unsigned(84,8) ,
2758	 => std_logic_vector(to_unsigned(84,8) ,
2759	 => std_logic_vector(to_unsigned(82,8) ,
2760	 => std_logic_vector(to_unsigned(80,8) ,
2761	 => std_logic_vector(to_unsigned(77,8) ,
2762	 => std_logic_vector(to_unsigned(78,8) ,
2763	 => std_logic_vector(to_unsigned(81,8) ,
2764	 => std_logic_vector(to_unsigned(81,8) ,
2765	 => std_logic_vector(to_unsigned(80,8) ,
2766	 => std_logic_vector(to_unsigned(80,8) ,
2767	 => std_logic_vector(to_unsigned(79,8) ,
2768	 => std_logic_vector(to_unsigned(78,8) ,
2769	 => std_logic_vector(to_unsigned(82,8) ,
2770	 => std_logic_vector(to_unsigned(85,8) ,
2771	 => std_logic_vector(to_unsigned(84,8) ,
2772	 => std_logic_vector(to_unsigned(78,8) ,
2773	 => std_logic_vector(to_unsigned(82,8) ,
2774	 => std_logic_vector(to_unsigned(86,8) ,
2775	 => std_logic_vector(to_unsigned(76,8) ,
2776	 => std_logic_vector(to_unsigned(72,8) ,
2777	 => std_logic_vector(to_unsigned(85,8) ,
2778	 => std_logic_vector(to_unsigned(86,8) ,
2779	 => std_logic_vector(to_unsigned(84,8) ,
2780	 => std_logic_vector(to_unsigned(82,8) ,
2781	 => std_logic_vector(to_unsigned(81,8) ,
2782	 => std_logic_vector(to_unsigned(85,8) ,
2783	 => std_logic_vector(to_unsigned(82,8) ,
2784	 => std_logic_vector(to_unsigned(79,8) ,
2785	 => std_logic_vector(to_unsigned(84,8) ,
2786	 => std_logic_vector(to_unsigned(88,8) ,
2787	 => std_logic_vector(to_unsigned(91,8) ,
2788	 => std_logic_vector(to_unsigned(92,8) ,
2789	 => std_logic_vector(to_unsigned(85,8) ,
2790	 => std_logic_vector(to_unsigned(86,8) ,
2791	 => std_logic_vector(to_unsigned(87,8) ,
2792	 => std_logic_vector(to_unsigned(87,8) ,
2793	 => std_logic_vector(to_unsigned(87,8) ,
2794	 => std_logic_vector(to_unsigned(84,8) ,
2795	 => std_logic_vector(to_unsigned(82,8) ,
2796	 => std_logic_vector(to_unsigned(81,8) ,
2797	 => std_logic_vector(to_unsigned(12,8) ,
2798	 => std_logic_vector(to_unsigned(0,8) ,
2799	 => std_logic_vector(to_unsigned(0,8) ,
2800	 => std_logic_vector(to_unsigned(9,8) ,
2801	 => std_logic_vector(to_unsigned(84,8) ,
2802	 => std_logic_vector(to_unsigned(84,8) ,
2803	 => std_logic_vector(to_unsigned(80,8) ,
2804	 => std_logic_vector(to_unsigned(91,8) ,
2805	 => std_logic_vector(to_unsigned(90,8) ,
2806	 => std_logic_vector(to_unsigned(90,8) ,
2807	 => std_logic_vector(to_unsigned(88,8) ,
2808	 => std_logic_vector(to_unsigned(91,8) ,
2809	 => std_logic_vector(to_unsigned(103,8) ,
2810	 => std_logic_vector(to_unsigned(111,8) ,
2811	 => std_logic_vector(to_unsigned(107,8) ,
2812	 => std_logic_vector(to_unsigned(105,8) ,
2813	 => std_logic_vector(to_unsigned(105,8) ,
2814	 => std_logic_vector(to_unsigned(104,8) ,
2815	 => std_logic_vector(to_unsigned(105,8) ,
2816	 => std_logic_vector(to_unsigned(103,8) ,
2817	 => std_logic_vector(to_unsigned(103,8) ,
2818	 => std_logic_vector(to_unsigned(100,8) ,
2819	 => std_logic_vector(to_unsigned(101,8) ,
2820	 => std_logic_vector(to_unsigned(108,8) ,
2821	 => std_logic_vector(to_unsigned(107,8) ,
2822	 => std_logic_vector(to_unsigned(108,8) ,
2823	 => std_logic_vector(to_unsigned(108,8) ,
2824	 => std_logic_vector(to_unsigned(103,8) ,
2825	 => std_logic_vector(to_unsigned(103,8) ,
2826	 => std_logic_vector(to_unsigned(107,8) ,
2827	 => std_logic_vector(to_unsigned(111,8) ,
2828	 => std_logic_vector(to_unsigned(105,8) ,
2829	 => std_logic_vector(to_unsigned(108,8) ,
2830	 => std_logic_vector(to_unsigned(111,8) ,
2831	 => std_logic_vector(to_unsigned(112,8) ,
2832	 => std_logic_vector(to_unsigned(112,8) ,
2833	 => std_logic_vector(to_unsigned(118,8) ,
2834	 => std_logic_vector(to_unsigned(127,8) ,
2835	 => std_logic_vector(to_unsigned(128,8) ,
2836	 => std_logic_vector(to_unsigned(130,8) ,
2837	 => std_logic_vector(to_unsigned(127,8) ,
2838	 => std_logic_vector(to_unsigned(128,8) ,
2839	 => std_logic_vector(to_unsigned(131,8) ,
2840	 => std_logic_vector(to_unsigned(136,8) ,
2841	 => std_logic_vector(to_unsigned(141,8) ,
2842	 => std_logic_vector(to_unsigned(142,8) ,
2843	 => std_logic_vector(to_unsigned(147,8) ,
2844	 => std_logic_vector(to_unsigned(142,8) ,
2845	 => std_logic_vector(to_unsigned(146,8) ,
2846	 => std_logic_vector(to_unsigned(151,8) ,
2847	 => std_logic_vector(to_unsigned(142,8) ,
2848	 => std_logic_vector(to_unsigned(139,8) ,
2849	 => std_logic_vector(to_unsigned(146,8) ,
2850	 => std_logic_vector(to_unsigned(149,8) ,
2851	 => std_logic_vector(to_unsigned(149,8) ,
2852	 => std_logic_vector(to_unsigned(152,8) ,
2853	 => std_logic_vector(to_unsigned(154,8) ,
2854	 => std_logic_vector(to_unsigned(154,8) ,
2855	 => std_logic_vector(to_unsigned(157,8) ,
2856	 => std_logic_vector(to_unsigned(156,8) ,
2857	 => std_logic_vector(to_unsigned(157,8) ,
2858	 => std_logic_vector(to_unsigned(159,8) ,
2859	 => std_logic_vector(to_unsigned(156,8) ,
2860	 => std_logic_vector(to_unsigned(154,8) ,
2861	 => std_logic_vector(to_unsigned(156,8) ,
2862	 => std_logic_vector(to_unsigned(157,8) ,
2863	 => std_logic_vector(to_unsigned(161,8) ,
2864	 => std_logic_vector(to_unsigned(161,8) ,
2865	 => std_logic_vector(to_unsigned(163,8) ,
2866	 => std_logic_vector(to_unsigned(163,8) ,
2867	 => std_logic_vector(to_unsigned(157,8) ,
2868	 => std_logic_vector(to_unsigned(156,8) ,
2869	 => std_logic_vector(to_unsigned(157,8) ,
2870	 => std_logic_vector(to_unsigned(159,8) ,
2871	 => std_logic_vector(to_unsigned(157,8) ,
2872	 => std_logic_vector(to_unsigned(157,8) ,
2873	 => std_logic_vector(to_unsigned(156,8) ,
2874	 => std_logic_vector(to_unsigned(157,8) ,
2875	 => std_logic_vector(to_unsigned(159,8) ,
2876	 => std_logic_vector(to_unsigned(159,8) ,
2877	 => std_logic_vector(to_unsigned(159,8) ,
2878	 => std_logic_vector(to_unsigned(159,8) ,
2879	 => std_logic_vector(to_unsigned(161,8) ,
2880	 => std_logic_vector(to_unsigned(159,8) ,
2881	 => std_logic_vector(to_unsigned(100,8) ,
2882	 => std_logic_vector(to_unsigned(93,8) ,
2883	 => std_logic_vector(to_unsigned(91,8) ,
2884	 => std_logic_vector(to_unsigned(95,8) ,
2885	 => std_logic_vector(to_unsigned(92,8) ,
2886	 => std_logic_vector(to_unsigned(87,8) ,
2887	 => std_logic_vector(to_unsigned(93,8) ,
2888	 => std_logic_vector(to_unsigned(93,8) ,
2889	 => std_logic_vector(to_unsigned(92,8) ,
2890	 => std_logic_vector(to_unsigned(95,8) ,
2891	 => std_logic_vector(to_unsigned(93,8) ,
2892	 => std_logic_vector(to_unsigned(90,8) ,
2893	 => std_logic_vector(to_unsigned(91,8) ,
2894	 => std_logic_vector(to_unsigned(95,8) ,
2895	 => std_logic_vector(to_unsigned(93,8) ,
2896	 => std_logic_vector(to_unsigned(86,8) ,
2897	 => std_logic_vector(to_unsigned(86,8) ,
2898	 => std_logic_vector(to_unsigned(87,8) ,
2899	 => std_logic_vector(to_unsigned(84,8) ,
2900	 => std_logic_vector(to_unsigned(86,8) ,
2901	 => std_logic_vector(to_unsigned(86,8) ,
2902	 => std_logic_vector(to_unsigned(86,8) ,
2903	 => std_logic_vector(to_unsigned(86,8) ,
2904	 => std_logic_vector(to_unsigned(86,8) ,
2905	 => std_logic_vector(to_unsigned(91,8) ,
2906	 => std_logic_vector(to_unsigned(91,8) ,
2907	 => std_logic_vector(to_unsigned(85,8) ,
2908	 => std_logic_vector(to_unsigned(88,8) ,
2909	 => std_logic_vector(to_unsigned(95,8) ,
2910	 => std_logic_vector(to_unsigned(95,8) ,
2911	 => std_logic_vector(to_unsigned(93,8) ,
2912	 => std_logic_vector(to_unsigned(85,8) ,
2913	 => std_logic_vector(to_unsigned(79,8) ,
2914	 => std_logic_vector(to_unsigned(87,8) ,
2915	 => std_logic_vector(to_unsigned(100,8) ,
2916	 => std_logic_vector(to_unsigned(96,8) ,
2917	 => std_logic_vector(to_unsigned(90,8) ,
2918	 => std_logic_vector(to_unsigned(91,8) ,
2919	 => std_logic_vector(to_unsigned(96,8) ,
2920	 => std_logic_vector(to_unsigned(95,8) ,
2921	 => std_logic_vector(to_unsigned(93,8) ,
2922	 => std_logic_vector(to_unsigned(99,8) ,
2923	 => std_logic_vector(to_unsigned(97,8) ,
2924	 => std_logic_vector(to_unsigned(96,8) ,
2925	 => std_logic_vector(to_unsigned(103,8) ,
2926	 => std_logic_vector(to_unsigned(104,8) ,
2927	 => std_logic_vector(to_unsigned(101,8) ,
2928	 => std_logic_vector(to_unsigned(101,8) ,
2929	 => std_logic_vector(to_unsigned(103,8) ,
2930	 => std_logic_vector(to_unsigned(104,8) ,
2931	 => std_logic_vector(to_unsigned(97,8) ,
2932	 => std_logic_vector(to_unsigned(100,8) ,
2933	 => std_logic_vector(to_unsigned(99,8) ,
2934	 => std_logic_vector(to_unsigned(100,8) ,
2935	 => std_logic_vector(to_unsigned(115,8) ,
2936	 => std_logic_vector(to_unsigned(111,8) ,
2937	 => std_logic_vector(to_unsigned(112,8) ,
2938	 => std_logic_vector(to_unsigned(115,8) ,
2939	 => std_logic_vector(to_unsigned(108,8) ,
2940	 => std_logic_vector(to_unsigned(108,8) ,
2941	 => std_logic_vector(to_unsigned(109,8) ,
2942	 => std_logic_vector(to_unsigned(108,8) ,
2943	 => std_logic_vector(to_unsigned(108,8) ,
2944	 => std_logic_vector(to_unsigned(103,8) ,
2945	 => std_logic_vector(to_unsigned(107,8) ,
2946	 => std_logic_vector(to_unsigned(111,8) ,
2947	 => std_logic_vector(to_unsigned(105,8) ,
2948	 => std_logic_vector(to_unsigned(107,8) ,
2949	 => std_logic_vector(to_unsigned(111,8) ,
2950	 => std_logic_vector(to_unsigned(107,8) ,
2951	 => std_logic_vector(to_unsigned(109,8) ,
2952	 => std_logic_vector(to_unsigned(116,8) ,
2953	 => std_logic_vector(to_unsigned(109,8) ,
2954	 => std_logic_vector(to_unsigned(112,8) ,
2955	 => std_logic_vector(to_unsigned(112,8) ,
2956	 => std_logic_vector(to_unsigned(114,8) ,
2957	 => std_logic_vector(to_unsigned(121,8) ,
2958	 => std_logic_vector(to_unsigned(112,8) ,
2959	 => std_logic_vector(to_unsigned(108,8) ,
2960	 => std_logic_vector(to_unsigned(105,8) ,
2961	 => std_logic_vector(to_unsigned(108,8) ,
2962	 => std_logic_vector(to_unsigned(103,8) ,
2963	 => std_logic_vector(to_unsigned(97,8) ,
2964	 => std_logic_vector(to_unsigned(101,8) ,
2965	 => std_logic_vector(to_unsigned(104,8) ,
2966	 => std_logic_vector(to_unsigned(103,8) ,
2967	 => std_logic_vector(to_unsigned(97,8) ,
2968	 => std_logic_vector(to_unsigned(99,8) ,
2969	 => std_logic_vector(to_unsigned(100,8) ,
2970	 => std_logic_vector(to_unsigned(97,8) ,
2971	 => std_logic_vector(to_unsigned(111,8) ,
2972	 => std_logic_vector(to_unsigned(104,8) ,
2973	 => std_logic_vector(to_unsigned(97,8) ,
2974	 => std_logic_vector(to_unsigned(99,8) ,
2975	 => std_logic_vector(to_unsigned(99,8) ,
2976	 => std_logic_vector(to_unsigned(95,8) ,
2977	 => std_logic_vector(to_unsigned(93,8) ,
2978	 => std_logic_vector(to_unsigned(96,8) ,
2979	 => std_logic_vector(to_unsigned(99,8) ,
2980	 => std_logic_vector(to_unsigned(97,8) ,
2981	 => std_logic_vector(to_unsigned(96,8) ,
2982	 => std_logic_vector(to_unsigned(97,8) ,
2983	 => std_logic_vector(to_unsigned(93,8) ,
2984	 => std_logic_vector(to_unsigned(93,8) ,
2985	 => std_logic_vector(to_unsigned(97,8) ,
2986	 => std_logic_vector(to_unsigned(97,8) ,
2987	 => std_logic_vector(to_unsigned(97,8) ,
2988	 => std_logic_vector(to_unsigned(97,8) ,
2989	 => std_logic_vector(to_unsigned(104,8) ,
2990	 => std_logic_vector(to_unsigned(103,8) ,
2991	 => std_logic_vector(to_unsigned(95,8) ,
2992	 => std_logic_vector(to_unsigned(97,8) ,
2993	 => std_logic_vector(to_unsigned(101,8) ,
2994	 => std_logic_vector(to_unsigned(103,8) ,
2995	 => std_logic_vector(to_unsigned(101,8) ,
2996	 => std_logic_vector(to_unsigned(95,8) ,
2997	 => std_logic_vector(to_unsigned(95,8) ,
2998	 => std_logic_vector(to_unsigned(101,8) ,
2999	 => std_logic_vector(to_unsigned(105,8) ,
3000	 => std_logic_vector(to_unsigned(104,8) ,
3001	 => std_logic_vector(to_unsigned(107,8) ,
3002	 => std_logic_vector(to_unsigned(104,8) ,
3003	 => std_logic_vector(to_unsigned(100,8) ,
3004	 => std_logic_vector(to_unsigned(100,8) ,
3005	 => std_logic_vector(to_unsigned(100,8) ,
3006	 => std_logic_vector(to_unsigned(100,8) ,
3007	 => std_logic_vector(to_unsigned(100,8) ,
3008	 => std_logic_vector(to_unsigned(99,8) ,
3009	 => std_logic_vector(to_unsigned(95,8) ,
3010	 => std_logic_vector(to_unsigned(95,8) ,
3011	 => std_logic_vector(to_unsigned(97,8) ,
3012	 => std_logic_vector(to_unsigned(93,8) ,
3013	 => std_logic_vector(to_unsigned(96,8) ,
3014	 => std_logic_vector(to_unsigned(99,8) ,
3015	 => std_logic_vector(to_unsigned(96,8) ,
3016	 => std_logic_vector(to_unsigned(96,8) ,
3017	 => std_logic_vector(to_unsigned(91,8) ,
3018	 => std_logic_vector(to_unsigned(96,8) ,
3019	 => std_logic_vector(to_unsigned(99,8) ,
3020	 => std_logic_vector(to_unsigned(96,8) ,
3021	 => std_logic_vector(to_unsigned(99,8) ,
3022	 => std_logic_vector(to_unsigned(105,8) ,
3023	 => std_logic_vector(to_unsigned(107,8) ,
3024	 => std_logic_vector(to_unsigned(104,8) ,
3025	 => std_logic_vector(to_unsigned(100,8) ,
3026	 => std_logic_vector(to_unsigned(95,8) ,
3027	 => std_logic_vector(to_unsigned(99,8) ,
3028	 => std_logic_vector(to_unsigned(101,8) ,
3029	 => std_logic_vector(to_unsigned(96,8) ,
3030	 => std_logic_vector(to_unsigned(97,8) ,
3031	 => std_logic_vector(to_unsigned(95,8) ,
3032	 => std_logic_vector(to_unsigned(90,8) ,
3033	 => std_logic_vector(to_unsigned(88,8) ,
3034	 => std_logic_vector(to_unsigned(84,8) ,
3035	 => std_logic_vector(to_unsigned(84,8) ,
3036	 => std_logic_vector(to_unsigned(80,8) ,
3037	 => std_logic_vector(to_unsigned(82,8) ,
3038	 => std_logic_vector(to_unsigned(81,8) ,
3039	 => std_logic_vector(to_unsigned(84,8) ,
3040	 => std_logic_vector(to_unsigned(81,8) ,
3041	 => std_logic_vector(to_unsigned(81,8) ,
3042	 => std_logic_vector(to_unsigned(79,8) ,
3043	 => std_logic_vector(to_unsigned(80,8) ,
3044	 => std_logic_vector(to_unsigned(84,8) ,
3045	 => std_logic_vector(to_unsigned(82,8) ,
3046	 => std_logic_vector(to_unsigned(82,8) ,
3047	 => std_logic_vector(to_unsigned(79,8) ,
3048	 => std_logic_vector(to_unsigned(79,8) ,
3049	 => std_logic_vector(to_unsigned(82,8) ,
3050	 => std_logic_vector(to_unsigned(86,8) ,
3051	 => std_logic_vector(to_unsigned(87,8) ,
3052	 => std_logic_vector(to_unsigned(87,8) ,
3053	 => std_logic_vector(to_unsigned(87,8) ,
3054	 => std_logic_vector(to_unsigned(86,8) ,
3055	 => std_logic_vector(to_unsigned(86,8) ,
3056	 => std_logic_vector(to_unsigned(85,8) ,
3057	 => std_logic_vector(to_unsigned(86,8) ,
3058	 => std_logic_vector(to_unsigned(82,8) ,
3059	 => std_logic_vector(to_unsigned(80,8) ,
3060	 => std_logic_vector(to_unsigned(78,8) ,
3061	 => std_logic_vector(to_unsigned(70,8) ,
3062	 => std_logic_vector(to_unsigned(71,8) ,
3063	 => std_logic_vector(to_unsigned(79,8) ,
3064	 => std_logic_vector(to_unsigned(78,8) ,
3065	 => std_logic_vector(to_unsigned(72,8) ,
3066	 => std_logic_vector(to_unsigned(74,8) ,
3067	 => std_logic_vector(to_unsigned(77,8) ,
3068	 => std_logic_vector(to_unsigned(77,8) ,
3069	 => std_logic_vector(to_unsigned(77,8) ,
3070	 => std_logic_vector(to_unsigned(67,8) ,
3071	 => std_logic_vector(to_unsigned(73,8) ,
3072	 => std_logic_vector(to_unsigned(73,8) ,
3073	 => std_logic_vector(to_unsigned(76,8) ,
3074	 => std_logic_vector(to_unsigned(74,8) ,
3075	 => std_logic_vector(to_unsigned(77,8) ,
3076	 => std_logic_vector(to_unsigned(78,8) ,
3077	 => std_logic_vector(to_unsigned(72,8) ,
3078	 => std_logic_vector(to_unsigned(78,8) ,
3079	 => std_logic_vector(to_unsigned(77,8) ,
3080	 => std_logic_vector(to_unsigned(77,8) ,
3081	 => std_logic_vector(to_unsigned(78,8) ,
3082	 => std_logic_vector(to_unsigned(74,8) ,
3083	 => std_logic_vector(to_unsigned(80,8) ,
3084	 => std_logic_vector(to_unsigned(80,8) ,
3085	 => std_logic_vector(to_unsigned(74,8) ,
3086	 => std_logic_vector(to_unsigned(72,8) ,
3087	 => std_logic_vector(to_unsigned(76,8) ,
3088	 => std_logic_vector(to_unsigned(79,8) ,
3089	 => std_logic_vector(to_unsigned(82,8) ,
3090	 => std_logic_vector(to_unsigned(87,8) ,
3091	 => std_logic_vector(to_unsigned(87,8) ,
3092	 => std_logic_vector(to_unsigned(81,8) ,
3093	 => std_logic_vector(to_unsigned(81,8) ,
3094	 => std_logic_vector(to_unsigned(82,8) ,
3095	 => std_logic_vector(to_unsigned(84,8) ,
3096	 => std_logic_vector(to_unsigned(81,8) ,
3097	 => std_logic_vector(to_unsigned(77,8) ,
3098	 => std_logic_vector(to_unsigned(82,8) ,
3099	 => std_logic_vector(to_unsigned(84,8) ,
3100	 => std_logic_vector(to_unsigned(81,8) ,
3101	 => std_logic_vector(to_unsigned(82,8) ,
3102	 => std_logic_vector(to_unsigned(81,8) ,
3103	 => std_logic_vector(to_unsigned(85,8) ,
3104	 => std_logic_vector(to_unsigned(86,8) ,
3105	 => std_logic_vector(to_unsigned(86,8) ,
3106	 => std_logic_vector(to_unsigned(84,8) ,
3107	 => std_logic_vector(to_unsigned(86,8) ,
3108	 => std_logic_vector(to_unsigned(87,8) ,
3109	 => std_logic_vector(to_unsigned(85,8) ,
3110	 => std_logic_vector(to_unsigned(85,8) ,
3111	 => std_logic_vector(to_unsigned(87,8) ,
3112	 => std_logic_vector(to_unsigned(91,8) ,
3113	 => std_logic_vector(to_unsigned(86,8) ,
3114	 => std_logic_vector(to_unsigned(84,8) ,
3115	 => std_logic_vector(to_unsigned(80,8) ,
3116	 => std_logic_vector(to_unsigned(81,8) ,
3117	 => std_logic_vector(to_unsigned(29,8) ,
3118	 => std_logic_vector(to_unsigned(1,8) ,
3119	 => std_logic_vector(to_unsigned(0,8) ,
3120	 => std_logic_vector(to_unsigned(2,8) ,
3121	 => std_logic_vector(to_unsigned(59,8) ,
3122	 => std_logic_vector(to_unsigned(88,8) ,
3123	 => std_logic_vector(to_unsigned(81,8) ,
3124	 => std_logic_vector(to_unsigned(85,8) ,
3125	 => std_logic_vector(to_unsigned(90,8) ,
3126	 => std_logic_vector(to_unsigned(92,8) ,
3127	 => std_logic_vector(to_unsigned(90,8) ,
3128	 => std_logic_vector(to_unsigned(95,8) ,
3129	 => std_logic_vector(to_unsigned(101,8) ,
3130	 => std_logic_vector(to_unsigned(118,8) ,
3131	 => std_logic_vector(to_unsigned(130,8) ,
3132	 => std_logic_vector(to_unsigned(122,8) ,
3133	 => std_logic_vector(to_unsigned(107,8) ,
3134	 => std_logic_vector(to_unsigned(97,8) ,
3135	 => std_logic_vector(to_unsigned(101,8) ,
3136	 => std_logic_vector(to_unsigned(101,8) ,
3137	 => std_logic_vector(to_unsigned(99,8) ,
3138	 => std_logic_vector(to_unsigned(97,8) ,
3139	 => std_logic_vector(to_unsigned(103,8) ,
3140	 => std_logic_vector(to_unsigned(111,8) ,
3141	 => std_logic_vector(to_unsigned(105,8) ,
3142	 => std_logic_vector(to_unsigned(101,8) ,
3143	 => std_logic_vector(to_unsigned(100,8) ,
3144	 => std_logic_vector(to_unsigned(93,8) ,
3145	 => std_logic_vector(to_unsigned(103,8) ,
3146	 => std_logic_vector(to_unsigned(109,8) ,
3147	 => std_logic_vector(to_unsigned(109,8) ,
3148	 => std_logic_vector(to_unsigned(107,8) ,
3149	 => std_logic_vector(to_unsigned(108,8) ,
3150	 => std_logic_vector(to_unsigned(109,8) ,
3151	 => std_logic_vector(to_unsigned(112,8) ,
3152	 => std_logic_vector(to_unsigned(115,8) ,
3153	 => std_logic_vector(to_unsigned(114,8) ,
3154	 => std_logic_vector(to_unsigned(121,8) ,
3155	 => std_logic_vector(to_unsigned(128,8) ,
3156	 => std_logic_vector(to_unsigned(128,8) ,
3157	 => std_logic_vector(to_unsigned(127,8) ,
3158	 => std_logic_vector(to_unsigned(133,8) ,
3159	 => std_logic_vector(to_unsigned(136,8) ,
3160	 => std_logic_vector(to_unsigned(136,8) ,
3161	 => std_logic_vector(to_unsigned(134,8) ,
3162	 => std_logic_vector(to_unsigned(136,8) ,
3163	 => std_logic_vector(to_unsigned(136,8) ,
3164	 => std_logic_vector(to_unsigned(141,8) ,
3165	 => std_logic_vector(to_unsigned(144,8) ,
3166	 => std_logic_vector(to_unsigned(146,8) ,
3167	 => std_logic_vector(to_unsigned(144,8) ,
3168	 => std_logic_vector(to_unsigned(141,8) ,
3169	 => std_logic_vector(to_unsigned(152,8) ,
3170	 => std_logic_vector(to_unsigned(157,8) ,
3171	 => std_logic_vector(to_unsigned(151,8) ,
3172	 => std_logic_vector(to_unsigned(149,8) ,
3173	 => std_logic_vector(to_unsigned(151,8) ,
3174	 => std_logic_vector(to_unsigned(154,8) ,
3175	 => std_logic_vector(to_unsigned(154,8) ,
3176	 => std_logic_vector(to_unsigned(156,8) ,
3177	 => std_logic_vector(to_unsigned(159,8) ,
3178	 => std_logic_vector(to_unsigned(159,8) ,
3179	 => std_logic_vector(to_unsigned(156,8) ,
3180	 => std_logic_vector(to_unsigned(156,8) ,
3181	 => std_logic_vector(to_unsigned(157,8) ,
3182	 => std_logic_vector(to_unsigned(159,8) ,
3183	 => std_logic_vector(to_unsigned(161,8) ,
3184	 => std_logic_vector(to_unsigned(159,8) ,
3185	 => std_logic_vector(to_unsigned(161,8) ,
3186	 => std_logic_vector(to_unsigned(161,8) ,
3187	 => std_logic_vector(to_unsigned(159,8) ,
3188	 => std_logic_vector(to_unsigned(159,8) ,
3189	 => std_logic_vector(to_unsigned(159,8) ,
3190	 => std_logic_vector(to_unsigned(161,8) ,
3191	 => std_logic_vector(to_unsigned(161,8) ,
3192	 => std_logic_vector(to_unsigned(159,8) ,
3193	 => std_logic_vector(to_unsigned(157,8) ,
3194	 => std_logic_vector(to_unsigned(157,8) ,
3195	 => std_logic_vector(to_unsigned(159,8) ,
3196	 => std_logic_vector(to_unsigned(161,8) ,
3197	 => std_logic_vector(to_unsigned(161,8) ,
3198	 => std_logic_vector(to_unsigned(163,8) ,
3199	 => std_logic_vector(to_unsigned(163,8) ,
3200	 => std_logic_vector(to_unsigned(163,8) ,
3201	 => std_logic_vector(to_unsigned(95,8) ,
3202	 => std_logic_vector(to_unsigned(96,8) ,
3203	 => std_logic_vector(to_unsigned(91,8) ,
3204	 => std_logic_vector(to_unsigned(91,8) ,
3205	 => std_logic_vector(to_unsigned(91,8) ,
3206	 => std_logic_vector(to_unsigned(90,8) ,
3207	 => std_logic_vector(to_unsigned(91,8) ,
3208	 => std_logic_vector(to_unsigned(87,8) ,
3209	 => std_logic_vector(to_unsigned(90,8) ,
3210	 => std_logic_vector(to_unsigned(92,8) ,
3211	 => std_logic_vector(to_unsigned(86,8) ,
3212	 => std_logic_vector(to_unsigned(82,8) ,
3213	 => std_logic_vector(to_unsigned(86,8) ,
3214	 => std_logic_vector(to_unsigned(86,8) ,
3215	 => std_logic_vector(to_unsigned(85,8) ,
3216	 => std_logic_vector(to_unsigned(85,8) ,
3217	 => std_logic_vector(to_unsigned(90,8) ,
3218	 => std_logic_vector(to_unsigned(85,8) ,
3219	 => std_logic_vector(to_unsigned(82,8) ,
3220	 => std_logic_vector(to_unsigned(85,8) ,
3221	 => std_logic_vector(to_unsigned(85,8) ,
3222	 => std_logic_vector(to_unsigned(86,8) ,
3223	 => std_logic_vector(to_unsigned(86,8) ,
3224	 => std_logic_vector(to_unsigned(84,8) ,
3225	 => std_logic_vector(to_unsigned(85,8) ,
3226	 => std_logic_vector(to_unsigned(84,8) ,
3227	 => std_logic_vector(to_unsigned(81,8) ,
3228	 => std_logic_vector(to_unsigned(86,8) ,
3229	 => std_logic_vector(to_unsigned(92,8) ,
3230	 => std_logic_vector(to_unsigned(88,8) ,
3231	 => std_logic_vector(to_unsigned(87,8) ,
3232	 => std_logic_vector(to_unsigned(86,8) ,
3233	 => std_logic_vector(to_unsigned(82,8) ,
3234	 => std_logic_vector(to_unsigned(86,8) ,
3235	 => std_logic_vector(to_unsigned(91,8) ,
3236	 => std_logic_vector(to_unsigned(88,8) ,
3237	 => std_logic_vector(to_unsigned(92,8) ,
3238	 => std_logic_vector(to_unsigned(91,8) ,
3239	 => std_logic_vector(to_unsigned(91,8) ,
3240	 => std_logic_vector(to_unsigned(92,8) ,
3241	 => std_logic_vector(to_unsigned(95,8) ,
3242	 => std_logic_vector(to_unsigned(96,8) ,
3243	 => std_logic_vector(to_unsigned(93,8) ,
3244	 => std_logic_vector(to_unsigned(96,8) ,
3245	 => std_logic_vector(to_unsigned(103,8) ,
3246	 => std_logic_vector(to_unsigned(107,8) ,
3247	 => std_logic_vector(to_unsigned(105,8) ,
3248	 => std_logic_vector(to_unsigned(103,8) ,
3249	 => std_logic_vector(to_unsigned(103,8) ,
3250	 => std_logic_vector(to_unsigned(107,8) ,
3251	 => std_logic_vector(to_unsigned(100,8) ,
3252	 => std_logic_vector(to_unsigned(99,8) ,
3253	 => std_logic_vector(to_unsigned(97,8) ,
3254	 => std_logic_vector(to_unsigned(101,8) ,
3255	 => std_logic_vector(to_unsigned(104,8) ,
3256	 => std_logic_vector(to_unsigned(105,8) ,
3257	 => std_logic_vector(to_unsigned(108,8) ,
3258	 => std_logic_vector(to_unsigned(112,8) ,
3259	 => std_logic_vector(to_unsigned(109,8) ,
3260	 => std_logic_vector(to_unsigned(107,8) ,
3261	 => std_logic_vector(to_unsigned(105,8) ,
3262	 => std_logic_vector(to_unsigned(107,8) ,
3263	 => std_logic_vector(to_unsigned(108,8) ,
3264	 => std_logic_vector(to_unsigned(105,8) ,
3265	 => std_logic_vector(to_unsigned(109,8) ,
3266	 => std_logic_vector(to_unsigned(105,8) ,
3267	 => std_logic_vector(to_unsigned(96,8) ,
3268	 => std_logic_vector(to_unsigned(103,8) ,
3269	 => std_logic_vector(to_unsigned(112,8) ,
3270	 => std_logic_vector(to_unsigned(107,8) ,
3271	 => std_logic_vector(to_unsigned(109,8) ,
3272	 => std_logic_vector(to_unsigned(112,8) ,
3273	 => std_logic_vector(to_unsigned(108,8) ,
3274	 => std_logic_vector(to_unsigned(112,8) ,
3275	 => std_logic_vector(to_unsigned(109,8) ,
3276	 => std_logic_vector(to_unsigned(109,8) ,
3277	 => std_logic_vector(to_unsigned(116,8) ,
3278	 => std_logic_vector(to_unsigned(111,8) ,
3279	 => std_logic_vector(to_unsigned(105,8) ,
3280	 => std_logic_vector(to_unsigned(105,8) ,
3281	 => std_logic_vector(to_unsigned(109,8) ,
3282	 => std_logic_vector(to_unsigned(104,8) ,
3283	 => std_logic_vector(to_unsigned(97,8) ,
3284	 => std_logic_vector(to_unsigned(101,8) ,
3285	 => std_logic_vector(to_unsigned(100,8) ,
3286	 => std_logic_vector(to_unsigned(100,8) ,
3287	 => std_logic_vector(to_unsigned(95,8) ,
3288	 => std_logic_vector(to_unsigned(92,8) ,
3289	 => std_logic_vector(to_unsigned(99,8) ,
3290	 => std_logic_vector(to_unsigned(96,8) ,
3291	 => std_logic_vector(to_unsigned(103,8) ,
3292	 => std_logic_vector(to_unsigned(97,8) ,
3293	 => std_logic_vector(to_unsigned(99,8) ,
3294	 => std_logic_vector(to_unsigned(100,8) ,
3295	 => std_logic_vector(to_unsigned(95,8) ,
3296	 => std_logic_vector(to_unsigned(91,8) ,
3297	 => std_logic_vector(to_unsigned(91,8) ,
3298	 => std_logic_vector(to_unsigned(93,8) ,
3299	 => std_logic_vector(to_unsigned(93,8) ,
3300	 => std_logic_vector(to_unsigned(88,8) ,
3301	 => std_logic_vector(to_unsigned(86,8) ,
3302	 => std_logic_vector(to_unsigned(91,8) ,
3303	 => std_logic_vector(to_unsigned(92,8) ,
3304	 => std_logic_vector(to_unsigned(92,8) ,
3305	 => std_logic_vector(to_unsigned(93,8) ,
3306	 => std_logic_vector(to_unsigned(93,8) ,
3307	 => std_logic_vector(to_unsigned(97,8) ,
3308	 => std_logic_vector(to_unsigned(95,8) ,
3309	 => std_logic_vector(to_unsigned(99,8) ,
3310	 => std_logic_vector(to_unsigned(101,8) ,
3311	 => std_logic_vector(to_unsigned(96,8) ,
3312	 => std_logic_vector(to_unsigned(97,8) ,
3313	 => std_logic_vector(to_unsigned(97,8) ,
3314	 => std_logic_vector(to_unsigned(93,8) ,
3315	 => std_logic_vector(to_unsigned(97,8) ,
3316	 => std_logic_vector(to_unsigned(92,8) ,
3317	 => std_logic_vector(to_unsigned(92,8) ,
3318	 => std_logic_vector(to_unsigned(93,8) ,
3319	 => std_logic_vector(to_unsigned(95,8) ,
3320	 => std_logic_vector(to_unsigned(97,8) ,
3321	 => std_logic_vector(to_unsigned(97,8) ,
3322	 => std_logic_vector(to_unsigned(101,8) ,
3323	 => std_logic_vector(to_unsigned(100,8) ,
3324	 => std_logic_vector(to_unsigned(97,8) ,
3325	 => std_logic_vector(to_unsigned(97,8) ,
3326	 => std_logic_vector(to_unsigned(99,8) ,
3327	 => std_logic_vector(to_unsigned(91,8) ,
3328	 => std_logic_vector(to_unsigned(92,8) ,
3329	 => std_logic_vector(to_unsigned(96,8) ,
3330	 => std_logic_vector(to_unsigned(95,8) ,
3331	 => std_logic_vector(to_unsigned(93,8) ,
3332	 => std_logic_vector(to_unsigned(90,8) ,
3333	 => std_logic_vector(to_unsigned(92,8) ,
3334	 => std_logic_vector(to_unsigned(91,8) ,
3335	 => std_logic_vector(to_unsigned(90,8) ,
3336	 => std_logic_vector(to_unsigned(93,8) ,
3337	 => std_logic_vector(to_unsigned(96,8) ,
3338	 => std_logic_vector(to_unsigned(99,8) ,
3339	 => std_logic_vector(to_unsigned(96,8) ,
3340	 => std_logic_vector(to_unsigned(91,8) ,
3341	 => std_logic_vector(to_unsigned(96,8) ,
3342	 => std_logic_vector(to_unsigned(103,8) ,
3343	 => std_logic_vector(to_unsigned(97,8) ,
3344	 => std_logic_vector(to_unsigned(99,8) ,
3345	 => std_logic_vector(to_unsigned(101,8) ,
3346	 => std_logic_vector(to_unsigned(99,8) ,
3347	 => std_logic_vector(to_unsigned(95,8) ,
3348	 => std_logic_vector(to_unsigned(91,8) ,
3349	 => std_logic_vector(to_unsigned(92,8) ,
3350	 => std_logic_vector(to_unsigned(91,8) ,
3351	 => std_logic_vector(to_unsigned(86,8) ,
3352	 => std_logic_vector(to_unsigned(86,8) ,
3353	 => std_logic_vector(to_unsigned(86,8) ,
3354	 => std_logic_vector(to_unsigned(76,8) ,
3355	 => std_logic_vector(to_unsigned(74,8) ,
3356	 => std_logic_vector(to_unsigned(81,8) ,
3357	 => std_logic_vector(to_unsigned(84,8) ,
3358	 => std_logic_vector(to_unsigned(80,8) ,
3359	 => std_logic_vector(to_unsigned(82,8) ,
3360	 => std_logic_vector(to_unsigned(85,8) ,
3361	 => std_logic_vector(to_unsigned(86,8) ,
3362	 => std_logic_vector(to_unsigned(84,8) ,
3363	 => std_logic_vector(to_unsigned(84,8) ,
3364	 => std_logic_vector(to_unsigned(86,8) ,
3365	 => std_logic_vector(to_unsigned(88,8) ,
3366	 => std_logic_vector(to_unsigned(90,8) ,
3367	 => std_logic_vector(to_unsigned(85,8) ,
3368	 => std_logic_vector(to_unsigned(82,8) ,
3369	 => std_logic_vector(to_unsigned(84,8) ,
3370	 => std_logic_vector(to_unsigned(88,8) ,
3371	 => std_logic_vector(to_unsigned(85,8) ,
3372	 => std_logic_vector(to_unsigned(86,8) ,
3373	 => std_logic_vector(to_unsigned(90,8) ,
3374	 => std_logic_vector(to_unsigned(88,8) ,
3375	 => std_logic_vector(to_unsigned(85,8) ,
3376	 => std_logic_vector(to_unsigned(85,8) ,
3377	 => std_logic_vector(to_unsigned(87,8) ,
3378	 => std_logic_vector(to_unsigned(82,8) ,
3379	 => std_logic_vector(to_unsigned(76,8) ,
3380	 => std_logic_vector(to_unsigned(77,8) ,
3381	 => std_logic_vector(to_unsigned(72,8) ,
3382	 => std_logic_vector(to_unsigned(71,8) ,
3383	 => std_logic_vector(to_unsigned(76,8) ,
3384	 => std_logic_vector(to_unsigned(77,8) ,
3385	 => std_logic_vector(to_unsigned(73,8) ,
3386	 => std_logic_vector(to_unsigned(72,8) ,
3387	 => std_logic_vector(to_unsigned(68,8) ,
3388	 => std_logic_vector(to_unsigned(71,8) ,
3389	 => std_logic_vector(to_unsigned(76,8) ,
3390	 => std_logic_vector(to_unsigned(69,8) ,
3391	 => std_logic_vector(to_unsigned(73,8) ,
3392	 => std_logic_vector(to_unsigned(73,8) ,
3393	 => std_logic_vector(to_unsigned(79,8) ,
3394	 => std_logic_vector(to_unsigned(84,8) ,
3395	 => std_logic_vector(to_unsigned(76,8) ,
3396	 => std_logic_vector(to_unsigned(70,8) ,
3397	 => std_logic_vector(to_unsigned(70,8) ,
3398	 => std_logic_vector(to_unsigned(79,8) ,
3399	 => std_logic_vector(to_unsigned(73,8) ,
3400	 => std_logic_vector(to_unsigned(72,8) ,
3401	 => std_logic_vector(to_unsigned(79,8) ,
3402	 => std_logic_vector(to_unsigned(76,8) ,
3403	 => std_logic_vector(to_unsigned(77,8) ,
3404	 => std_logic_vector(to_unsigned(73,8) ,
3405	 => std_logic_vector(to_unsigned(78,8) ,
3406	 => std_logic_vector(to_unsigned(80,8) ,
3407	 => std_logic_vector(to_unsigned(78,8) ,
3408	 => std_logic_vector(to_unsigned(80,8) ,
3409	 => std_logic_vector(to_unsigned(87,8) ,
3410	 => std_logic_vector(to_unsigned(85,8) ,
3411	 => std_logic_vector(to_unsigned(80,8) ,
3412	 => std_logic_vector(to_unsigned(84,8) ,
3413	 => std_logic_vector(to_unsigned(82,8) ,
3414	 => std_logic_vector(to_unsigned(78,8) ,
3415	 => std_logic_vector(to_unsigned(82,8) ,
3416	 => std_logic_vector(to_unsigned(81,8) ,
3417	 => std_logic_vector(to_unsigned(74,8) ,
3418	 => std_logic_vector(to_unsigned(82,8) ,
3419	 => std_logic_vector(to_unsigned(84,8) ,
3420	 => std_logic_vector(to_unsigned(84,8) ,
3421	 => std_logic_vector(to_unsigned(90,8) ,
3422	 => std_logic_vector(to_unsigned(86,8) ,
3423	 => std_logic_vector(to_unsigned(85,8) ,
3424	 => std_logic_vector(to_unsigned(90,8) ,
3425	 => std_logic_vector(to_unsigned(88,8) ,
3426	 => std_logic_vector(to_unsigned(86,8) ,
3427	 => std_logic_vector(to_unsigned(87,8) ,
3428	 => std_logic_vector(to_unsigned(86,8) ,
3429	 => std_logic_vector(to_unsigned(88,8) ,
3430	 => std_logic_vector(to_unsigned(88,8) ,
3431	 => std_logic_vector(to_unsigned(84,8) ,
3432	 => std_logic_vector(to_unsigned(88,8) ,
3433	 => std_logic_vector(to_unsigned(85,8) ,
3434	 => std_logic_vector(to_unsigned(85,8) ,
3435	 => std_logic_vector(to_unsigned(81,8) ,
3436	 => std_logic_vector(to_unsigned(85,8) ,
3437	 => std_logic_vector(to_unsigned(58,8) ,
3438	 => std_logic_vector(to_unsigned(2,8) ,
3439	 => std_logic_vector(to_unsigned(0,8) ,
3440	 => std_logic_vector(to_unsigned(0,8) ,
3441	 => std_logic_vector(to_unsigned(39,8) ,
3442	 => std_logic_vector(to_unsigned(103,8) ,
3443	 => std_logic_vector(to_unsigned(91,8) ,
3444	 => std_logic_vector(to_unsigned(87,8) ,
3445	 => std_logic_vector(to_unsigned(92,8) ,
3446	 => std_logic_vector(to_unsigned(99,8) ,
3447	 => std_logic_vector(to_unsigned(96,8) ,
3448	 => std_logic_vector(to_unsigned(93,8) ,
3449	 => std_logic_vector(to_unsigned(96,8) ,
3450	 => std_logic_vector(to_unsigned(105,8) ,
3451	 => std_logic_vector(to_unsigned(131,8) ,
3452	 => std_logic_vector(to_unsigned(131,8) ,
3453	 => std_logic_vector(to_unsigned(109,8) ,
3454	 => std_logic_vector(to_unsigned(104,8) ,
3455	 => std_logic_vector(to_unsigned(109,8) ,
3456	 => std_logic_vector(to_unsigned(100,8) ,
3457	 => std_logic_vector(to_unsigned(97,8) ,
3458	 => std_logic_vector(to_unsigned(100,8) ,
3459	 => std_logic_vector(to_unsigned(101,8) ,
3460	 => std_logic_vector(to_unsigned(104,8) ,
3461	 => std_logic_vector(to_unsigned(103,8) ,
3462	 => std_logic_vector(to_unsigned(103,8) ,
3463	 => std_logic_vector(to_unsigned(99,8) ,
3464	 => std_logic_vector(to_unsigned(100,8) ,
3465	 => std_logic_vector(to_unsigned(103,8) ,
3466	 => std_logic_vector(to_unsigned(104,8) ,
3467	 => std_logic_vector(to_unsigned(105,8) ,
3468	 => std_logic_vector(to_unsigned(107,8) ,
3469	 => std_logic_vector(to_unsigned(101,8) ,
3470	 => std_logic_vector(to_unsigned(108,8) ,
3471	 => std_logic_vector(to_unsigned(108,8) ,
3472	 => std_logic_vector(to_unsigned(109,8) ,
3473	 => std_logic_vector(to_unsigned(115,8) ,
3474	 => std_logic_vector(to_unsigned(119,8) ,
3475	 => std_logic_vector(to_unsigned(125,8) ,
3476	 => std_logic_vector(to_unsigned(131,8) ,
3477	 => std_logic_vector(to_unsigned(128,8) ,
3478	 => std_logic_vector(to_unsigned(128,8) ,
3479	 => std_logic_vector(to_unsigned(133,8) ,
3480	 => std_logic_vector(to_unsigned(133,8) ,
3481	 => std_logic_vector(to_unsigned(134,8) ,
3482	 => std_logic_vector(to_unsigned(136,8) ,
3483	 => std_logic_vector(to_unsigned(133,8) ,
3484	 => std_logic_vector(to_unsigned(141,8) ,
3485	 => std_logic_vector(to_unsigned(141,8) ,
3486	 => std_logic_vector(to_unsigned(138,8) ,
3487	 => std_logic_vector(to_unsigned(138,8) ,
3488	 => std_logic_vector(to_unsigned(136,8) ,
3489	 => std_logic_vector(to_unsigned(146,8) ,
3490	 => std_logic_vector(to_unsigned(154,8) ,
3491	 => std_logic_vector(to_unsigned(149,8) ,
3492	 => std_logic_vector(to_unsigned(147,8) ,
3493	 => std_logic_vector(to_unsigned(149,8) ,
3494	 => std_logic_vector(to_unsigned(154,8) ,
3495	 => std_logic_vector(to_unsigned(156,8) ,
3496	 => std_logic_vector(to_unsigned(157,8) ,
3497	 => std_logic_vector(to_unsigned(159,8) ,
3498	 => std_logic_vector(to_unsigned(157,8) ,
3499	 => std_logic_vector(to_unsigned(157,8) ,
3500	 => std_logic_vector(to_unsigned(159,8) ,
3501	 => std_logic_vector(to_unsigned(159,8) ,
3502	 => std_logic_vector(to_unsigned(161,8) ,
3503	 => std_logic_vector(to_unsigned(161,8) ,
3504	 => std_logic_vector(to_unsigned(159,8) ,
3505	 => std_logic_vector(to_unsigned(159,8) ,
3506	 => std_logic_vector(to_unsigned(161,8) ,
3507	 => std_logic_vector(to_unsigned(163,8) ,
3508	 => std_logic_vector(to_unsigned(163,8) ,
3509	 => std_logic_vector(to_unsigned(159,8) ,
3510	 => std_logic_vector(to_unsigned(159,8) ,
3511	 => std_logic_vector(to_unsigned(159,8) ,
3512	 => std_logic_vector(to_unsigned(157,8) ,
3513	 => std_logic_vector(to_unsigned(157,8) ,
3514	 => std_logic_vector(to_unsigned(156,8) ,
3515	 => std_logic_vector(to_unsigned(159,8) ,
3516	 => std_logic_vector(to_unsigned(163,8) ,
3517	 => std_logic_vector(to_unsigned(161,8) ,
3518	 => std_logic_vector(to_unsigned(161,8) ,
3519	 => std_logic_vector(to_unsigned(163,8) ,
3520	 => std_logic_vector(to_unsigned(163,8) ,
3521	 => std_logic_vector(to_unsigned(96,8) ,
3522	 => std_logic_vector(to_unsigned(93,8) ,
3523	 => std_logic_vector(to_unsigned(86,8) ,
3524	 => std_logic_vector(to_unsigned(86,8) ,
3525	 => std_logic_vector(to_unsigned(84,8) ,
3526	 => std_logic_vector(to_unsigned(82,8) ,
3527	 => std_logic_vector(to_unsigned(85,8) ,
3528	 => std_logic_vector(to_unsigned(79,8) ,
3529	 => std_logic_vector(to_unsigned(82,8) ,
3530	 => std_logic_vector(to_unsigned(88,8) ,
3531	 => std_logic_vector(to_unsigned(87,8) ,
3532	 => std_logic_vector(to_unsigned(82,8) ,
3533	 => std_logic_vector(to_unsigned(80,8) ,
3534	 => std_logic_vector(to_unsigned(82,8) ,
3535	 => std_logic_vector(to_unsigned(80,8) ,
3536	 => std_logic_vector(to_unsigned(80,8) ,
3537	 => std_logic_vector(to_unsigned(84,8) ,
3538	 => std_logic_vector(to_unsigned(80,8) ,
3539	 => std_logic_vector(to_unsigned(82,8) ,
3540	 => std_logic_vector(to_unsigned(82,8) ,
3541	 => std_logic_vector(to_unsigned(80,8) ,
3542	 => std_logic_vector(to_unsigned(80,8) ,
3543	 => std_logic_vector(to_unsigned(79,8) ,
3544	 => std_logic_vector(to_unsigned(79,8) ,
3545	 => std_logic_vector(to_unsigned(81,8) ,
3546	 => std_logic_vector(to_unsigned(84,8) ,
3547	 => std_logic_vector(to_unsigned(79,8) ,
3548	 => std_logic_vector(to_unsigned(86,8) ,
3549	 => std_logic_vector(to_unsigned(95,8) ,
3550	 => std_logic_vector(to_unsigned(88,8) ,
3551	 => std_logic_vector(to_unsigned(84,8) ,
3552	 => std_logic_vector(to_unsigned(84,8) ,
3553	 => std_logic_vector(to_unsigned(88,8) ,
3554	 => std_logic_vector(to_unsigned(88,8) ,
3555	 => std_logic_vector(to_unsigned(86,8) ,
3556	 => std_logic_vector(to_unsigned(82,8) ,
3557	 => std_logic_vector(to_unsigned(87,8) ,
3558	 => std_logic_vector(to_unsigned(87,8) ,
3559	 => std_logic_vector(to_unsigned(88,8) ,
3560	 => std_logic_vector(to_unsigned(91,8) ,
3561	 => std_logic_vector(to_unsigned(93,8) ,
3562	 => std_logic_vector(to_unsigned(93,8) ,
3563	 => std_logic_vector(to_unsigned(93,8) ,
3564	 => std_logic_vector(to_unsigned(97,8) ,
3565	 => std_logic_vector(to_unsigned(96,8) ,
3566	 => std_logic_vector(to_unsigned(100,8) ,
3567	 => std_logic_vector(to_unsigned(107,8) ,
3568	 => std_logic_vector(to_unsigned(104,8) ,
3569	 => std_logic_vector(to_unsigned(99,8) ,
3570	 => std_logic_vector(to_unsigned(101,8) ,
3571	 => std_logic_vector(to_unsigned(100,8) ,
3572	 => std_logic_vector(to_unsigned(100,8) ,
3573	 => std_logic_vector(to_unsigned(101,8) ,
3574	 => std_logic_vector(to_unsigned(107,8) ,
3575	 => std_logic_vector(to_unsigned(100,8) ,
3576	 => std_logic_vector(to_unsigned(105,8) ,
3577	 => std_logic_vector(to_unsigned(111,8) ,
3578	 => std_logic_vector(to_unsigned(108,8) ,
3579	 => std_logic_vector(to_unsigned(105,8) ,
3580	 => std_logic_vector(to_unsigned(107,8) ,
3581	 => std_logic_vector(to_unsigned(105,8) ,
3582	 => std_logic_vector(to_unsigned(104,8) ,
3583	 => std_logic_vector(to_unsigned(105,8) ,
3584	 => std_logic_vector(to_unsigned(107,8) ,
3585	 => std_logic_vector(to_unsigned(112,8) ,
3586	 => std_logic_vector(to_unsigned(111,8) ,
3587	 => std_logic_vector(to_unsigned(105,8) ,
3588	 => std_logic_vector(to_unsigned(107,8) ,
3589	 => std_logic_vector(to_unsigned(111,8) ,
3590	 => std_logic_vector(to_unsigned(105,8) ,
3591	 => std_logic_vector(to_unsigned(108,8) ,
3592	 => std_logic_vector(to_unsigned(109,8) ,
3593	 => std_logic_vector(to_unsigned(105,8) ,
3594	 => std_logic_vector(to_unsigned(112,8) ,
3595	 => std_logic_vector(to_unsigned(108,8) ,
3596	 => std_logic_vector(to_unsigned(109,8) ,
3597	 => std_logic_vector(to_unsigned(112,8) ,
3598	 => std_logic_vector(to_unsigned(105,8) ,
3599	 => std_logic_vector(to_unsigned(101,8) ,
3600	 => std_logic_vector(to_unsigned(107,8) ,
3601	 => std_logic_vector(to_unsigned(104,8) ,
3602	 => std_logic_vector(to_unsigned(101,8) ,
3603	 => std_logic_vector(to_unsigned(101,8) ,
3604	 => std_logic_vector(to_unsigned(97,8) ,
3605	 => std_logic_vector(to_unsigned(101,8) ,
3606	 => std_logic_vector(to_unsigned(103,8) ,
3607	 => std_logic_vector(to_unsigned(97,8) ,
3608	 => std_logic_vector(to_unsigned(95,8) ,
3609	 => std_logic_vector(to_unsigned(95,8) ,
3610	 => std_logic_vector(to_unsigned(95,8) ,
3611	 => std_logic_vector(to_unsigned(96,8) ,
3612	 => std_logic_vector(to_unsigned(97,8) ,
3613	 => std_logic_vector(to_unsigned(100,8) ,
3614	 => std_logic_vector(to_unsigned(100,8) ,
3615	 => std_logic_vector(to_unsigned(99,8) ,
3616	 => std_logic_vector(to_unsigned(90,8) ,
3617	 => std_logic_vector(to_unsigned(84,8) ,
3618	 => std_logic_vector(to_unsigned(85,8) ,
3619	 => std_logic_vector(to_unsigned(82,8) ,
3620	 => std_logic_vector(to_unsigned(80,8) ,
3621	 => std_logic_vector(to_unsigned(84,8) ,
3622	 => std_logic_vector(to_unsigned(86,8) ,
3623	 => std_logic_vector(to_unsigned(86,8) ,
3624	 => std_logic_vector(to_unsigned(90,8) ,
3625	 => std_logic_vector(to_unsigned(92,8) ,
3626	 => std_logic_vector(to_unsigned(92,8) ,
3627	 => std_logic_vector(to_unsigned(95,8) ,
3628	 => std_logic_vector(to_unsigned(95,8) ,
3629	 => std_logic_vector(to_unsigned(97,8) ,
3630	 => std_logic_vector(to_unsigned(99,8) ,
3631	 => std_logic_vector(to_unsigned(92,8) ,
3632	 => std_logic_vector(to_unsigned(93,8) ,
3633	 => std_logic_vector(to_unsigned(90,8) ,
3634	 => std_logic_vector(to_unsigned(91,8) ,
3635	 => std_logic_vector(to_unsigned(107,8) ,
3636	 => std_logic_vector(to_unsigned(95,8) ,
3637	 => std_logic_vector(to_unsigned(86,8) ,
3638	 => std_logic_vector(to_unsigned(91,8) ,
3639	 => std_logic_vector(to_unsigned(90,8) ,
3640	 => std_logic_vector(to_unsigned(92,8) ,
3641	 => std_logic_vector(to_unsigned(96,8) ,
3642	 => std_logic_vector(to_unsigned(96,8) ,
3643	 => std_logic_vector(to_unsigned(93,8) ,
3644	 => std_logic_vector(to_unsigned(91,8) ,
3645	 => std_logic_vector(to_unsigned(95,8) ,
3646	 => std_logic_vector(to_unsigned(95,8) ,
3647	 => std_logic_vector(to_unsigned(91,8) ,
3648	 => std_logic_vector(to_unsigned(92,8) ,
3649	 => std_logic_vector(to_unsigned(93,8) ,
3650	 => std_logic_vector(to_unsigned(93,8) ,
3651	 => std_logic_vector(to_unsigned(95,8) ,
3652	 => std_logic_vector(to_unsigned(92,8) ,
3653	 => std_logic_vector(to_unsigned(93,8) ,
3654	 => std_logic_vector(to_unsigned(91,8) ,
3655	 => std_logic_vector(to_unsigned(86,8) ,
3656	 => std_logic_vector(to_unsigned(91,8) ,
3657	 => std_logic_vector(to_unsigned(97,8) ,
3658	 => std_logic_vector(to_unsigned(97,8) ,
3659	 => std_logic_vector(to_unsigned(91,8) ,
3660	 => std_logic_vector(to_unsigned(93,8) ,
3661	 => std_logic_vector(to_unsigned(101,8) ,
3662	 => std_logic_vector(to_unsigned(101,8) ,
3663	 => std_logic_vector(to_unsigned(97,8) ,
3664	 => std_logic_vector(to_unsigned(95,8) ,
3665	 => std_logic_vector(to_unsigned(99,8) ,
3666	 => std_logic_vector(to_unsigned(100,8) ,
3667	 => std_logic_vector(to_unsigned(93,8) ,
3668	 => std_logic_vector(to_unsigned(92,8) ,
3669	 => std_logic_vector(to_unsigned(96,8) ,
3670	 => std_logic_vector(to_unsigned(91,8) ,
3671	 => std_logic_vector(to_unsigned(90,8) ,
3672	 => std_logic_vector(to_unsigned(88,8) ,
3673	 => std_logic_vector(to_unsigned(85,8) ,
3674	 => std_logic_vector(to_unsigned(80,8) ,
3675	 => std_logic_vector(to_unsigned(79,8) ,
3676	 => std_logic_vector(to_unsigned(85,8) ,
3677	 => std_logic_vector(to_unsigned(82,8) ,
3678	 => std_logic_vector(to_unsigned(82,8) ,
3679	 => std_logic_vector(to_unsigned(79,8) ,
3680	 => std_logic_vector(to_unsigned(85,8) ,
3681	 => std_logic_vector(to_unsigned(88,8) ,
3682	 => std_logic_vector(to_unsigned(82,8) ,
3683	 => std_logic_vector(to_unsigned(81,8) ,
3684	 => std_logic_vector(to_unsigned(80,8) ,
3685	 => std_logic_vector(to_unsigned(82,8) ,
3686	 => std_logic_vector(to_unsigned(87,8) ,
3687	 => std_logic_vector(to_unsigned(85,8) ,
3688	 => std_logic_vector(to_unsigned(86,8) ,
3689	 => std_logic_vector(to_unsigned(87,8) ,
3690	 => std_logic_vector(to_unsigned(85,8) ,
3691	 => std_logic_vector(to_unsigned(80,8) ,
3692	 => std_logic_vector(to_unsigned(85,8) ,
3693	 => std_logic_vector(to_unsigned(86,8) ,
3694	 => std_logic_vector(to_unsigned(87,8) ,
3695	 => std_logic_vector(to_unsigned(85,8) ,
3696	 => std_logic_vector(to_unsigned(78,8) ,
3697	 => std_logic_vector(to_unsigned(79,8) ,
3698	 => std_logic_vector(to_unsigned(80,8) ,
3699	 => std_logic_vector(to_unsigned(72,8) ,
3700	 => std_logic_vector(to_unsigned(78,8) ,
3701	 => std_logic_vector(to_unsigned(80,8) ,
3702	 => std_logic_vector(to_unsigned(72,8) ,
3703	 => std_logic_vector(to_unsigned(66,8) ,
3704	 => std_logic_vector(to_unsigned(69,8) ,
3705	 => std_logic_vector(to_unsigned(70,8) ,
3706	 => std_logic_vector(to_unsigned(71,8) ,
3707	 => std_logic_vector(to_unsigned(73,8) ,
3708	 => std_logic_vector(to_unsigned(67,8) ,
3709	 => std_logic_vector(to_unsigned(68,8) ,
3710	 => std_logic_vector(to_unsigned(73,8) ,
3711	 => std_logic_vector(to_unsigned(69,8) ,
3712	 => std_logic_vector(to_unsigned(67,8) ,
3713	 => std_logic_vector(to_unsigned(74,8) ,
3714	 => std_logic_vector(to_unsigned(77,8) ,
3715	 => std_logic_vector(to_unsigned(72,8) ,
3716	 => std_logic_vector(to_unsigned(71,8) ,
3717	 => std_logic_vector(to_unsigned(70,8) ,
3718	 => std_logic_vector(to_unsigned(73,8) ,
3719	 => std_logic_vector(to_unsigned(72,8) ,
3720	 => std_logic_vector(to_unsigned(73,8) ,
3721	 => std_logic_vector(to_unsigned(74,8) ,
3722	 => std_logic_vector(to_unsigned(76,8) ,
3723	 => std_logic_vector(to_unsigned(81,8) ,
3724	 => std_logic_vector(to_unsigned(74,8) ,
3725	 => std_logic_vector(to_unsigned(76,8) ,
3726	 => std_logic_vector(to_unsigned(78,8) ,
3727	 => std_logic_vector(to_unsigned(81,8) ,
3728	 => std_logic_vector(to_unsigned(78,8) ,
3729	 => std_logic_vector(to_unsigned(79,8) ,
3730	 => std_logic_vector(to_unsigned(84,8) ,
3731	 => std_logic_vector(to_unsigned(82,8) ,
3732	 => std_logic_vector(to_unsigned(79,8) ,
3733	 => std_logic_vector(to_unsigned(78,8) ,
3734	 => std_logic_vector(to_unsigned(81,8) ,
3735	 => std_logic_vector(to_unsigned(78,8) ,
3736	 => std_logic_vector(to_unsigned(77,8) ,
3737	 => std_logic_vector(to_unsigned(79,8) ,
3738	 => std_logic_vector(to_unsigned(80,8) ,
3739	 => std_logic_vector(to_unsigned(81,8) ,
3740	 => std_logic_vector(to_unsigned(84,8) ,
3741	 => std_logic_vector(to_unsigned(88,8) ,
3742	 => std_logic_vector(to_unsigned(86,8) ,
3743	 => std_logic_vector(to_unsigned(82,8) ,
3744	 => std_logic_vector(to_unsigned(87,8) ,
3745	 => std_logic_vector(to_unsigned(90,8) ,
3746	 => std_logic_vector(to_unsigned(91,8) ,
3747	 => std_logic_vector(to_unsigned(93,8) ,
3748	 => std_logic_vector(to_unsigned(86,8) ,
3749	 => std_logic_vector(to_unsigned(86,8) ,
3750	 => std_logic_vector(to_unsigned(80,8) ,
3751	 => std_logic_vector(to_unsigned(72,8) ,
3752	 => std_logic_vector(to_unsigned(86,8) ,
3753	 => std_logic_vector(to_unsigned(90,8) ,
3754	 => std_logic_vector(to_unsigned(81,8) ,
3755	 => std_logic_vector(to_unsigned(80,8) ,
3756	 => std_logic_vector(to_unsigned(86,8) ,
3757	 => std_logic_vector(to_unsigned(70,8) ,
3758	 => std_logic_vector(to_unsigned(3,8) ,
3759	 => std_logic_vector(to_unsigned(0,8) ,
3760	 => std_logic_vector(to_unsigned(0,8) ,
3761	 => std_logic_vector(to_unsigned(23,8) ,
3762	 => std_logic_vector(to_unsigned(103,8) ,
3763	 => std_logic_vector(to_unsigned(90,8) ,
3764	 => std_logic_vector(to_unsigned(91,8) ,
3765	 => std_logic_vector(to_unsigned(92,8) ,
3766	 => std_logic_vector(to_unsigned(97,8) ,
3767	 => std_logic_vector(to_unsigned(97,8) ,
3768	 => std_logic_vector(to_unsigned(92,8) ,
3769	 => std_logic_vector(to_unsigned(99,8) ,
3770	 => std_logic_vector(to_unsigned(104,8) ,
3771	 => std_logic_vector(to_unsigned(115,8) ,
3772	 => std_logic_vector(to_unsigned(118,8) ,
3773	 => std_logic_vector(to_unsigned(104,8) ,
3774	 => std_logic_vector(to_unsigned(107,8) ,
3775	 => std_logic_vector(to_unsigned(114,8) ,
3776	 => std_logic_vector(to_unsigned(109,8) ,
3777	 => std_logic_vector(to_unsigned(103,8) ,
3778	 => std_logic_vector(to_unsigned(101,8) ,
3779	 => std_logic_vector(to_unsigned(97,8) ,
3780	 => std_logic_vector(to_unsigned(95,8) ,
3781	 => std_logic_vector(to_unsigned(99,8) ,
3782	 => std_logic_vector(to_unsigned(104,8) ,
3783	 => std_logic_vector(to_unsigned(101,8) ,
3784	 => std_logic_vector(to_unsigned(105,8) ,
3785	 => std_logic_vector(to_unsigned(105,8) ,
3786	 => std_logic_vector(to_unsigned(101,8) ,
3787	 => std_logic_vector(to_unsigned(101,8) ,
3788	 => std_logic_vector(to_unsigned(96,8) ,
3789	 => std_logic_vector(to_unsigned(95,8) ,
3790	 => std_logic_vector(to_unsigned(105,8) ,
3791	 => std_logic_vector(to_unsigned(107,8) ,
3792	 => std_logic_vector(to_unsigned(108,8) ,
3793	 => std_logic_vector(to_unsigned(114,8) ,
3794	 => std_logic_vector(to_unsigned(115,8) ,
3795	 => std_logic_vector(to_unsigned(116,8) ,
3796	 => std_logic_vector(to_unsigned(124,8) ,
3797	 => std_logic_vector(to_unsigned(130,8) ,
3798	 => std_logic_vector(to_unsigned(121,8) ,
3799	 => std_logic_vector(to_unsigned(122,8) ,
3800	 => std_logic_vector(to_unsigned(128,8) ,
3801	 => std_logic_vector(to_unsigned(128,8) ,
3802	 => std_logic_vector(to_unsigned(130,8) ,
3803	 => std_logic_vector(to_unsigned(125,8) ,
3804	 => std_logic_vector(to_unsigned(131,8) ,
3805	 => std_logic_vector(to_unsigned(136,8) ,
3806	 => std_logic_vector(to_unsigned(136,8) ,
3807	 => std_logic_vector(to_unsigned(133,8) ,
3808	 => std_logic_vector(to_unsigned(127,8) ,
3809	 => std_logic_vector(to_unsigned(128,8) ,
3810	 => std_logic_vector(to_unsigned(139,8) ,
3811	 => std_logic_vector(to_unsigned(146,8) ,
3812	 => std_logic_vector(to_unsigned(147,8) ,
3813	 => std_logic_vector(to_unsigned(147,8) ,
3814	 => std_logic_vector(to_unsigned(151,8) ,
3815	 => std_logic_vector(to_unsigned(154,8) ,
3816	 => std_logic_vector(to_unsigned(152,8) ,
3817	 => std_logic_vector(to_unsigned(154,8) ,
3818	 => std_logic_vector(to_unsigned(152,8) ,
3819	 => std_logic_vector(to_unsigned(159,8) ,
3820	 => std_logic_vector(to_unsigned(159,8) ,
3821	 => std_logic_vector(to_unsigned(157,8) ,
3822	 => std_logic_vector(to_unsigned(159,8) ,
3823	 => std_logic_vector(to_unsigned(159,8) ,
3824	 => std_logic_vector(to_unsigned(159,8) ,
3825	 => std_logic_vector(to_unsigned(159,8) ,
3826	 => std_logic_vector(to_unsigned(159,8) ,
3827	 => std_logic_vector(to_unsigned(159,8) ,
3828	 => std_logic_vector(to_unsigned(159,8) ,
3829	 => std_logic_vector(to_unsigned(159,8) ,
3830	 => std_logic_vector(to_unsigned(163,8) ,
3831	 => std_logic_vector(to_unsigned(159,8) ,
3832	 => std_logic_vector(to_unsigned(157,8) ,
3833	 => std_logic_vector(to_unsigned(157,8) ,
3834	 => std_logic_vector(to_unsigned(154,8) ,
3835	 => std_logic_vector(to_unsigned(161,8) ,
3836	 => std_logic_vector(to_unsigned(161,8) ,
3837	 => std_logic_vector(to_unsigned(156,8) ,
3838	 => std_logic_vector(to_unsigned(157,8) ,
3839	 => std_logic_vector(to_unsigned(159,8) ,
3840	 => std_logic_vector(to_unsigned(157,8) ,
3841	 => std_logic_vector(to_unsigned(93,8) ,
3842	 => std_logic_vector(to_unsigned(90,8) ,
3843	 => std_logic_vector(to_unsigned(87,8) ,
3844	 => std_logic_vector(to_unsigned(84,8) ,
3845	 => std_logic_vector(to_unsigned(81,8) ,
3846	 => std_logic_vector(to_unsigned(86,8) ,
3847	 => std_logic_vector(to_unsigned(88,8) ,
3848	 => std_logic_vector(to_unsigned(85,8) ,
3849	 => std_logic_vector(to_unsigned(81,8) ,
3850	 => std_logic_vector(to_unsigned(80,8) ,
3851	 => std_logic_vector(to_unsigned(86,8) ,
3852	 => std_logic_vector(to_unsigned(82,8) ,
3853	 => std_logic_vector(to_unsigned(81,8) ,
3854	 => std_logic_vector(to_unsigned(78,8) ,
3855	 => std_logic_vector(to_unsigned(74,8) ,
3856	 => std_logic_vector(to_unsigned(81,8) ,
3857	 => std_logic_vector(to_unsigned(84,8) ,
3858	 => std_logic_vector(to_unsigned(78,8) ,
3859	 => std_logic_vector(to_unsigned(73,8) ,
3860	 => std_logic_vector(to_unsigned(81,8) ,
3861	 => std_logic_vector(to_unsigned(82,8) ,
3862	 => std_logic_vector(to_unsigned(80,8) ,
3863	 => std_logic_vector(to_unsigned(80,8) ,
3864	 => std_logic_vector(to_unsigned(77,8) ,
3865	 => std_logic_vector(to_unsigned(77,8) ,
3866	 => std_logic_vector(to_unsigned(82,8) ,
3867	 => std_logic_vector(to_unsigned(80,8) ,
3868	 => std_logic_vector(to_unsigned(82,8) ,
3869	 => std_logic_vector(to_unsigned(85,8) ,
3870	 => std_logic_vector(to_unsigned(78,8) ,
3871	 => std_logic_vector(to_unsigned(81,8) ,
3872	 => std_logic_vector(to_unsigned(85,8) ,
3873	 => std_logic_vector(to_unsigned(90,8) ,
3874	 => std_logic_vector(to_unsigned(87,8) ,
3875	 => std_logic_vector(to_unsigned(86,8) ,
3876	 => std_logic_vector(to_unsigned(87,8) ,
3877	 => std_logic_vector(to_unsigned(87,8) ,
3878	 => std_logic_vector(to_unsigned(87,8) ,
3879	 => std_logic_vector(to_unsigned(85,8) ,
3880	 => std_logic_vector(to_unsigned(91,8) ,
3881	 => std_logic_vector(to_unsigned(91,8) ,
3882	 => std_logic_vector(to_unsigned(87,8) ,
3883	 => std_logic_vector(to_unsigned(92,8) ,
3884	 => std_logic_vector(to_unsigned(93,8) ,
3885	 => std_logic_vector(to_unsigned(92,8) ,
3886	 => std_logic_vector(to_unsigned(96,8) ,
3887	 => std_logic_vector(to_unsigned(100,8) ,
3888	 => std_logic_vector(to_unsigned(99,8) ,
3889	 => std_logic_vector(to_unsigned(99,8) ,
3890	 => std_logic_vector(to_unsigned(100,8) ,
3891	 => std_logic_vector(to_unsigned(93,8) ,
3892	 => std_logic_vector(to_unsigned(101,8) ,
3893	 => std_logic_vector(to_unsigned(104,8) ,
3894	 => std_logic_vector(to_unsigned(107,8) ,
3895	 => std_logic_vector(to_unsigned(104,8) ,
3896	 => std_logic_vector(to_unsigned(104,8) ,
3897	 => std_logic_vector(to_unsigned(107,8) ,
3898	 => std_logic_vector(to_unsigned(109,8) ,
3899	 => std_logic_vector(to_unsigned(104,8) ,
3900	 => std_logic_vector(to_unsigned(108,8) ,
3901	 => std_logic_vector(to_unsigned(115,8) ,
3902	 => std_logic_vector(to_unsigned(107,8) ,
3903	 => std_logic_vector(to_unsigned(104,8) ,
3904	 => std_logic_vector(to_unsigned(108,8) ,
3905	 => std_logic_vector(to_unsigned(112,8) ,
3906	 => std_logic_vector(to_unsigned(116,8) ,
3907	 => std_logic_vector(to_unsigned(112,8) ,
3908	 => std_logic_vector(to_unsigned(114,8) ,
3909	 => std_logic_vector(to_unsigned(112,8) ,
3910	 => std_logic_vector(to_unsigned(108,8) ,
3911	 => std_logic_vector(to_unsigned(109,8) ,
3912	 => std_logic_vector(to_unsigned(109,8) ,
3913	 => std_logic_vector(to_unsigned(107,8) ,
3914	 => std_logic_vector(to_unsigned(108,8) ,
3915	 => std_logic_vector(to_unsigned(109,8) ,
3916	 => std_logic_vector(to_unsigned(111,8) ,
3917	 => std_logic_vector(to_unsigned(107,8) ,
3918	 => std_logic_vector(to_unsigned(103,8) ,
3919	 => std_logic_vector(to_unsigned(100,8) ,
3920	 => std_logic_vector(to_unsigned(99,8) ,
3921	 => std_logic_vector(to_unsigned(96,8) ,
3922	 => std_logic_vector(to_unsigned(96,8) ,
3923	 => std_logic_vector(to_unsigned(101,8) ,
3924	 => std_logic_vector(to_unsigned(99,8) ,
3925	 => std_logic_vector(to_unsigned(99,8) ,
3926	 => std_logic_vector(to_unsigned(100,8) ,
3927	 => std_logic_vector(to_unsigned(96,8) ,
3928	 => std_logic_vector(to_unsigned(97,8) ,
3929	 => std_logic_vector(to_unsigned(93,8) ,
3930	 => std_logic_vector(to_unsigned(91,8) ,
3931	 => std_logic_vector(to_unsigned(95,8) ,
3932	 => std_logic_vector(to_unsigned(93,8) ,
3933	 => std_logic_vector(to_unsigned(93,8) ,
3934	 => std_logic_vector(to_unsigned(95,8) ,
3935	 => std_logic_vector(to_unsigned(91,8) ,
3936	 => std_logic_vector(to_unsigned(84,8) ,
3937	 => std_logic_vector(to_unsigned(77,8) ,
3938	 => std_logic_vector(to_unsigned(77,8) ,
3939	 => std_logic_vector(to_unsigned(82,8) ,
3940	 => std_logic_vector(to_unsigned(85,8) ,
3941	 => std_logic_vector(to_unsigned(82,8) ,
3942	 => std_logic_vector(to_unsigned(85,8) ,
3943	 => std_logic_vector(to_unsigned(85,8) ,
3944	 => std_logic_vector(to_unsigned(87,8) ,
3945	 => std_logic_vector(to_unsigned(88,8) ,
3946	 => std_logic_vector(to_unsigned(87,8) ,
3947	 => std_logic_vector(to_unsigned(92,8) ,
3948	 => std_logic_vector(to_unsigned(88,8) ,
3949	 => std_logic_vector(to_unsigned(87,8) ,
3950	 => std_logic_vector(to_unsigned(91,8) ,
3951	 => std_logic_vector(to_unsigned(88,8) ,
3952	 => std_logic_vector(to_unsigned(90,8) ,
3953	 => std_logic_vector(to_unsigned(90,8) ,
3954	 => std_logic_vector(to_unsigned(93,8) ,
3955	 => std_logic_vector(to_unsigned(107,8) ,
3956	 => std_logic_vector(to_unsigned(93,8) ,
3957	 => std_logic_vector(to_unsigned(80,8) ,
3958	 => std_logic_vector(to_unsigned(90,8) ,
3959	 => std_logic_vector(to_unsigned(91,8) ,
3960	 => std_logic_vector(to_unsigned(91,8) ,
3961	 => std_logic_vector(to_unsigned(93,8) ,
3962	 => std_logic_vector(to_unsigned(93,8) ,
3963	 => std_logic_vector(to_unsigned(92,8) ,
3964	 => std_logic_vector(to_unsigned(91,8) ,
3965	 => std_logic_vector(to_unsigned(91,8) ,
3966	 => std_logic_vector(to_unsigned(87,8) ,
3967	 => std_logic_vector(to_unsigned(86,8) ,
3968	 => std_logic_vector(to_unsigned(90,8) ,
3969	 => std_logic_vector(to_unsigned(91,8) ,
3970	 => std_logic_vector(to_unsigned(91,8) ,
3971	 => std_logic_vector(to_unsigned(93,8) ,
3972	 => std_logic_vector(to_unsigned(96,8) ,
3973	 => std_logic_vector(to_unsigned(91,8) ,
3974	 => std_logic_vector(to_unsigned(87,8) ,
3975	 => std_logic_vector(to_unsigned(88,8) ,
3976	 => std_logic_vector(to_unsigned(96,8) ,
3977	 => std_logic_vector(to_unsigned(95,8) ,
3978	 => std_logic_vector(to_unsigned(93,8) ,
3979	 => std_logic_vector(to_unsigned(91,8) ,
3980	 => std_logic_vector(to_unsigned(96,8) ,
3981	 => std_logic_vector(to_unsigned(99,8) ,
3982	 => std_logic_vector(to_unsigned(99,8) ,
3983	 => std_logic_vector(to_unsigned(99,8) ,
3984	 => std_logic_vector(to_unsigned(95,8) ,
3985	 => std_logic_vector(to_unsigned(97,8) ,
3986	 => std_logic_vector(to_unsigned(96,8) ,
3987	 => std_logic_vector(to_unsigned(93,8) ,
3988	 => std_logic_vector(to_unsigned(92,8) ,
3989	 => std_logic_vector(to_unsigned(91,8) ,
3990	 => std_logic_vector(to_unsigned(88,8) ,
3991	 => std_logic_vector(to_unsigned(90,8) ,
3992	 => std_logic_vector(to_unsigned(88,8) ,
3993	 => std_logic_vector(to_unsigned(88,8) ,
3994	 => std_logic_vector(to_unsigned(87,8) ,
3995	 => std_logic_vector(to_unsigned(85,8) ,
3996	 => std_logic_vector(to_unsigned(85,8) ,
3997	 => std_logic_vector(to_unsigned(81,8) ,
3998	 => std_logic_vector(to_unsigned(82,8) ,
3999	 => std_logic_vector(to_unsigned(82,8) ,
4000	 => std_logic_vector(to_unsigned(88,8) ,
4001	 => std_logic_vector(to_unsigned(88,8) ,
4002	 => std_logic_vector(to_unsigned(82,8) ,
4003	 => std_logic_vector(to_unsigned(82,8) ,
4004	 => std_logic_vector(to_unsigned(85,8) ,
4005	 => std_logic_vector(to_unsigned(87,8) ,
4006	 => std_logic_vector(to_unsigned(85,8) ,
4007	 => std_logic_vector(to_unsigned(84,8) ,
4008	 => std_logic_vector(to_unsigned(84,8) ,
4009	 => std_logic_vector(to_unsigned(85,8) ,
4010	 => std_logic_vector(to_unsigned(84,8) ,
4011	 => std_logic_vector(to_unsigned(79,8) ,
4012	 => std_logic_vector(to_unsigned(77,8) ,
4013	 => std_logic_vector(to_unsigned(79,8) ,
4014	 => std_logic_vector(to_unsigned(80,8) ,
4015	 => std_logic_vector(to_unsigned(81,8) ,
4016	 => std_logic_vector(to_unsigned(81,8) ,
4017	 => std_logic_vector(to_unsigned(79,8) ,
4018	 => std_logic_vector(to_unsigned(78,8) ,
4019	 => std_logic_vector(to_unsigned(73,8) ,
4020	 => std_logic_vector(to_unsigned(76,8) ,
4021	 => std_logic_vector(to_unsigned(77,8) ,
4022	 => std_logic_vector(to_unsigned(78,8) ,
4023	 => std_logic_vector(to_unsigned(71,8) ,
4024	 => std_logic_vector(to_unsigned(66,8) ,
4025	 => std_logic_vector(to_unsigned(63,8) ,
4026	 => std_logic_vector(to_unsigned(62,8) ,
4027	 => std_logic_vector(to_unsigned(71,8) ,
4028	 => std_logic_vector(to_unsigned(73,8) ,
4029	 => std_logic_vector(to_unsigned(64,8) ,
4030	 => std_logic_vector(to_unsigned(70,8) ,
4031	 => std_logic_vector(to_unsigned(73,8) ,
4032	 => std_logic_vector(to_unsigned(74,8) ,
4033	 => std_logic_vector(to_unsigned(77,8) ,
4034	 => std_logic_vector(to_unsigned(74,8) ,
4035	 => std_logic_vector(to_unsigned(73,8) ,
4036	 => std_logic_vector(to_unsigned(74,8) ,
4037	 => std_logic_vector(to_unsigned(71,8) ,
4038	 => std_logic_vector(to_unsigned(70,8) ,
4039	 => std_logic_vector(to_unsigned(73,8) ,
4040	 => std_logic_vector(to_unsigned(77,8) ,
4041	 => std_logic_vector(to_unsigned(77,8) ,
4042	 => std_logic_vector(to_unsigned(73,8) ,
4043	 => std_logic_vector(to_unsigned(71,8) ,
4044	 => std_logic_vector(to_unsigned(70,8) ,
4045	 => std_logic_vector(to_unsigned(74,8) ,
4046	 => std_logic_vector(to_unsigned(73,8) ,
4047	 => std_logic_vector(to_unsigned(77,8) ,
4048	 => std_logic_vector(to_unsigned(80,8) ,
4049	 => std_logic_vector(to_unsigned(78,8) ,
4050	 => std_logic_vector(to_unsigned(82,8) ,
4051	 => std_logic_vector(to_unsigned(82,8) ,
4052	 => std_logic_vector(to_unsigned(78,8) ,
4053	 => std_logic_vector(to_unsigned(77,8) ,
4054	 => std_logic_vector(to_unsigned(79,8) ,
4055	 => std_logic_vector(to_unsigned(82,8) ,
4056	 => std_logic_vector(to_unsigned(81,8) ,
4057	 => std_logic_vector(to_unsigned(77,8) ,
4058	 => std_logic_vector(to_unsigned(76,8) ,
4059	 => std_logic_vector(to_unsigned(78,8) ,
4060	 => std_logic_vector(to_unsigned(79,8) ,
4061	 => std_logic_vector(to_unsigned(85,8) ,
4062	 => std_logic_vector(to_unsigned(81,8) ,
4063	 => std_logic_vector(to_unsigned(80,8) ,
4064	 => std_logic_vector(to_unsigned(81,8) ,
4065	 => std_logic_vector(to_unsigned(82,8) ,
4066	 => std_logic_vector(to_unsigned(85,8) ,
4067	 => std_logic_vector(to_unsigned(85,8) ,
4068	 => std_logic_vector(to_unsigned(85,8) ,
4069	 => std_logic_vector(to_unsigned(88,8) ,
4070	 => std_logic_vector(to_unsigned(80,8) ,
4071	 => std_logic_vector(to_unsigned(69,8) ,
4072	 => std_logic_vector(to_unsigned(82,8) ,
4073	 => std_logic_vector(to_unsigned(88,8) ,
4074	 => std_logic_vector(to_unsigned(81,8) ,
4075	 => std_logic_vector(to_unsigned(80,8) ,
4076	 => std_logic_vector(to_unsigned(87,8) ,
4077	 => std_logic_vector(to_unsigned(82,8) ,
4078	 => std_logic_vector(to_unsigned(12,8) ,
4079	 => std_logic_vector(to_unsigned(0,8) ,
4080	 => std_logic_vector(to_unsigned(0,8) ,
4081	 => std_logic_vector(to_unsigned(9,8) ,
4082	 => std_logic_vector(to_unsigned(86,8) ,
4083	 => std_logic_vector(to_unsigned(93,8) ,
4084	 => std_logic_vector(to_unsigned(88,8) ,
4085	 => std_logic_vector(to_unsigned(90,8) ,
4086	 => std_logic_vector(to_unsigned(92,8) ,
4087	 => std_logic_vector(to_unsigned(91,8) ,
4088	 => std_logic_vector(to_unsigned(99,8) ,
4089	 => std_logic_vector(to_unsigned(105,8) ,
4090	 => std_logic_vector(to_unsigned(105,8) ,
4091	 => std_logic_vector(to_unsigned(114,8) ,
4092	 => std_logic_vector(to_unsigned(118,8) ,
4093	 => std_logic_vector(to_unsigned(108,8) ,
4094	 => std_logic_vector(to_unsigned(104,8) ,
4095	 => std_logic_vector(to_unsigned(112,8) ,
4096	 => std_logic_vector(to_unsigned(114,8) ,
4097	 => std_logic_vector(to_unsigned(104,8) ,
4098	 => std_logic_vector(to_unsigned(96,8) ,
4099	 => std_logic_vector(to_unsigned(92,8) ,
4100	 => std_logic_vector(to_unsigned(93,8) ,
4101	 => std_logic_vector(to_unsigned(96,8) ,
4102	 => std_logic_vector(to_unsigned(103,8) ,
4103	 => std_logic_vector(to_unsigned(97,8) ,
4104	 => std_logic_vector(to_unsigned(100,8) ,
4105	 => std_logic_vector(to_unsigned(107,8) ,
4106	 => std_logic_vector(to_unsigned(100,8) ,
4107	 => std_logic_vector(to_unsigned(96,8) ,
4108	 => std_logic_vector(to_unsigned(99,8) ,
4109	 => std_logic_vector(to_unsigned(99,8) ,
4110	 => std_logic_vector(to_unsigned(101,8) ,
4111	 => std_logic_vector(to_unsigned(103,8) ,
4112	 => std_logic_vector(to_unsigned(108,8) ,
4113	 => std_logic_vector(to_unsigned(107,8) ,
4114	 => std_logic_vector(to_unsigned(108,8) ,
4115	 => std_logic_vector(to_unsigned(112,8) ,
4116	 => std_logic_vector(to_unsigned(116,8) ,
4117	 => std_logic_vector(to_unsigned(122,8) ,
4118	 => std_logic_vector(to_unsigned(118,8) ,
4119	 => std_logic_vector(to_unsigned(116,8) ,
4120	 => std_logic_vector(to_unsigned(122,8) ,
4121	 => std_logic_vector(to_unsigned(122,8) ,
4122	 => std_logic_vector(to_unsigned(124,8) ,
4123	 => std_logic_vector(to_unsigned(125,8) ,
4124	 => std_logic_vector(to_unsigned(125,8) ,
4125	 => std_logic_vector(to_unsigned(128,8) ,
4126	 => std_logic_vector(to_unsigned(141,8) ,
4127	 => std_logic_vector(to_unsigned(136,8) ,
4128	 => std_logic_vector(to_unsigned(121,8) ,
4129	 => std_logic_vector(to_unsigned(121,8) ,
4130	 => std_logic_vector(to_unsigned(130,8) ,
4131	 => std_logic_vector(to_unsigned(134,8) ,
4132	 => std_logic_vector(to_unsigned(136,8) ,
4133	 => std_logic_vector(to_unsigned(144,8) ,
4134	 => std_logic_vector(to_unsigned(146,8) ,
4135	 => std_logic_vector(to_unsigned(147,8) ,
4136	 => std_logic_vector(to_unsigned(147,8) ,
4137	 => std_logic_vector(to_unsigned(151,8) ,
4138	 => std_logic_vector(to_unsigned(154,8) ,
4139	 => std_logic_vector(to_unsigned(156,8) ,
4140	 => std_logic_vector(to_unsigned(157,8) ,
4141	 => std_logic_vector(to_unsigned(154,8) ,
4142	 => std_logic_vector(to_unsigned(156,8) ,
4143	 => std_logic_vector(to_unsigned(161,8) ,
4144	 => std_logic_vector(to_unsigned(161,8) ,
4145	 => std_logic_vector(to_unsigned(161,8) ,
4146	 => std_logic_vector(to_unsigned(159,8) ,
4147	 => std_logic_vector(to_unsigned(157,8) ,
4148	 => std_logic_vector(to_unsigned(157,8) ,
4149	 => std_logic_vector(to_unsigned(159,8) ,
4150	 => std_logic_vector(to_unsigned(163,8) ,
4151	 => std_logic_vector(to_unsigned(163,8) ,
4152	 => std_logic_vector(to_unsigned(156,8) ,
4153	 => std_logic_vector(to_unsigned(157,8) ,
4154	 => std_logic_vector(to_unsigned(161,8) ,
4155	 => std_logic_vector(to_unsigned(157,8) ,
4156	 => std_logic_vector(to_unsigned(157,8) ,
4157	 => std_logic_vector(to_unsigned(161,8) ,
4158	 => std_logic_vector(to_unsigned(161,8) ,
4159	 => std_logic_vector(to_unsigned(163,8) ,
4160	 => std_logic_vector(to_unsigned(161,8) ,
4161	 => std_logic_vector(to_unsigned(92,8) ,
4162	 => std_logic_vector(to_unsigned(90,8) ,
4163	 => std_logic_vector(to_unsigned(86,8) ,
4164	 => std_logic_vector(to_unsigned(79,8) ,
4165	 => std_logic_vector(to_unsigned(82,8) ,
4166	 => std_logic_vector(to_unsigned(90,8) ,
4167	 => std_logic_vector(to_unsigned(90,8) ,
4168	 => std_logic_vector(to_unsigned(86,8) ,
4169	 => std_logic_vector(to_unsigned(79,8) ,
4170	 => std_logic_vector(to_unsigned(73,8) ,
4171	 => std_logic_vector(to_unsigned(81,8) ,
4172	 => std_logic_vector(to_unsigned(82,8) ,
4173	 => std_logic_vector(to_unsigned(85,8) ,
4174	 => std_logic_vector(to_unsigned(79,8) ,
4175	 => std_logic_vector(to_unsigned(77,8) ,
4176	 => std_logic_vector(to_unsigned(79,8) ,
4177	 => std_logic_vector(to_unsigned(79,8) ,
4178	 => std_logic_vector(to_unsigned(81,8) ,
4179	 => std_logic_vector(to_unsigned(79,8) ,
4180	 => std_logic_vector(to_unsigned(80,8) ,
4181	 => std_logic_vector(to_unsigned(82,8) ,
4182	 => std_logic_vector(to_unsigned(85,8) ,
4183	 => std_logic_vector(to_unsigned(84,8) ,
4184	 => std_logic_vector(to_unsigned(81,8) ,
4185	 => std_logic_vector(to_unsigned(73,8) ,
4186	 => std_logic_vector(to_unsigned(80,8) ,
4187	 => std_logic_vector(to_unsigned(81,8) ,
4188	 => std_logic_vector(to_unsigned(81,8) ,
4189	 => std_logic_vector(to_unsigned(82,8) ,
4190	 => std_logic_vector(to_unsigned(72,8) ,
4191	 => std_logic_vector(to_unsigned(76,8) ,
4192	 => std_logic_vector(to_unsigned(84,8) ,
4193	 => std_logic_vector(to_unsigned(81,8) ,
4194	 => std_logic_vector(to_unsigned(80,8) ,
4195	 => std_logic_vector(to_unsigned(82,8) ,
4196	 => std_logic_vector(to_unsigned(84,8) ,
4197	 => std_logic_vector(to_unsigned(81,8) ,
4198	 => std_logic_vector(to_unsigned(88,8) ,
4199	 => std_logic_vector(to_unsigned(88,8) ,
4200	 => std_logic_vector(to_unsigned(88,8) ,
4201	 => std_logic_vector(to_unsigned(93,8) ,
4202	 => std_logic_vector(to_unsigned(91,8) ,
4203	 => std_logic_vector(to_unsigned(90,8) ,
4204	 => std_logic_vector(to_unsigned(88,8) ,
4205	 => std_logic_vector(to_unsigned(91,8) ,
4206	 => std_logic_vector(to_unsigned(96,8) ,
4207	 => std_logic_vector(to_unsigned(96,8) ,
4208	 => std_logic_vector(to_unsigned(96,8) ,
4209	 => std_logic_vector(to_unsigned(97,8) ,
4210	 => std_logic_vector(to_unsigned(104,8) ,
4211	 => std_logic_vector(to_unsigned(100,8) ,
4212	 => std_logic_vector(to_unsigned(97,8) ,
4213	 => std_logic_vector(to_unsigned(104,8) ,
4214	 => std_logic_vector(to_unsigned(105,8) ,
4215	 => std_logic_vector(to_unsigned(107,8) ,
4216	 => std_logic_vector(to_unsigned(107,8) ,
4217	 => std_logic_vector(to_unsigned(105,8) ,
4218	 => std_logic_vector(to_unsigned(112,8) ,
4219	 => std_logic_vector(to_unsigned(112,8) ,
4220	 => std_logic_vector(to_unsigned(118,8) ,
4221	 => std_logic_vector(to_unsigned(116,8) ,
4222	 => std_logic_vector(to_unsigned(108,8) ,
4223	 => std_logic_vector(to_unsigned(105,8) ,
4224	 => std_logic_vector(to_unsigned(107,8) ,
4225	 => std_logic_vector(to_unsigned(108,8) ,
4226	 => std_logic_vector(to_unsigned(112,8) ,
4227	 => std_logic_vector(to_unsigned(111,8) ,
4228	 => std_logic_vector(to_unsigned(109,8) ,
4229	 => std_logic_vector(to_unsigned(107,8) ,
4230	 => std_logic_vector(to_unsigned(107,8) ,
4231	 => std_logic_vector(to_unsigned(107,8) ,
4232	 => std_logic_vector(to_unsigned(108,8) ,
4233	 => std_logic_vector(to_unsigned(105,8) ,
4234	 => std_logic_vector(to_unsigned(104,8) ,
4235	 => std_logic_vector(to_unsigned(104,8) ,
4236	 => std_logic_vector(to_unsigned(100,8) ,
4237	 => std_logic_vector(to_unsigned(104,8) ,
4238	 => std_logic_vector(to_unsigned(101,8) ,
4239	 => std_logic_vector(to_unsigned(101,8) ,
4240	 => std_logic_vector(to_unsigned(97,8) ,
4241	 => std_logic_vector(to_unsigned(90,8) ,
4242	 => std_logic_vector(to_unsigned(91,8) ,
4243	 => std_logic_vector(to_unsigned(95,8) ,
4244	 => std_logic_vector(to_unsigned(96,8) ,
4245	 => std_logic_vector(to_unsigned(95,8) ,
4246	 => std_logic_vector(to_unsigned(95,8) ,
4247	 => std_logic_vector(to_unsigned(92,8) ,
4248	 => std_logic_vector(to_unsigned(91,8) ,
4249	 => std_logic_vector(to_unsigned(91,8) ,
4250	 => std_logic_vector(to_unsigned(88,8) ,
4251	 => std_logic_vector(to_unsigned(92,8) ,
4252	 => std_logic_vector(to_unsigned(90,8) ,
4253	 => std_logic_vector(to_unsigned(90,8) ,
4254	 => std_logic_vector(to_unsigned(87,8) ,
4255	 => std_logic_vector(to_unsigned(86,8) ,
4256	 => std_logic_vector(to_unsigned(82,8) ,
4257	 => std_logic_vector(to_unsigned(81,8) ,
4258	 => std_logic_vector(to_unsigned(81,8) ,
4259	 => std_logic_vector(to_unsigned(90,8) ,
4260	 => std_logic_vector(to_unsigned(90,8) ,
4261	 => std_logic_vector(to_unsigned(81,8) ,
4262	 => std_logic_vector(to_unsigned(84,8) ,
4263	 => std_logic_vector(to_unsigned(82,8) ,
4264	 => std_logic_vector(to_unsigned(80,8) ,
4265	 => std_logic_vector(to_unsigned(80,8) ,
4266	 => std_logic_vector(to_unsigned(80,8) ,
4267	 => std_logic_vector(to_unsigned(84,8) ,
4268	 => std_logic_vector(to_unsigned(81,8) ,
4269	 => std_logic_vector(to_unsigned(80,8) ,
4270	 => std_logic_vector(to_unsigned(80,8) ,
4271	 => std_logic_vector(to_unsigned(84,8) ,
4272	 => std_logic_vector(to_unsigned(87,8) ,
4273	 => std_logic_vector(to_unsigned(88,8) ,
4274	 => std_logic_vector(to_unsigned(86,8) ,
4275	 => std_logic_vector(to_unsigned(91,8) ,
4276	 => std_logic_vector(to_unsigned(85,8) ,
4277	 => std_logic_vector(to_unsigned(81,8) ,
4278	 => std_logic_vector(to_unsigned(90,8) ,
4279	 => std_logic_vector(to_unsigned(90,8) ,
4280	 => std_logic_vector(to_unsigned(91,8) ,
4281	 => std_logic_vector(to_unsigned(86,8) ,
4282	 => std_logic_vector(to_unsigned(90,8) ,
4283	 => std_logic_vector(to_unsigned(96,8) ,
4284	 => std_logic_vector(to_unsigned(90,8) ,
4285	 => std_logic_vector(to_unsigned(91,8) ,
4286	 => std_logic_vector(to_unsigned(88,8) ,
4287	 => std_logic_vector(to_unsigned(84,8) ,
4288	 => std_logic_vector(to_unsigned(84,8) ,
4289	 => std_logic_vector(to_unsigned(87,8) ,
4290	 => std_logic_vector(to_unsigned(92,8) ,
4291	 => std_logic_vector(to_unsigned(93,8) ,
4292	 => std_logic_vector(to_unsigned(93,8) ,
4293	 => std_logic_vector(to_unsigned(88,8) ,
4294	 => std_logic_vector(to_unsigned(88,8) ,
4295	 => std_logic_vector(to_unsigned(91,8) ,
4296	 => std_logic_vector(to_unsigned(93,8) ,
4297	 => std_logic_vector(to_unsigned(91,8) ,
4298	 => std_logic_vector(to_unsigned(92,8) ,
4299	 => std_logic_vector(to_unsigned(95,8) ,
4300	 => std_logic_vector(to_unsigned(95,8) ,
4301	 => std_logic_vector(to_unsigned(92,8) ,
4302	 => std_logic_vector(to_unsigned(99,8) ,
4303	 => std_logic_vector(to_unsigned(103,8) ,
4304	 => std_logic_vector(to_unsigned(97,8) ,
4305	 => std_logic_vector(to_unsigned(99,8) ,
4306	 => std_logic_vector(to_unsigned(96,8) ,
4307	 => std_logic_vector(to_unsigned(95,8) ,
4308	 => std_logic_vector(to_unsigned(92,8) ,
4309	 => std_logic_vector(to_unsigned(91,8) ,
4310	 => std_logic_vector(to_unsigned(86,8) ,
4311	 => std_logic_vector(to_unsigned(86,8) ,
4312	 => std_logic_vector(to_unsigned(90,8) ,
4313	 => std_logic_vector(to_unsigned(91,8) ,
4314	 => std_logic_vector(to_unsigned(85,8) ,
4315	 => std_logic_vector(to_unsigned(84,8) ,
4316	 => std_logic_vector(to_unsigned(86,8) ,
4317	 => std_logic_vector(to_unsigned(82,8) ,
4318	 => std_logic_vector(to_unsigned(76,8) ,
4319	 => std_logic_vector(to_unsigned(85,8) ,
4320	 => std_logic_vector(to_unsigned(88,8) ,
4321	 => std_logic_vector(to_unsigned(85,8) ,
4322	 => std_logic_vector(to_unsigned(84,8) ,
4323	 => std_logic_vector(to_unsigned(80,8) ,
4324	 => std_logic_vector(to_unsigned(85,8) ,
4325	 => std_logic_vector(to_unsigned(86,8) ,
4326	 => std_logic_vector(to_unsigned(82,8) ,
4327	 => std_logic_vector(to_unsigned(84,8) ,
4328	 => std_logic_vector(to_unsigned(82,8) ,
4329	 => std_logic_vector(to_unsigned(85,8) ,
4330	 => std_logic_vector(to_unsigned(82,8) ,
4331	 => std_logic_vector(to_unsigned(81,8) ,
4332	 => std_logic_vector(to_unsigned(84,8) ,
4333	 => std_logic_vector(to_unsigned(81,8) ,
4334	 => std_logic_vector(to_unsigned(79,8) ,
4335	 => std_logic_vector(to_unsigned(79,8) ,
4336	 => std_logic_vector(to_unsigned(82,8) ,
4337	 => std_logic_vector(to_unsigned(79,8) ,
4338	 => std_logic_vector(to_unsigned(80,8) ,
4339	 => std_logic_vector(to_unsigned(81,8) ,
4340	 => std_logic_vector(to_unsigned(77,8) ,
4341	 => std_logic_vector(to_unsigned(73,8) ,
4342	 => std_logic_vector(to_unsigned(74,8) ,
4343	 => std_logic_vector(to_unsigned(72,8) ,
4344	 => std_logic_vector(to_unsigned(67,8) ,
4345	 => std_logic_vector(to_unsigned(65,8) ,
4346	 => std_logic_vector(to_unsigned(63,8) ,
4347	 => std_logic_vector(to_unsigned(68,8) ,
4348	 => std_logic_vector(to_unsigned(69,8) ,
4349	 => std_logic_vector(to_unsigned(65,8) ,
4350	 => std_logic_vector(to_unsigned(70,8) ,
4351	 => std_logic_vector(to_unsigned(74,8) ,
4352	 => std_logic_vector(to_unsigned(79,8) ,
4353	 => std_logic_vector(to_unsigned(77,8) ,
4354	 => std_logic_vector(to_unsigned(69,8) ,
4355	 => std_logic_vector(to_unsigned(69,8) ,
4356	 => std_logic_vector(to_unsigned(71,8) ,
4357	 => std_logic_vector(to_unsigned(69,8) ,
4358	 => std_logic_vector(to_unsigned(70,8) ,
4359	 => std_logic_vector(to_unsigned(76,8) ,
4360	 => std_logic_vector(to_unsigned(74,8) ,
4361	 => std_logic_vector(to_unsigned(71,8) ,
4362	 => std_logic_vector(to_unsigned(73,8) ,
4363	 => std_logic_vector(to_unsigned(72,8) ,
4364	 => std_logic_vector(to_unsigned(74,8) ,
4365	 => std_logic_vector(to_unsigned(81,8) ,
4366	 => std_logic_vector(to_unsigned(81,8) ,
4367	 => std_logic_vector(to_unsigned(76,8) ,
4368	 => std_logic_vector(to_unsigned(82,8) ,
4369	 => std_logic_vector(to_unsigned(84,8) ,
4370	 => std_logic_vector(to_unsigned(86,8) ,
4371	 => std_logic_vector(to_unsigned(80,8) ,
4372	 => std_logic_vector(to_unsigned(78,8) ,
4373	 => std_logic_vector(to_unsigned(80,8) ,
4374	 => std_logic_vector(to_unsigned(80,8) ,
4375	 => std_logic_vector(to_unsigned(82,8) ,
4376	 => std_logic_vector(to_unsigned(84,8) ,
4377	 => std_logic_vector(to_unsigned(82,8) ,
4378	 => std_logic_vector(to_unsigned(82,8) ,
4379	 => std_logic_vector(to_unsigned(82,8) ,
4380	 => std_logic_vector(to_unsigned(80,8) ,
4381	 => std_logic_vector(to_unsigned(84,8) ,
4382	 => std_logic_vector(to_unsigned(85,8) ,
4383	 => std_logic_vector(to_unsigned(86,8) ,
4384	 => std_logic_vector(to_unsigned(81,8) ,
4385	 => std_logic_vector(to_unsigned(81,8) ,
4386	 => std_logic_vector(to_unsigned(86,8) ,
4387	 => std_logic_vector(to_unsigned(84,8) ,
4388	 => std_logic_vector(to_unsigned(85,8) ,
4389	 => std_logic_vector(to_unsigned(87,8) ,
4390	 => std_logic_vector(to_unsigned(72,8) ,
4391	 => std_logic_vector(to_unsigned(65,8) ,
4392	 => std_logic_vector(to_unsigned(78,8) ,
4393	 => std_logic_vector(to_unsigned(86,8) ,
4394	 => std_logic_vector(to_unsigned(86,8) ,
4395	 => std_logic_vector(to_unsigned(81,8) ,
4396	 => std_logic_vector(to_unsigned(84,8) ,
4397	 => std_logic_vector(to_unsigned(93,8) ,
4398	 => std_logic_vector(to_unsigned(31,8) ,
4399	 => std_logic_vector(to_unsigned(0,8) ,
4400	 => std_logic_vector(to_unsigned(0,8) ,
4401	 => std_logic_vector(to_unsigned(2,8) ,
4402	 => std_logic_vector(to_unsigned(63,8) ,
4403	 => std_logic_vector(to_unsigned(100,8) ,
4404	 => std_logic_vector(to_unsigned(87,8) ,
4405	 => std_logic_vector(to_unsigned(90,8) ,
4406	 => std_logic_vector(to_unsigned(93,8) ,
4407	 => std_logic_vector(to_unsigned(93,8) ,
4408	 => std_logic_vector(to_unsigned(100,8) ,
4409	 => std_logic_vector(to_unsigned(107,8) ,
4410	 => std_logic_vector(to_unsigned(108,8) ,
4411	 => std_logic_vector(to_unsigned(114,8) ,
4412	 => std_logic_vector(to_unsigned(116,8) ,
4413	 => std_logic_vector(to_unsigned(107,8) ,
4414	 => std_logic_vector(to_unsigned(103,8) ,
4415	 => std_logic_vector(to_unsigned(111,8) ,
4416	 => std_logic_vector(to_unsigned(109,8) ,
4417	 => std_logic_vector(to_unsigned(96,8) ,
4418	 => std_logic_vector(to_unsigned(90,8) ,
4419	 => std_logic_vector(to_unsigned(92,8) ,
4420	 => std_logic_vector(to_unsigned(96,8) ,
4421	 => std_logic_vector(to_unsigned(93,8) ,
4422	 => std_logic_vector(to_unsigned(95,8) ,
4423	 => std_logic_vector(to_unsigned(96,8) ,
4424	 => std_logic_vector(to_unsigned(101,8) ,
4425	 => std_logic_vector(to_unsigned(103,8) ,
4426	 => std_logic_vector(to_unsigned(96,8) ,
4427	 => std_logic_vector(to_unsigned(93,8) ,
4428	 => std_logic_vector(to_unsigned(100,8) ,
4429	 => std_logic_vector(to_unsigned(101,8) ,
4430	 => std_logic_vector(to_unsigned(96,8) ,
4431	 => std_logic_vector(to_unsigned(101,8) ,
4432	 => std_logic_vector(to_unsigned(109,8) ,
4433	 => std_logic_vector(to_unsigned(111,8) ,
4434	 => std_logic_vector(to_unsigned(105,8) ,
4435	 => std_logic_vector(to_unsigned(111,8) ,
4436	 => std_logic_vector(to_unsigned(116,8) ,
4437	 => std_logic_vector(to_unsigned(115,8) ,
4438	 => std_logic_vector(to_unsigned(115,8) ,
4439	 => std_logic_vector(to_unsigned(118,8) ,
4440	 => std_logic_vector(to_unsigned(119,8) ,
4441	 => std_logic_vector(to_unsigned(122,8) ,
4442	 => std_logic_vector(to_unsigned(128,8) ,
4443	 => std_logic_vector(to_unsigned(136,8) ,
4444	 => std_logic_vector(to_unsigned(127,8) ,
4445	 => std_logic_vector(to_unsigned(131,8) ,
4446	 => std_logic_vector(to_unsigned(144,8) ,
4447	 => std_logic_vector(to_unsigned(136,8) ,
4448	 => std_logic_vector(to_unsigned(125,8) ,
4449	 => std_logic_vector(to_unsigned(128,8) ,
4450	 => std_logic_vector(to_unsigned(133,8) ,
4451	 => std_logic_vector(to_unsigned(134,8) ,
4452	 => std_logic_vector(to_unsigned(138,8) ,
4453	 => std_logic_vector(to_unsigned(142,8) ,
4454	 => std_logic_vector(to_unsigned(141,8) ,
4455	 => std_logic_vector(to_unsigned(142,8) ,
4456	 => std_logic_vector(to_unsigned(146,8) ,
4457	 => std_logic_vector(to_unsigned(149,8) ,
4458	 => std_logic_vector(to_unsigned(154,8) ,
4459	 => std_logic_vector(to_unsigned(156,8) ,
4460	 => std_logic_vector(to_unsigned(154,8) ,
4461	 => std_logic_vector(to_unsigned(156,8) ,
4462	 => std_logic_vector(to_unsigned(157,8) ,
4463	 => std_logic_vector(to_unsigned(159,8) ,
4464	 => std_logic_vector(to_unsigned(161,8) ,
4465	 => std_logic_vector(to_unsigned(161,8) ,
4466	 => std_logic_vector(to_unsigned(161,8) ,
4467	 => std_logic_vector(to_unsigned(159,8) ,
4468	 => std_logic_vector(to_unsigned(159,8) ,
4469	 => std_logic_vector(to_unsigned(163,8) ,
4470	 => std_logic_vector(to_unsigned(161,8) ,
4471	 => std_logic_vector(to_unsigned(163,8) ,
4472	 => std_logic_vector(to_unsigned(161,8) ,
4473	 => std_logic_vector(to_unsigned(161,8) ,
4474	 => std_logic_vector(to_unsigned(161,8) ,
4475	 => std_logic_vector(to_unsigned(154,8) ,
4476	 => std_logic_vector(to_unsigned(156,8) ,
4477	 => std_logic_vector(to_unsigned(161,8) ,
4478	 => std_logic_vector(to_unsigned(163,8) ,
4479	 => std_logic_vector(to_unsigned(164,8) ,
4480	 => std_logic_vector(to_unsigned(163,8) ,
4481	 => std_logic_vector(to_unsigned(85,8) ,
4482	 => std_logic_vector(to_unsigned(85,8) ,
4483	 => std_logic_vector(to_unsigned(77,8) ,
4484	 => std_logic_vector(to_unsigned(81,8) ,
4485	 => std_logic_vector(to_unsigned(74,8) ,
4486	 => std_logic_vector(to_unsigned(80,8) ,
4487	 => std_logic_vector(to_unsigned(88,8) ,
4488	 => std_logic_vector(to_unsigned(79,8) ,
4489	 => std_logic_vector(to_unsigned(76,8) ,
4490	 => std_logic_vector(to_unsigned(72,8) ,
4491	 => std_logic_vector(to_unsigned(78,8) ,
4492	 => std_logic_vector(to_unsigned(80,8) ,
4493	 => std_logic_vector(to_unsigned(80,8) ,
4494	 => std_logic_vector(to_unsigned(77,8) ,
4495	 => std_logic_vector(to_unsigned(78,8) ,
4496	 => std_logic_vector(to_unsigned(81,8) ,
4497	 => std_logic_vector(to_unsigned(82,8) ,
4498	 => std_logic_vector(to_unsigned(79,8) ,
4499	 => std_logic_vector(to_unsigned(80,8) ,
4500	 => std_logic_vector(to_unsigned(84,8) ,
4501	 => std_logic_vector(to_unsigned(79,8) ,
4502	 => std_logic_vector(to_unsigned(81,8) ,
4503	 => std_logic_vector(to_unsigned(81,8) ,
4504	 => std_logic_vector(to_unsigned(78,8) ,
4505	 => std_logic_vector(to_unsigned(74,8) ,
4506	 => std_logic_vector(to_unsigned(76,8) ,
4507	 => std_logic_vector(to_unsigned(76,8) ,
4508	 => std_logic_vector(to_unsigned(80,8) ,
4509	 => std_logic_vector(to_unsigned(71,8) ,
4510	 => std_logic_vector(to_unsigned(73,8) ,
4511	 => std_logic_vector(to_unsigned(77,8) ,
4512	 => std_logic_vector(to_unsigned(78,8) ,
4513	 => std_logic_vector(to_unsigned(81,8) ,
4514	 => std_logic_vector(to_unsigned(84,8) ,
4515	 => std_logic_vector(to_unsigned(82,8) ,
4516	 => std_logic_vector(to_unsigned(78,8) ,
4517	 => std_logic_vector(to_unsigned(72,8) ,
4518	 => std_logic_vector(to_unsigned(78,8) ,
4519	 => std_logic_vector(to_unsigned(87,8) ,
4520	 => std_logic_vector(to_unsigned(86,8) ,
4521	 => std_logic_vector(to_unsigned(84,8) ,
4522	 => std_logic_vector(to_unsigned(87,8) ,
4523	 => std_logic_vector(to_unsigned(88,8) ,
4524	 => std_logic_vector(to_unsigned(92,8) ,
4525	 => std_logic_vector(to_unsigned(92,8) ,
4526	 => std_logic_vector(to_unsigned(96,8) ,
4527	 => std_logic_vector(to_unsigned(96,8) ,
4528	 => std_logic_vector(to_unsigned(97,8) ,
4529	 => std_logic_vector(to_unsigned(96,8) ,
4530	 => std_logic_vector(to_unsigned(100,8) ,
4531	 => std_logic_vector(to_unsigned(101,8) ,
4532	 => std_logic_vector(to_unsigned(100,8) ,
4533	 => std_logic_vector(to_unsigned(109,8) ,
4534	 => std_logic_vector(to_unsigned(111,8) ,
4535	 => std_logic_vector(to_unsigned(105,8) ,
4536	 => std_logic_vector(to_unsigned(107,8) ,
4537	 => std_logic_vector(to_unsigned(107,8) ,
4538	 => std_logic_vector(to_unsigned(109,8) ,
4539	 => std_logic_vector(to_unsigned(112,8) ,
4540	 => std_logic_vector(to_unsigned(115,8) ,
4541	 => std_logic_vector(to_unsigned(109,8) ,
4542	 => std_logic_vector(to_unsigned(105,8) ,
4543	 => std_logic_vector(to_unsigned(103,8) ,
4544	 => std_logic_vector(to_unsigned(103,8) ,
4545	 => std_logic_vector(to_unsigned(103,8) ,
4546	 => std_logic_vector(to_unsigned(109,8) ,
4547	 => std_logic_vector(to_unsigned(111,8) ,
4548	 => std_logic_vector(to_unsigned(108,8) ,
4549	 => std_logic_vector(to_unsigned(105,8) ,
4550	 => std_logic_vector(to_unsigned(104,8) ,
4551	 => std_logic_vector(to_unsigned(105,8) ,
4552	 => std_logic_vector(to_unsigned(105,8) ,
4553	 => std_logic_vector(to_unsigned(104,8) ,
4554	 => std_logic_vector(to_unsigned(105,8) ,
4555	 => std_logic_vector(to_unsigned(104,8) ,
4556	 => std_logic_vector(to_unsigned(96,8) ,
4557	 => std_logic_vector(to_unsigned(99,8) ,
4558	 => std_logic_vector(to_unsigned(99,8) ,
4559	 => std_logic_vector(to_unsigned(99,8) ,
4560	 => std_logic_vector(to_unsigned(92,8) ,
4561	 => std_logic_vector(to_unsigned(86,8) ,
4562	 => std_logic_vector(to_unsigned(87,8) ,
4563	 => std_logic_vector(to_unsigned(85,8) ,
4564	 => std_logic_vector(to_unsigned(86,8) ,
4565	 => std_logic_vector(to_unsigned(90,8) ,
4566	 => std_logic_vector(to_unsigned(87,8) ,
4567	 => std_logic_vector(to_unsigned(86,8) ,
4568	 => std_logic_vector(to_unsigned(82,8) ,
4569	 => std_logic_vector(to_unsigned(87,8) ,
4570	 => std_logic_vector(to_unsigned(87,8) ,
4571	 => std_logic_vector(to_unsigned(88,8) ,
4572	 => std_logic_vector(to_unsigned(90,8) ,
4573	 => std_logic_vector(to_unsigned(88,8) ,
4574	 => std_logic_vector(to_unsigned(82,8) ,
4575	 => std_logic_vector(to_unsigned(85,8) ,
4576	 => std_logic_vector(to_unsigned(85,8) ,
4577	 => std_logic_vector(to_unsigned(85,8) ,
4578	 => std_logic_vector(to_unsigned(82,8) ,
4579	 => std_logic_vector(to_unsigned(85,8) ,
4580	 => std_logic_vector(to_unsigned(81,8) ,
4581	 => std_logic_vector(to_unsigned(80,8) ,
4582	 => std_logic_vector(to_unsigned(80,8) ,
4583	 => std_logic_vector(to_unsigned(77,8) ,
4584	 => std_logic_vector(to_unsigned(80,8) ,
4585	 => std_logic_vector(to_unsigned(79,8) ,
4586	 => std_logic_vector(to_unsigned(79,8) ,
4587	 => std_logic_vector(to_unsigned(79,8) ,
4588	 => std_logic_vector(to_unsigned(81,8) ,
4589	 => std_logic_vector(to_unsigned(79,8) ,
4590	 => std_logic_vector(to_unsigned(74,8) ,
4591	 => std_logic_vector(to_unsigned(76,8) ,
4592	 => std_logic_vector(to_unsigned(76,8) ,
4593	 => std_logic_vector(to_unsigned(80,8) ,
4594	 => std_logic_vector(to_unsigned(81,8) ,
4595	 => std_logic_vector(to_unsigned(85,8) ,
4596	 => std_logic_vector(to_unsigned(85,8) ,
4597	 => std_logic_vector(to_unsigned(85,8) ,
4598	 => std_logic_vector(to_unsigned(91,8) ,
4599	 => std_logic_vector(to_unsigned(87,8) ,
4600	 => std_logic_vector(to_unsigned(91,8) ,
4601	 => std_logic_vector(to_unsigned(88,8) ,
4602	 => std_logic_vector(to_unsigned(90,8) ,
4603	 => std_logic_vector(to_unsigned(90,8) ,
4604	 => std_logic_vector(to_unsigned(84,8) ,
4605	 => std_logic_vector(to_unsigned(88,8) ,
4606	 => std_logic_vector(to_unsigned(87,8) ,
4607	 => std_logic_vector(to_unsigned(82,8) ,
4608	 => std_logic_vector(to_unsigned(82,8) ,
4609	 => std_logic_vector(to_unsigned(86,8) ,
4610	 => std_logic_vector(to_unsigned(91,8) ,
4611	 => std_logic_vector(to_unsigned(92,8) ,
4612	 => std_logic_vector(to_unsigned(91,8) ,
4613	 => std_logic_vector(to_unsigned(90,8) ,
4614	 => std_logic_vector(to_unsigned(93,8) ,
4615	 => std_logic_vector(to_unsigned(95,8) ,
4616	 => std_logic_vector(to_unsigned(92,8) ,
4617	 => std_logic_vector(to_unsigned(90,8) ,
4618	 => std_logic_vector(to_unsigned(93,8) ,
4619	 => std_logic_vector(to_unsigned(99,8) ,
4620	 => std_logic_vector(to_unsigned(95,8) ,
4621	 => std_logic_vector(to_unsigned(92,8) ,
4622	 => std_logic_vector(to_unsigned(97,8) ,
4623	 => std_logic_vector(to_unsigned(103,8) ,
4624	 => std_logic_vector(to_unsigned(97,8) ,
4625	 => std_logic_vector(to_unsigned(101,8) ,
4626	 => std_logic_vector(to_unsigned(97,8) ,
4627	 => std_logic_vector(to_unsigned(92,8) ,
4628	 => std_logic_vector(to_unsigned(95,8) ,
4629	 => std_logic_vector(to_unsigned(100,8) ,
4630	 => std_logic_vector(to_unsigned(95,8) ,
4631	 => std_logic_vector(to_unsigned(93,8) ,
4632	 => std_logic_vector(to_unsigned(92,8) ,
4633	 => std_logic_vector(to_unsigned(86,8) ,
4634	 => std_logic_vector(to_unsigned(88,8) ,
4635	 => std_logic_vector(to_unsigned(91,8) ,
4636	 => std_logic_vector(to_unsigned(90,8) ,
4637	 => std_logic_vector(to_unsigned(87,8) ,
4638	 => std_logic_vector(to_unsigned(80,8) ,
4639	 => std_logic_vector(to_unsigned(87,8) ,
4640	 => std_logic_vector(to_unsigned(91,8) ,
4641	 => std_logic_vector(to_unsigned(88,8) ,
4642	 => std_logic_vector(to_unsigned(87,8) ,
4643	 => std_logic_vector(to_unsigned(86,8) ,
4644	 => std_logic_vector(to_unsigned(85,8) ,
4645	 => std_logic_vector(to_unsigned(85,8) ,
4646	 => std_logic_vector(to_unsigned(86,8) ,
4647	 => std_logic_vector(to_unsigned(85,8) ,
4648	 => std_logic_vector(to_unsigned(82,8) ,
4649	 => std_logic_vector(to_unsigned(84,8) ,
4650	 => std_logic_vector(to_unsigned(80,8) ,
4651	 => std_logic_vector(to_unsigned(84,8) ,
4652	 => std_logic_vector(to_unsigned(86,8) ,
4653	 => std_logic_vector(to_unsigned(84,8) ,
4654	 => std_logic_vector(to_unsigned(85,8) ,
4655	 => std_logic_vector(to_unsigned(82,8) ,
4656	 => std_logic_vector(to_unsigned(80,8) ,
4657	 => std_logic_vector(to_unsigned(80,8) ,
4658	 => std_logic_vector(to_unsigned(80,8) ,
4659	 => std_logic_vector(to_unsigned(82,8) ,
4660	 => std_logic_vector(to_unsigned(80,8) ,
4661	 => std_logic_vector(to_unsigned(71,8) ,
4662	 => std_logic_vector(to_unsigned(70,8) ,
4663	 => std_logic_vector(to_unsigned(70,8) ,
4664	 => std_logic_vector(to_unsigned(68,8) ,
4665	 => std_logic_vector(to_unsigned(72,8) ,
4666	 => std_logic_vector(to_unsigned(70,8) ,
4667	 => std_logic_vector(to_unsigned(66,8) ,
4668	 => std_logic_vector(to_unsigned(64,8) ,
4669	 => std_logic_vector(to_unsigned(66,8) ,
4670	 => std_logic_vector(to_unsigned(70,8) ,
4671	 => std_logic_vector(to_unsigned(72,8) ,
4672	 => std_logic_vector(to_unsigned(71,8) ,
4673	 => std_logic_vector(to_unsigned(67,8) ,
4674	 => std_logic_vector(to_unsigned(69,8) ,
4675	 => std_logic_vector(to_unsigned(71,8) ,
4676	 => std_logic_vector(to_unsigned(68,8) ,
4677	 => std_logic_vector(to_unsigned(68,8) ,
4678	 => std_logic_vector(to_unsigned(71,8) ,
4679	 => std_logic_vector(to_unsigned(73,8) ,
4680	 => std_logic_vector(to_unsigned(74,8) ,
4681	 => std_logic_vector(to_unsigned(73,8) ,
4682	 => std_logic_vector(to_unsigned(72,8) ,
4683	 => std_logic_vector(to_unsigned(72,8) ,
4684	 => std_logic_vector(to_unsigned(76,8) ,
4685	 => std_logic_vector(to_unsigned(79,8) ,
4686	 => std_logic_vector(to_unsigned(77,8) ,
4687	 => std_logic_vector(to_unsigned(81,8) ,
4688	 => std_logic_vector(to_unsigned(85,8) ,
4689	 => std_logic_vector(to_unsigned(85,8) ,
4690	 => std_logic_vector(to_unsigned(86,8) ,
4691	 => std_logic_vector(to_unsigned(87,8) ,
4692	 => std_logic_vector(to_unsigned(81,8) ,
4693	 => std_logic_vector(to_unsigned(85,8) ,
4694	 => std_logic_vector(to_unsigned(87,8) ,
4695	 => std_logic_vector(to_unsigned(82,8) ,
4696	 => std_logic_vector(to_unsigned(81,8) ,
4697	 => std_logic_vector(to_unsigned(84,8) ,
4698	 => std_logic_vector(to_unsigned(85,8) ,
4699	 => std_logic_vector(to_unsigned(86,8) ,
4700	 => std_logic_vector(to_unsigned(88,8) ,
4701	 => std_logic_vector(to_unsigned(84,8) ,
4702	 => std_logic_vector(to_unsigned(82,8) ,
4703	 => std_logic_vector(to_unsigned(81,8) ,
4704	 => std_logic_vector(to_unsigned(85,8) ,
4705	 => std_logic_vector(to_unsigned(87,8) ,
4706	 => std_logic_vector(to_unsigned(87,8) ,
4707	 => std_logic_vector(to_unsigned(91,8) ,
4708	 => std_logic_vector(to_unsigned(90,8) ,
4709	 => std_logic_vector(to_unsigned(88,8) ,
4710	 => std_logic_vector(to_unsigned(74,8) ,
4711	 => std_logic_vector(to_unsigned(68,8) ,
4712	 => std_logic_vector(to_unsigned(80,8) ,
4713	 => std_logic_vector(to_unsigned(88,8) ,
4714	 => std_logic_vector(to_unsigned(90,8) ,
4715	 => std_logic_vector(to_unsigned(81,8) ,
4716	 => std_logic_vector(to_unsigned(82,8) ,
4717	 => std_logic_vector(to_unsigned(90,8) ,
4718	 => std_logic_vector(to_unsigned(53,8) ,
4719	 => std_logic_vector(to_unsigned(2,8) ,
4720	 => std_logic_vector(to_unsigned(0,8) ,
4721	 => std_logic_vector(to_unsigned(1,8) ,
4722	 => std_logic_vector(to_unsigned(41,8) ,
4723	 => std_logic_vector(to_unsigned(101,8) ,
4724	 => std_logic_vector(to_unsigned(82,8) ,
4725	 => std_logic_vector(to_unsigned(88,8) ,
4726	 => std_logic_vector(to_unsigned(93,8) ,
4727	 => std_logic_vector(to_unsigned(96,8) ,
4728	 => std_logic_vector(to_unsigned(99,8) ,
4729	 => std_logic_vector(to_unsigned(101,8) ,
4730	 => std_logic_vector(to_unsigned(107,8) ,
4731	 => std_logic_vector(to_unsigned(111,8) ,
4732	 => std_logic_vector(to_unsigned(105,8) ,
4733	 => std_logic_vector(to_unsigned(101,8) ,
4734	 => std_logic_vector(to_unsigned(101,8) ,
4735	 => std_logic_vector(to_unsigned(99,8) ,
4736	 => std_logic_vector(to_unsigned(103,8) ,
4737	 => std_logic_vector(to_unsigned(95,8) ,
4738	 => std_logic_vector(to_unsigned(91,8) ,
4739	 => std_logic_vector(to_unsigned(97,8) ,
4740	 => std_logic_vector(to_unsigned(96,8) ,
4741	 => std_logic_vector(to_unsigned(92,8) ,
4742	 => std_logic_vector(to_unsigned(90,8) ,
4743	 => std_logic_vector(to_unsigned(92,8) ,
4744	 => std_logic_vector(to_unsigned(96,8) ,
4745	 => std_logic_vector(to_unsigned(96,8) ,
4746	 => std_logic_vector(to_unsigned(99,8) ,
4747	 => std_logic_vector(to_unsigned(96,8) ,
4748	 => std_logic_vector(to_unsigned(104,8) ,
4749	 => std_logic_vector(to_unsigned(103,8) ,
4750	 => std_logic_vector(to_unsigned(97,8) ,
4751	 => std_logic_vector(to_unsigned(107,8) ,
4752	 => std_logic_vector(to_unsigned(105,8) ,
4753	 => std_logic_vector(to_unsigned(109,8) ,
4754	 => std_logic_vector(to_unsigned(107,8) ,
4755	 => std_logic_vector(to_unsigned(105,8) ,
4756	 => std_logic_vector(to_unsigned(109,8) ,
4757	 => std_logic_vector(to_unsigned(112,8) ,
4758	 => std_logic_vector(to_unsigned(111,8) ,
4759	 => std_logic_vector(to_unsigned(114,8) ,
4760	 => std_logic_vector(to_unsigned(121,8) ,
4761	 => std_logic_vector(to_unsigned(125,8) ,
4762	 => std_logic_vector(to_unsigned(122,8) ,
4763	 => std_logic_vector(to_unsigned(125,8) ,
4764	 => std_logic_vector(to_unsigned(130,8) ,
4765	 => std_logic_vector(to_unsigned(134,8) ,
4766	 => std_logic_vector(to_unsigned(136,8) ,
4767	 => std_logic_vector(to_unsigned(138,8) ,
4768	 => std_logic_vector(to_unsigned(136,8) ,
4769	 => std_logic_vector(to_unsigned(127,8) ,
4770	 => std_logic_vector(to_unsigned(122,8) ,
4771	 => std_logic_vector(to_unsigned(127,8) ,
4772	 => std_logic_vector(to_unsigned(133,8) ,
4773	 => std_logic_vector(to_unsigned(136,8) ,
4774	 => std_logic_vector(to_unsigned(136,8) ,
4775	 => std_logic_vector(to_unsigned(139,8) ,
4776	 => std_logic_vector(to_unsigned(146,8) ,
4777	 => std_logic_vector(to_unsigned(144,8) ,
4778	 => std_logic_vector(to_unsigned(147,8) ,
4779	 => std_logic_vector(to_unsigned(154,8) ,
4780	 => std_logic_vector(to_unsigned(156,8) ,
4781	 => std_logic_vector(to_unsigned(156,8) ,
4782	 => std_logic_vector(to_unsigned(157,8) ,
4783	 => std_logic_vector(to_unsigned(157,8) ,
4784	 => std_logic_vector(to_unsigned(159,8) ,
4785	 => std_logic_vector(to_unsigned(159,8) ,
4786	 => std_logic_vector(to_unsigned(159,8) ,
4787	 => std_logic_vector(to_unsigned(159,8) ,
4788	 => std_logic_vector(to_unsigned(161,8) ,
4789	 => std_logic_vector(to_unsigned(164,8) ,
4790	 => std_logic_vector(to_unsigned(161,8) ,
4791	 => std_logic_vector(to_unsigned(159,8) ,
4792	 => std_logic_vector(to_unsigned(163,8) ,
4793	 => std_logic_vector(to_unsigned(161,8) ,
4794	 => std_logic_vector(to_unsigned(157,8) ,
4795	 => std_logic_vector(to_unsigned(157,8) ,
4796	 => std_logic_vector(to_unsigned(159,8) ,
4797	 => std_logic_vector(to_unsigned(157,8) ,
4798	 => std_logic_vector(to_unsigned(157,8) ,
4799	 => std_logic_vector(to_unsigned(163,8) ,
4800	 => std_logic_vector(to_unsigned(161,8) ,
4801	 => std_logic_vector(to_unsigned(79,8) ,
4802	 => std_logic_vector(to_unsigned(80,8) ,
4803	 => std_logic_vector(to_unsigned(78,8) ,
4804	 => std_logic_vector(to_unsigned(71,8) ,
4805	 => std_logic_vector(to_unsigned(70,8) ,
4806	 => std_logic_vector(to_unsigned(80,8) ,
4807	 => std_logic_vector(to_unsigned(77,8) ,
4808	 => std_logic_vector(to_unsigned(73,8) ,
4809	 => std_logic_vector(to_unsigned(77,8) ,
4810	 => std_logic_vector(to_unsigned(73,8) ,
4811	 => std_logic_vector(to_unsigned(70,8) ,
4812	 => std_logic_vector(to_unsigned(71,8) ,
4813	 => std_logic_vector(to_unsigned(77,8) ,
4814	 => std_logic_vector(to_unsigned(74,8) ,
4815	 => std_logic_vector(to_unsigned(69,8) ,
4816	 => std_logic_vector(to_unsigned(71,8) ,
4817	 => std_logic_vector(to_unsigned(77,8) ,
4818	 => std_logic_vector(to_unsigned(77,8) ,
4819	 => std_logic_vector(to_unsigned(74,8) ,
4820	 => std_logic_vector(to_unsigned(77,8) ,
4821	 => std_logic_vector(to_unsigned(73,8) ,
4822	 => std_logic_vector(to_unsigned(78,8) ,
4823	 => std_logic_vector(to_unsigned(82,8) ,
4824	 => std_logic_vector(to_unsigned(73,8) ,
4825	 => std_logic_vector(to_unsigned(72,8) ,
4826	 => std_logic_vector(to_unsigned(77,8) ,
4827	 => std_logic_vector(to_unsigned(72,8) ,
4828	 => std_logic_vector(to_unsigned(69,8) ,
4829	 => std_logic_vector(to_unsigned(71,8) ,
4830	 => std_logic_vector(to_unsigned(76,8) ,
4831	 => std_logic_vector(to_unsigned(74,8) ,
4832	 => std_logic_vector(to_unsigned(76,8) ,
4833	 => std_logic_vector(to_unsigned(80,8) ,
4834	 => std_logic_vector(to_unsigned(76,8) ,
4835	 => std_logic_vector(to_unsigned(72,8) ,
4836	 => std_logic_vector(to_unsigned(78,8) ,
4837	 => std_logic_vector(to_unsigned(73,8) ,
4838	 => std_logic_vector(to_unsigned(73,8) ,
4839	 => std_logic_vector(to_unsigned(81,8) ,
4840	 => std_logic_vector(to_unsigned(84,8) ,
4841	 => std_logic_vector(to_unsigned(79,8) ,
4842	 => std_logic_vector(to_unsigned(79,8) ,
4843	 => std_logic_vector(to_unsigned(81,8) ,
4844	 => std_logic_vector(to_unsigned(87,8) ,
4845	 => std_logic_vector(to_unsigned(91,8) ,
4846	 => std_logic_vector(to_unsigned(90,8) ,
4847	 => std_logic_vector(to_unsigned(93,8) ,
4848	 => std_logic_vector(to_unsigned(93,8) ,
4849	 => std_logic_vector(to_unsigned(90,8) ,
4850	 => std_logic_vector(to_unsigned(93,8) ,
4851	 => std_logic_vector(to_unsigned(97,8) ,
4852	 => std_logic_vector(to_unsigned(100,8) ,
4853	 => std_logic_vector(to_unsigned(107,8) ,
4854	 => std_logic_vector(to_unsigned(112,8) ,
4855	 => std_logic_vector(to_unsigned(112,8) ,
4856	 => std_logic_vector(to_unsigned(108,8) ,
4857	 => std_logic_vector(to_unsigned(109,8) ,
4858	 => std_logic_vector(to_unsigned(107,8) ,
4859	 => std_logic_vector(to_unsigned(101,8) ,
4860	 => std_logic_vector(to_unsigned(109,8) ,
4861	 => std_logic_vector(to_unsigned(109,8) ,
4862	 => std_logic_vector(to_unsigned(108,8) ,
4863	 => std_logic_vector(to_unsigned(105,8) ,
4864	 => std_logic_vector(to_unsigned(104,8) ,
4865	 => std_logic_vector(to_unsigned(105,8) ,
4866	 => std_logic_vector(to_unsigned(107,8) ,
4867	 => std_logic_vector(to_unsigned(109,8) ,
4868	 => std_logic_vector(to_unsigned(115,8) ,
4869	 => std_logic_vector(to_unsigned(112,8) ,
4870	 => std_logic_vector(to_unsigned(114,8) ,
4871	 => std_logic_vector(to_unsigned(112,8) ,
4872	 => std_logic_vector(to_unsigned(105,8) ,
4873	 => std_logic_vector(to_unsigned(104,8) ,
4874	 => std_logic_vector(to_unsigned(111,8) ,
4875	 => std_logic_vector(to_unsigned(112,8) ,
4876	 => std_logic_vector(to_unsigned(104,8) ,
4877	 => std_logic_vector(to_unsigned(95,8) ,
4878	 => std_logic_vector(to_unsigned(100,8) ,
4879	 => std_logic_vector(to_unsigned(96,8) ,
4880	 => std_logic_vector(to_unsigned(91,8) ,
4881	 => std_logic_vector(to_unsigned(90,8) ,
4882	 => std_logic_vector(to_unsigned(88,8) ,
4883	 => std_logic_vector(to_unsigned(87,8) ,
4884	 => std_logic_vector(to_unsigned(88,8) ,
4885	 => std_logic_vector(to_unsigned(90,8) ,
4886	 => std_logic_vector(to_unsigned(85,8) ,
4887	 => std_logic_vector(to_unsigned(81,8) ,
4888	 => std_logic_vector(to_unsigned(82,8) ,
4889	 => std_logic_vector(to_unsigned(85,8) ,
4890	 => std_logic_vector(to_unsigned(85,8) ,
4891	 => std_logic_vector(to_unsigned(85,8) ,
4892	 => std_logic_vector(to_unsigned(82,8) ,
4893	 => std_logic_vector(to_unsigned(80,8) ,
4894	 => std_logic_vector(to_unsigned(82,8) ,
4895	 => std_logic_vector(to_unsigned(87,8) ,
4896	 => std_logic_vector(to_unsigned(81,8) ,
4897	 => std_logic_vector(to_unsigned(80,8) ,
4898	 => std_logic_vector(to_unsigned(79,8) ,
4899	 => std_logic_vector(to_unsigned(78,8) ,
4900	 => std_logic_vector(to_unsigned(77,8) ,
4901	 => std_logic_vector(to_unsigned(84,8) ,
4902	 => std_logic_vector(to_unsigned(80,8) ,
4903	 => std_logic_vector(to_unsigned(78,8) ,
4904	 => std_logic_vector(to_unsigned(80,8) ,
4905	 => std_logic_vector(to_unsigned(77,8) ,
4906	 => std_logic_vector(to_unsigned(79,8) ,
4907	 => std_logic_vector(to_unsigned(77,8) ,
4908	 => std_logic_vector(to_unsigned(78,8) ,
4909	 => std_logic_vector(to_unsigned(76,8) ,
4910	 => std_logic_vector(to_unsigned(73,8) ,
4911	 => std_logic_vector(to_unsigned(72,8) ,
4912	 => std_logic_vector(to_unsigned(74,8) ,
4913	 => std_logic_vector(to_unsigned(76,8) ,
4914	 => std_logic_vector(to_unsigned(80,8) ,
4915	 => std_logic_vector(to_unsigned(87,8) ,
4916	 => std_logic_vector(to_unsigned(86,8) ,
4917	 => std_logic_vector(to_unsigned(85,8) ,
4918	 => std_logic_vector(to_unsigned(87,8) ,
4919	 => std_logic_vector(to_unsigned(87,8) ,
4920	 => std_logic_vector(to_unsigned(86,8) ,
4921	 => std_logic_vector(to_unsigned(93,8) ,
4922	 => std_logic_vector(to_unsigned(96,8) ,
4923	 => std_logic_vector(to_unsigned(90,8) ,
4924	 => std_logic_vector(to_unsigned(91,8) ,
4925	 => std_logic_vector(to_unsigned(91,8) ,
4926	 => std_logic_vector(to_unsigned(88,8) ,
4927	 => std_logic_vector(to_unsigned(86,8) ,
4928	 => std_logic_vector(to_unsigned(87,8) ,
4929	 => std_logic_vector(to_unsigned(91,8) ,
4930	 => std_logic_vector(to_unsigned(92,8) ,
4931	 => std_logic_vector(to_unsigned(90,8) ,
4932	 => std_logic_vector(to_unsigned(88,8) ,
4933	 => std_logic_vector(to_unsigned(87,8) ,
4934	 => std_logic_vector(to_unsigned(91,8) ,
4935	 => std_logic_vector(to_unsigned(95,8) ,
4936	 => std_logic_vector(to_unsigned(95,8) ,
4937	 => std_logic_vector(to_unsigned(92,8) ,
4938	 => std_logic_vector(to_unsigned(91,8) ,
4939	 => std_logic_vector(to_unsigned(96,8) ,
4940	 => std_logic_vector(to_unsigned(95,8) ,
4941	 => std_logic_vector(to_unsigned(95,8) ,
4942	 => std_logic_vector(to_unsigned(97,8) ,
4943	 => std_logic_vector(to_unsigned(99,8) ,
4944	 => std_logic_vector(to_unsigned(100,8) ,
4945	 => std_logic_vector(to_unsigned(103,8) ,
4946	 => std_logic_vector(to_unsigned(99,8) ,
4947	 => std_logic_vector(to_unsigned(95,8) ,
4948	 => std_logic_vector(to_unsigned(91,8) ,
4949	 => std_logic_vector(to_unsigned(101,8) ,
4950	 => std_logic_vector(to_unsigned(101,8) ,
4951	 => std_logic_vector(to_unsigned(92,8) ,
4952	 => std_logic_vector(to_unsigned(93,8) ,
4953	 => std_logic_vector(to_unsigned(90,8) ,
4954	 => std_logic_vector(to_unsigned(90,8) ,
4955	 => std_logic_vector(to_unsigned(96,8) ,
4956	 => std_logic_vector(to_unsigned(92,8) ,
4957	 => std_logic_vector(to_unsigned(90,8) ,
4958	 => std_logic_vector(to_unsigned(91,8) ,
4959	 => std_logic_vector(to_unsigned(86,8) ,
4960	 => std_logic_vector(to_unsigned(85,8) ,
4961	 => std_logic_vector(to_unsigned(88,8) ,
4962	 => std_logic_vector(to_unsigned(80,8) ,
4963	 => std_logic_vector(to_unsigned(84,8) ,
4964	 => std_logic_vector(to_unsigned(87,8) ,
4965	 => std_logic_vector(to_unsigned(84,8) ,
4966	 => std_logic_vector(to_unsigned(85,8) ,
4967	 => std_logic_vector(to_unsigned(85,8) ,
4968	 => std_logic_vector(to_unsigned(84,8) ,
4969	 => std_logic_vector(to_unsigned(87,8) ,
4970	 => std_logic_vector(to_unsigned(81,8) ,
4971	 => std_logic_vector(to_unsigned(81,8) ,
4972	 => std_logic_vector(to_unsigned(82,8) ,
4973	 => std_logic_vector(to_unsigned(84,8) ,
4974	 => std_logic_vector(to_unsigned(84,8) ,
4975	 => std_logic_vector(to_unsigned(77,8) ,
4976	 => std_logic_vector(to_unsigned(78,8) ,
4977	 => std_logic_vector(to_unsigned(79,8) ,
4978	 => std_logic_vector(to_unsigned(74,8) ,
4979	 => std_logic_vector(to_unsigned(78,8) ,
4980	 => std_logic_vector(to_unsigned(81,8) ,
4981	 => std_logic_vector(to_unsigned(76,8) ,
4982	 => std_logic_vector(to_unsigned(77,8) ,
4983	 => std_logic_vector(to_unsigned(70,8) ,
4984	 => std_logic_vector(to_unsigned(68,8) ,
4985	 => std_logic_vector(to_unsigned(71,8) ,
4986	 => std_logic_vector(to_unsigned(72,8) ,
4987	 => std_logic_vector(to_unsigned(74,8) ,
4988	 => std_logic_vector(to_unsigned(73,8) ,
4989	 => std_logic_vector(to_unsigned(72,8) ,
4990	 => std_logic_vector(to_unsigned(74,8) ,
4991	 => std_logic_vector(to_unsigned(78,8) ,
4992	 => std_logic_vector(to_unsigned(76,8) ,
4993	 => std_logic_vector(to_unsigned(77,8) ,
4994	 => std_logic_vector(to_unsigned(77,8) ,
4995	 => std_logic_vector(to_unsigned(76,8) ,
4996	 => std_logic_vector(to_unsigned(77,8) ,
4997	 => std_logic_vector(to_unsigned(74,8) ,
4998	 => std_logic_vector(to_unsigned(71,8) ,
4999	 => std_logic_vector(to_unsigned(72,8) ,
5000	 => std_logic_vector(to_unsigned(77,8) ,
5001	 => std_logic_vector(to_unsigned(80,8) ,
5002	 => std_logic_vector(to_unsigned(79,8) ,
5003	 => std_logic_vector(to_unsigned(70,8) ,
5004	 => std_logic_vector(to_unsigned(77,8) ,
5005	 => std_logic_vector(to_unsigned(81,8) ,
5006	 => std_logic_vector(to_unsigned(80,8) ,
5007	 => std_logic_vector(to_unsigned(82,8) ,
5008	 => std_logic_vector(to_unsigned(80,8) ,
5009	 => std_logic_vector(to_unsigned(82,8) ,
5010	 => std_logic_vector(to_unsigned(79,8) ,
5011	 => std_logic_vector(to_unsigned(85,8) ,
5012	 => std_logic_vector(to_unsigned(88,8) ,
5013	 => std_logic_vector(to_unsigned(85,8) ,
5014	 => std_logic_vector(to_unsigned(86,8) ,
5015	 => std_logic_vector(to_unsigned(87,8) ,
5016	 => std_logic_vector(to_unsigned(82,8) ,
5017	 => std_logic_vector(to_unsigned(87,8) ,
5018	 => std_logic_vector(to_unsigned(87,8) ,
5019	 => std_logic_vector(to_unsigned(85,8) ,
5020	 => std_logic_vector(to_unsigned(86,8) ,
5021	 => std_logic_vector(to_unsigned(84,8) ,
5022	 => std_logic_vector(to_unsigned(86,8) ,
5023	 => std_logic_vector(to_unsigned(85,8) ,
5024	 => std_logic_vector(to_unsigned(82,8) ,
5025	 => std_logic_vector(to_unsigned(86,8) ,
5026	 => std_logic_vector(to_unsigned(85,8) ,
5027	 => std_logic_vector(to_unsigned(88,8) ,
5028	 => std_logic_vector(to_unsigned(82,8) ,
5029	 => std_logic_vector(to_unsigned(86,8) ,
5030	 => std_logic_vector(to_unsigned(77,8) ,
5031	 => std_logic_vector(to_unsigned(71,8) ,
5032	 => std_logic_vector(to_unsigned(84,8) ,
5033	 => std_logic_vector(to_unsigned(91,8) ,
5034	 => std_logic_vector(to_unsigned(90,8) ,
5035	 => std_logic_vector(to_unsigned(84,8) ,
5036	 => std_logic_vector(to_unsigned(77,8) ,
5037	 => std_logic_vector(to_unsigned(82,8) ,
5038	 => std_logic_vector(to_unsigned(73,8) ,
5039	 => std_logic_vector(to_unsigned(8,8) ,
5040	 => std_logic_vector(to_unsigned(0,8) ,
5041	 => std_logic_vector(to_unsigned(0,8) ,
5042	 => std_logic_vector(to_unsigned(21,8) ,
5043	 => std_logic_vector(to_unsigned(96,8) ,
5044	 => std_logic_vector(to_unsigned(85,8) ,
5045	 => std_logic_vector(to_unsigned(84,8) ,
5046	 => std_logic_vector(to_unsigned(92,8) ,
5047	 => std_logic_vector(to_unsigned(96,8) ,
5048	 => std_logic_vector(to_unsigned(99,8) ,
5049	 => std_logic_vector(to_unsigned(96,8) ,
5050	 => std_logic_vector(to_unsigned(103,8) ,
5051	 => std_logic_vector(to_unsigned(105,8) ,
5052	 => std_logic_vector(to_unsigned(118,8) ,
5053	 => std_logic_vector(to_unsigned(114,8) ,
5054	 => std_logic_vector(to_unsigned(100,8) ,
5055	 => std_logic_vector(to_unsigned(95,8) ,
5056	 => std_logic_vector(to_unsigned(90,8) ,
5057	 => std_logic_vector(to_unsigned(88,8) ,
5058	 => std_logic_vector(to_unsigned(91,8) ,
5059	 => std_logic_vector(to_unsigned(90,8) ,
5060	 => std_logic_vector(to_unsigned(90,8) ,
5061	 => std_logic_vector(to_unsigned(96,8) ,
5062	 => std_logic_vector(to_unsigned(93,8) ,
5063	 => std_logic_vector(to_unsigned(96,8) ,
5064	 => std_logic_vector(to_unsigned(92,8) ,
5065	 => std_logic_vector(to_unsigned(92,8) ,
5066	 => std_logic_vector(to_unsigned(93,8) ,
5067	 => std_logic_vector(to_unsigned(90,8) ,
5068	 => std_logic_vector(to_unsigned(90,8) ,
5069	 => std_logic_vector(to_unsigned(91,8) ,
5070	 => std_logic_vector(to_unsigned(96,8) ,
5071	 => std_logic_vector(to_unsigned(103,8) ,
5072	 => std_logic_vector(to_unsigned(97,8) ,
5073	 => std_logic_vector(to_unsigned(99,8) ,
5074	 => std_logic_vector(to_unsigned(101,8) ,
5075	 => std_logic_vector(to_unsigned(105,8) ,
5076	 => std_logic_vector(to_unsigned(107,8) ,
5077	 => std_logic_vector(to_unsigned(105,8) ,
5078	 => std_logic_vector(to_unsigned(104,8) ,
5079	 => std_logic_vector(to_unsigned(108,8) ,
5080	 => std_logic_vector(to_unsigned(112,8) ,
5081	 => std_logic_vector(to_unsigned(119,8) ,
5082	 => std_logic_vector(to_unsigned(121,8) ,
5083	 => std_logic_vector(to_unsigned(121,8) ,
5084	 => std_logic_vector(to_unsigned(124,8) ,
5085	 => std_logic_vector(to_unsigned(127,8) ,
5086	 => std_logic_vector(to_unsigned(127,8) ,
5087	 => std_logic_vector(to_unsigned(131,8) ,
5088	 => std_logic_vector(to_unsigned(136,8) ,
5089	 => std_logic_vector(to_unsigned(130,8) ,
5090	 => std_logic_vector(to_unsigned(124,8) ,
5091	 => std_logic_vector(to_unsigned(125,8) ,
5092	 => std_logic_vector(to_unsigned(130,8) ,
5093	 => std_logic_vector(to_unsigned(134,8) ,
5094	 => std_logic_vector(to_unsigned(134,8) ,
5095	 => std_logic_vector(to_unsigned(139,8) ,
5096	 => std_logic_vector(to_unsigned(142,8) ,
5097	 => std_logic_vector(to_unsigned(139,8) ,
5098	 => std_logic_vector(to_unsigned(141,8) ,
5099	 => std_logic_vector(to_unsigned(149,8) ,
5100	 => std_logic_vector(to_unsigned(154,8) ,
5101	 => std_logic_vector(to_unsigned(156,8) ,
5102	 => std_logic_vector(to_unsigned(154,8) ,
5103	 => std_logic_vector(to_unsigned(154,8) ,
5104	 => std_logic_vector(to_unsigned(157,8) ,
5105	 => std_logic_vector(to_unsigned(161,8) ,
5106	 => std_logic_vector(to_unsigned(157,8) ,
5107	 => std_logic_vector(to_unsigned(156,8) ,
5108	 => std_logic_vector(to_unsigned(161,8) ,
5109	 => std_logic_vector(to_unsigned(159,8) ,
5110	 => std_logic_vector(to_unsigned(157,8) ,
5111	 => std_logic_vector(to_unsigned(157,8) ,
5112	 => std_logic_vector(to_unsigned(159,8) ,
5113	 => std_logic_vector(to_unsigned(159,8) ,
5114	 => std_logic_vector(to_unsigned(156,8) ,
5115	 => std_logic_vector(to_unsigned(156,8) ,
5116	 => std_logic_vector(to_unsigned(161,8) ,
5117	 => std_logic_vector(to_unsigned(156,8) ,
5118	 => std_logic_vector(to_unsigned(156,8) ,
5119	 => std_logic_vector(to_unsigned(159,8) ,
5120	 => std_logic_vector(to_unsigned(157,8) ,
5121	 => std_logic_vector(to_unsigned(79,8) ,
5122	 => std_logic_vector(to_unsigned(76,8) ,
5123	 => std_logic_vector(to_unsigned(79,8) ,
5124	 => std_logic_vector(to_unsigned(71,8) ,
5125	 => std_logic_vector(to_unsigned(69,8) ,
5126	 => std_logic_vector(to_unsigned(80,8) ,
5127	 => std_logic_vector(to_unsigned(73,8) ,
5128	 => std_logic_vector(to_unsigned(71,8) ,
5129	 => std_logic_vector(to_unsigned(76,8) ,
5130	 => std_logic_vector(to_unsigned(67,8) ,
5131	 => std_logic_vector(to_unsigned(67,8) ,
5132	 => std_logic_vector(to_unsigned(71,8) ,
5133	 => std_logic_vector(to_unsigned(73,8) ,
5134	 => std_logic_vector(to_unsigned(76,8) ,
5135	 => std_logic_vector(to_unsigned(74,8) ,
5136	 => std_logic_vector(to_unsigned(67,8) ,
5137	 => std_logic_vector(to_unsigned(68,8) ,
5138	 => std_logic_vector(to_unsigned(71,8) ,
5139	 => std_logic_vector(to_unsigned(69,8) ,
5140	 => std_logic_vector(to_unsigned(67,8) ,
5141	 => std_logic_vector(to_unsigned(73,8) ,
5142	 => std_logic_vector(to_unsigned(79,8) ,
5143	 => std_logic_vector(to_unsigned(78,8) ,
5144	 => std_logic_vector(to_unsigned(76,8) ,
5145	 => std_logic_vector(to_unsigned(71,8) ,
5146	 => std_logic_vector(to_unsigned(76,8) ,
5147	 => std_logic_vector(to_unsigned(73,8) ,
5148	 => std_logic_vector(to_unsigned(64,8) ,
5149	 => std_logic_vector(to_unsigned(66,8) ,
5150	 => std_logic_vector(to_unsigned(69,8) ,
5151	 => std_logic_vector(to_unsigned(72,8) ,
5152	 => std_logic_vector(to_unsigned(76,8) ,
5153	 => std_logic_vector(to_unsigned(76,8) ,
5154	 => std_logic_vector(to_unsigned(68,8) ,
5155	 => std_logic_vector(to_unsigned(63,8) ,
5156	 => std_logic_vector(to_unsigned(74,8) ,
5157	 => std_logic_vector(to_unsigned(73,8) ,
5158	 => std_logic_vector(to_unsigned(78,8) ,
5159	 => std_logic_vector(to_unsigned(79,8) ,
5160	 => std_logic_vector(to_unsigned(80,8) ,
5161	 => std_logic_vector(to_unsigned(78,8) ,
5162	 => std_logic_vector(to_unsigned(81,8) ,
5163	 => std_logic_vector(to_unsigned(86,8) ,
5164	 => std_logic_vector(to_unsigned(82,8) ,
5165	 => std_logic_vector(to_unsigned(87,8) ,
5166	 => std_logic_vector(to_unsigned(91,8) ,
5167	 => std_logic_vector(to_unsigned(96,8) ,
5168	 => std_logic_vector(to_unsigned(97,8) ,
5169	 => std_logic_vector(to_unsigned(91,8) ,
5170	 => std_logic_vector(to_unsigned(92,8) ,
5171	 => std_logic_vector(to_unsigned(97,8) ,
5172	 => std_logic_vector(to_unsigned(97,8) ,
5173	 => std_logic_vector(to_unsigned(97,8) ,
5174	 => std_logic_vector(to_unsigned(105,8) ,
5175	 => std_logic_vector(to_unsigned(114,8) ,
5176	 => std_logic_vector(to_unsigned(107,8) ,
5177	 => std_logic_vector(to_unsigned(109,8) ,
5178	 => std_logic_vector(to_unsigned(105,8) ,
5179	 => std_logic_vector(to_unsigned(100,8) ,
5180	 => std_logic_vector(to_unsigned(108,8) ,
5181	 => std_logic_vector(to_unsigned(114,8) ,
5182	 => std_logic_vector(to_unsigned(108,8) ,
5183	 => std_logic_vector(to_unsigned(105,8) ,
5184	 => std_logic_vector(to_unsigned(108,8) ,
5185	 => std_logic_vector(to_unsigned(109,8) ,
5186	 => std_logic_vector(to_unsigned(111,8) ,
5187	 => std_logic_vector(to_unsigned(107,8) ,
5188	 => std_logic_vector(to_unsigned(111,8) ,
5189	 => std_logic_vector(to_unsigned(114,8) ,
5190	 => std_logic_vector(to_unsigned(115,8) ,
5191	 => std_logic_vector(to_unsigned(112,8) ,
5192	 => std_logic_vector(to_unsigned(107,8) ,
5193	 => std_logic_vector(to_unsigned(112,8) ,
5194	 => std_logic_vector(to_unsigned(115,8) ,
5195	 => std_logic_vector(to_unsigned(107,8) ,
5196	 => std_logic_vector(to_unsigned(105,8) ,
5197	 => std_logic_vector(to_unsigned(103,8) ,
5198	 => std_logic_vector(to_unsigned(99,8) ,
5199	 => std_logic_vector(to_unsigned(103,8) ,
5200	 => std_logic_vector(to_unsigned(104,8) ,
5201	 => std_logic_vector(to_unsigned(99,8) ,
5202	 => std_logic_vector(to_unsigned(90,8) ,
5203	 => std_logic_vector(to_unsigned(93,8) ,
5204	 => std_logic_vector(to_unsigned(100,8) ,
5205	 => std_logic_vector(to_unsigned(100,8) ,
5206	 => std_logic_vector(to_unsigned(92,8) ,
5207	 => std_logic_vector(to_unsigned(84,8) ,
5208	 => std_logic_vector(to_unsigned(85,8) ,
5209	 => std_logic_vector(to_unsigned(87,8) ,
5210	 => std_logic_vector(to_unsigned(88,8) ,
5211	 => std_logic_vector(to_unsigned(92,8) ,
5212	 => std_logic_vector(to_unsigned(84,8) ,
5213	 => std_logic_vector(to_unsigned(82,8) ,
5214	 => std_logic_vector(to_unsigned(84,8) ,
5215	 => std_logic_vector(to_unsigned(86,8) ,
5216	 => std_logic_vector(to_unsigned(79,8) ,
5217	 => std_logic_vector(to_unsigned(78,8) ,
5218	 => std_logic_vector(to_unsigned(77,8) ,
5219	 => std_logic_vector(to_unsigned(79,8) ,
5220	 => std_logic_vector(to_unsigned(80,8) ,
5221	 => std_logic_vector(to_unsigned(82,8) ,
5222	 => std_logic_vector(to_unsigned(77,8) ,
5223	 => std_logic_vector(to_unsigned(72,8) ,
5224	 => std_logic_vector(to_unsigned(74,8) ,
5225	 => std_logic_vector(to_unsigned(74,8) ,
5226	 => std_logic_vector(to_unsigned(76,8) ,
5227	 => std_logic_vector(to_unsigned(71,8) ,
5228	 => std_logic_vector(to_unsigned(71,8) ,
5229	 => std_logic_vector(to_unsigned(72,8) ,
5230	 => std_logic_vector(to_unsigned(72,8) ,
5231	 => std_logic_vector(to_unsigned(71,8) ,
5232	 => std_logic_vector(to_unsigned(74,8) ,
5233	 => std_logic_vector(to_unsigned(77,8) ,
5234	 => std_logic_vector(to_unsigned(80,8) ,
5235	 => std_logic_vector(to_unsigned(85,8) ,
5236	 => std_logic_vector(to_unsigned(86,8) ,
5237	 => std_logic_vector(to_unsigned(90,8) ,
5238	 => std_logic_vector(to_unsigned(84,8) ,
5239	 => std_logic_vector(to_unsigned(84,8) ,
5240	 => std_logic_vector(to_unsigned(82,8) ,
5241	 => std_logic_vector(to_unsigned(87,8) ,
5242	 => std_logic_vector(to_unsigned(87,8) ,
5243	 => std_logic_vector(to_unsigned(84,8) ,
5244	 => std_logic_vector(to_unsigned(92,8) ,
5245	 => std_logic_vector(to_unsigned(90,8) ,
5246	 => std_logic_vector(to_unsigned(91,8) ,
5247	 => std_logic_vector(to_unsigned(90,8) ,
5248	 => std_logic_vector(to_unsigned(93,8) ,
5249	 => std_logic_vector(to_unsigned(97,8) ,
5250	 => std_logic_vector(to_unsigned(95,8) ,
5251	 => std_logic_vector(to_unsigned(90,8) ,
5252	 => std_logic_vector(to_unsigned(91,8) ,
5253	 => std_logic_vector(to_unsigned(91,8) ,
5254	 => std_logic_vector(to_unsigned(92,8) ,
5255	 => std_logic_vector(to_unsigned(90,8) ,
5256	 => std_logic_vector(to_unsigned(90,8) ,
5257	 => std_logic_vector(to_unsigned(92,8) ,
5258	 => std_logic_vector(to_unsigned(90,8) ,
5259	 => std_logic_vector(to_unsigned(87,8) ,
5260	 => std_logic_vector(to_unsigned(87,8) ,
5261	 => std_logic_vector(to_unsigned(93,8) ,
5262	 => std_logic_vector(to_unsigned(95,8) ,
5263	 => std_logic_vector(to_unsigned(100,8) ,
5264	 => std_logic_vector(to_unsigned(104,8) ,
5265	 => std_logic_vector(to_unsigned(97,8) ,
5266	 => std_logic_vector(to_unsigned(96,8) ,
5267	 => std_logic_vector(to_unsigned(97,8) ,
5268	 => std_logic_vector(to_unsigned(93,8) ,
5269	 => std_logic_vector(to_unsigned(93,8) ,
5270	 => std_logic_vector(to_unsigned(95,8) ,
5271	 => std_logic_vector(to_unsigned(91,8) ,
5272	 => std_logic_vector(to_unsigned(93,8) ,
5273	 => std_logic_vector(to_unsigned(92,8) ,
5274	 => std_logic_vector(to_unsigned(92,8) ,
5275	 => std_logic_vector(to_unsigned(95,8) ,
5276	 => std_logic_vector(to_unsigned(92,8) ,
5277	 => std_logic_vector(to_unsigned(91,8) ,
5278	 => std_logic_vector(to_unsigned(92,8) ,
5279	 => std_logic_vector(to_unsigned(88,8) ,
5280	 => std_logic_vector(to_unsigned(86,8) ,
5281	 => std_logic_vector(to_unsigned(85,8) ,
5282	 => std_logic_vector(to_unsigned(80,8) ,
5283	 => std_logic_vector(to_unsigned(79,8) ,
5284	 => std_logic_vector(to_unsigned(82,8) ,
5285	 => std_logic_vector(to_unsigned(81,8) ,
5286	 => std_logic_vector(to_unsigned(79,8) ,
5287	 => std_logic_vector(to_unsigned(79,8) ,
5288	 => std_logic_vector(to_unsigned(81,8) ,
5289	 => std_logic_vector(to_unsigned(82,8) ,
5290	 => std_logic_vector(to_unsigned(79,8) ,
5291	 => std_logic_vector(to_unsigned(82,8) ,
5292	 => std_logic_vector(to_unsigned(80,8) ,
5293	 => std_logic_vector(to_unsigned(79,8) ,
5294	 => std_logic_vector(to_unsigned(80,8) ,
5295	 => std_logic_vector(to_unsigned(73,8) ,
5296	 => std_logic_vector(to_unsigned(74,8) ,
5297	 => std_logic_vector(to_unsigned(74,8) ,
5298	 => std_logic_vector(to_unsigned(76,8) ,
5299	 => std_logic_vector(to_unsigned(73,8) ,
5300	 => std_logic_vector(to_unsigned(72,8) ,
5301	 => std_logic_vector(to_unsigned(76,8) ,
5302	 => std_logic_vector(to_unsigned(78,8) ,
5303	 => std_logic_vector(to_unsigned(71,8) ,
5304	 => std_logic_vector(to_unsigned(71,8) ,
5305	 => std_logic_vector(to_unsigned(70,8) ,
5306	 => std_logic_vector(to_unsigned(70,8) ,
5307	 => std_logic_vector(to_unsigned(78,8) ,
5308	 => std_logic_vector(to_unsigned(77,8) ,
5309	 => std_logic_vector(to_unsigned(79,8) ,
5310	 => std_logic_vector(to_unsigned(77,8) ,
5311	 => std_logic_vector(to_unsigned(79,8) ,
5312	 => std_logic_vector(to_unsigned(81,8) ,
5313	 => std_logic_vector(to_unsigned(77,8) ,
5314	 => std_logic_vector(to_unsigned(70,8) ,
5315	 => std_logic_vector(to_unsigned(82,8) ,
5316	 => std_logic_vector(to_unsigned(82,8) ,
5317	 => std_logic_vector(to_unsigned(77,8) ,
5318	 => std_logic_vector(to_unsigned(73,8) ,
5319	 => std_logic_vector(to_unsigned(77,8) ,
5320	 => std_logic_vector(to_unsigned(81,8) ,
5321	 => std_logic_vector(to_unsigned(82,8) ,
5322	 => std_logic_vector(to_unsigned(79,8) ,
5323	 => std_logic_vector(to_unsigned(80,8) ,
5324	 => std_logic_vector(to_unsigned(84,8) ,
5325	 => std_logic_vector(to_unsigned(82,8) ,
5326	 => std_logic_vector(to_unsigned(81,8) ,
5327	 => std_logic_vector(to_unsigned(82,8) ,
5328	 => std_logic_vector(to_unsigned(86,8) ,
5329	 => std_logic_vector(to_unsigned(82,8) ,
5330	 => std_logic_vector(to_unsigned(78,8) ,
5331	 => std_logic_vector(to_unsigned(85,8) ,
5332	 => std_logic_vector(to_unsigned(88,8) ,
5333	 => std_logic_vector(to_unsigned(84,8) ,
5334	 => std_logic_vector(to_unsigned(87,8) ,
5335	 => std_logic_vector(to_unsigned(88,8) ,
5336	 => std_logic_vector(to_unsigned(87,8) ,
5337	 => std_logic_vector(to_unsigned(87,8) ,
5338	 => std_logic_vector(to_unsigned(85,8) ,
5339	 => std_logic_vector(to_unsigned(84,8) ,
5340	 => std_logic_vector(to_unsigned(81,8) ,
5341	 => std_logic_vector(to_unsigned(86,8) ,
5342	 => std_logic_vector(to_unsigned(91,8) ,
5343	 => std_logic_vector(to_unsigned(88,8) ,
5344	 => std_logic_vector(to_unsigned(85,8) ,
5345	 => std_logic_vector(to_unsigned(88,8) ,
5346	 => std_logic_vector(to_unsigned(87,8) ,
5347	 => std_logic_vector(to_unsigned(87,8) ,
5348	 => std_logic_vector(to_unsigned(74,8) ,
5349	 => std_logic_vector(to_unsigned(73,8) ,
5350	 => std_logic_vector(to_unsigned(69,8) ,
5351	 => std_logic_vector(to_unsigned(64,8) ,
5352	 => std_logic_vector(to_unsigned(71,8) ,
5353	 => std_logic_vector(to_unsigned(82,8) ,
5354	 => std_logic_vector(to_unsigned(84,8) ,
5355	 => std_logic_vector(to_unsigned(86,8) ,
5356	 => std_logic_vector(to_unsigned(74,8) ,
5357	 => std_logic_vector(to_unsigned(77,8) ,
5358	 => std_logic_vector(to_unsigned(74,8) ,
5359	 => std_logic_vector(to_unsigned(13,8) ,
5360	 => std_logic_vector(to_unsigned(0,8) ,
5361	 => std_logic_vector(to_unsigned(0,8) ,
5362	 => std_logic_vector(to_unsigned(8,8) ,
5363	 => std_logic_vector(to_unsigned(78,8) ,
5364	 => std_logic_vector(to_unsigned(84,8) ,
5365	 => std_logic_vector(to_unsigned(81,8) ,
5366	 => std_logic_vector(to_unsigned(91,8) ,
5367	 => std_logic_vector(to_unsigned(96,8) ,
5368	 => std_logic_vector(to_unsigned(93,8) ,
5369	 => std_logic_vector(to_unsigned(87,8) ,
5370	 => std_logic_vector(to_unsigned(93,8) ,
5371	 => std_logic_vector(to_unsigned(103,8) ,
5372	 => std_logic_vector(to_unsigned(133,8) ,
5373	 => std_logic_vector(to_unsigned(116,8) ,
5374	 => std_logic_vector(to_unsigned(92,8) ,
5375	 => std_logic_vector(to_unsigned(101,8) ,
5376	 => std_logic_vector(to_unsigned(95,8) ,
5377	 => std_logic_vector(to_unsigned(86,8) ,
5378	 => std_logic_vector(to_unsigned(86,8) ,
5379	 => std_logic_vector(to_unsigned(80,8) ,
5380	 => std_logic_vector(to_unsigned(80,8) ,
5381	 => std_logic_vector(to_unsigned(88,8) ,
5382	 => std_logic_vector(to_unsigned(92,8) ,
5383	 => std_logic_vector(to_unsigned(91,8) ,
5384	 => std_logic_vector(to_unsigned(85,8) ,
5385	 => std_logic_vector(to_unsigned(91,8) ,
5386	 => std_logic_vector(to_unsigned(88,8) ,
5387	 => std_logic_vector(to_unsigned(85,8) ,
5388	 => std_logic_vector(to_unsigned(78,8) ,
5389	 => std_logic_vector(to_unsigned(77,8) ,
5390	 => std_logic_vector(to_unsigned(85,8) ,
5391	 => std_logic_vector(to_unsigned(87,8) ,
5392	 => std_logic_vector(to_unsigned(93,8) ,
5393	 => std_logic_vector(to_unsigned(93,8) ,
5394	 => std_logic_vector(to_unsigned(92,8) ,
5395	 => std_logic_vector(to_unsigned(103,8) ,
5396	 => std_logic_vector(to_unsigned(105,8) ,
5397	 => std_logic_vector(to_unsigned(105,8) ,
5398	 => std_logic_vector(to_unsigned(103,8) ,
5399	 => std_logic_vector(to_unsigned(108,8) ,
5400	 => std_logic_vector(to_unsigned(111,8) ,
5401	 => std_logic_vector(to_unsigned(114,8) ,
5402	 => std_logic_vector(to_unsigned(121,8) ,
5403	 => std_logic_vector(to_unsigned(124,8) ,
5404	 => std_logic_vector(to_unsigned(125,8) ,
5405	 => std_logic_vector(to_unsigned(130,8) ,
5406	 => std_logic_vector(to_unsigned(130,8) ,
5407	 => std_logic_vector(to_unsigned(133,8) ,
5408	 => std_logic_vector(to_unsigned(133,8) ,
5409	 => std_logic_vector(to_unsigned(133,8) ,
5410	 => std_logic_vector(to_unsigned(131,8) ,
5411	 => std_logic_vector(to_unsigned(138,8) ,
5412	 => std_logic_vector(to_unsigned(141,8) ,
5413	 => std_logic_vector(to_unsigned(141,8) ,
5414	 => std_logic_vector(to_unsigned(141,8) ,
5415	 => std_logic_vector(to_unsigned(149,8) ,
5416	 => std_logic_vector(to_unsigned(147,8) ,
5417	 => std_logic_vector(to_unsigned(141,8) ,
5418	 => std_logic_vector(to_unsigned(144,8) ,
5419	 => std_logic_vector(to_unsigned(149,8) ,
5420	 => std_logic_vector(to_unsigned(149,8) ,
5421	 => std_logic_vector(to_unsigned(154,8) ,
5422	 => std_logic_vector(to_unsigned(154,8) ,
5423	 => std_logic_vector(to_unsigned(154,8) ,
5424	 => std_logic_vector(to_unsigned(154,8) ,
5425	 => std_logic_vector(to_unsigned(156,8) ,
5426	 => std_logic_vector(to_unsigned(157,8) ,
5427	 => std_logic_vector(to_unsigned(157,8) ,
5428	 => std_logic_vector(to_unsigned(161,8) ,
5429	 => std_logic_vector(to_unsigned(157,8) ,
5430	 => std_logic_vector(to_unsigned(157,8) ,
5431	 => std_logic_vector(to_unsigned(156,8) ,
5432	 => std_logic_vector(to_unsigned(157,8) ,
5433	 => std_logic_vector(to_unsigned(159,8) ,
5434	 => std_logic_vector(to_unsigned(157,8) ,
5435	 => std_logic_vector(to_unsigned(159,8) ,
5436	 => std_logic_vector(to_unsigned(159,8) ,
5437	 => std_logic_vector(to_unsigned(159,8) ,
5438	 => std_logic_vector(to_unsigned(157,8) ,
5439	 => std_logic_vector(to_unsigned(157,8) ,
5440	 => std_logic_vector(to_unsigned(159,8) ,
5441	 => std_logic_vector(to_unsigned(77,8) ,
5442	 => std_logic_vector(to_unsigned(72,8) ,
5443	 => std_logic_vector(to_unsigned(70,8) ,
5444	 => std_logic_vector(to_unsigned(74,8) ,
5445	 => std_logic_vector(to_unsigned(65,8) ,
5446	 => std_logic_vector(to_unsigned(73,8) ,
5447	 => std_logic_vector(to_unsigned(73,8) ,
5448	 => std_logic_vector(to_unsigned(73,8) ,
5449	 => std_logic_vector(to_unsigned(78,8) ,
5450	 => std_logic_vector(to_unsigned(67,8) ,
5451	 => std_logic_vector(to_unsigned(66,8) ,
5452	 => std_logic_vector(to_unsigned(68,8) ,
5453	 => std_logic_vector(to_unsigned(66,8) ,
5454	 => std_logic_vector(to_unsigned(70,8) ,
5455	 => std_logic_vector(to_unsigned(76,8) ,
5456	 => std_logic_vector(to_unsigned(71,8) ,
5457	 => std_logic_vector(to_unsigned(70,8) ,
5458	 => std_logic_vector(to_unsigned(69,8) ,
5459	 => std_logic_vector(to_unsigned(71,8) ,
5460	 => std_logic_vector(to_unsigned(68,8) ,
5461	 => std_logic_vector(to_unsigned(72,8) ,
5462	 => std_logic_vector(to_unsigned(72,8) ,
5463	 => std_logic_vector(to_unsigned(71,8) ,
5464	 => std_logic_vector(to_unsigned(77,8) ,
5465	 => std_logic_vector(to_unsigned(77,8) ,
5466	 => std_logic_vector(to_unsigned(74,8) ,
5467	 => std_logic_vector(to_unsigned(67,8) ,
5468	 => std_logic_vector(to_unsigned(66,8) ,
5469	 => std_logic_vector(to_unsigned(59,8) ,
5470	 => std_logic_vector(to_unsigned(66,8) ,
5471	 => std_logic_vector(to_unsigned(70,8) ,
5472	 => std_logic_vector(to_unsigned(69,8) ,
5473	 => std_logic_vector(to_unsigned(73,8) ,
5474	 => std_logic_vector(to_unsigned(72,8) ,
5475	 => std_logic_vector(to_unsigned(68,8) ,
5476	 => std_logic_vector(to_unsigned(71,8) ,
5477	 => std_logic_vector(to_unsigned(68,8) ,
5478	 => std_logic_vector(to_unsigned(70,8) ,
5479	 => std_logic_vector(to_unsigned(73,8) ,
5480	 => std_logic_vector(to_unsigned(73,8) ,
5481	 => std_logic_vector(to_unsigned(74,8) ,
5482	 => std_logic_vector(to_unsigned(79,8) ,
5483	 => std_logic_vector(to_unsigned(87,8) ,
5484	 => std_logic_vector(to_unsigned(85,8) ,
5485	 => std_logic_vector(to_unsigned(85,8) ,
5486	 => std_logic_vector(to_unsigned(91,8) ,
5487	 => std_logic_vector(to_unsigned(88,8) ,
5488	 => std_logic_vector(to_unsigned(91,8) ,
5489	 => std_logic_vector(to_unsigned(92,8) ,
5490	 => std_logic_vector(to_unsigned(96,8) ,
5491	 => std_logic_vector(to_unsigned(97,8) ,
5492	 => std_logic_vector(to_unsigned(97,8) ,
5493	 => std_logic_vector(to_unsigned(103,8) ,
5494	 => std_logic_vector(to_unsigned(104,8) ,
5495	 => std_logic_vector(to_unsigned(109,8) ,
5496	 => std_logic_vector(to_unsigned(105,8) ,
5497	 => std_logic_vector(to_unsigned(105,8) ,
5498	 => std_logic_vector(to_unsigned(109,8) ,
5499	 => std_logic_vector(to_unsigned(103,8) ,
5500	 => std_logic_vector(to_unsigned(107,8) ,
5501	 => std_logic_vector(to_unsigned(112,8) ,
5502	 => std_logic_vector(to_unsigned(99,8) ,
5503	 => std_logic_vector(to_unsigned(96,8) ,
5504	 => std_logic_vector(to_unsigned(103,8) ,
5505	 => std_logic_vector(to_unsigned(107,8) ,
5506	 => std_logic_vector(to_unsigned(112,8) ,
5507	 => std_logic_vector(to_unsigned(103,8) ,
5508	 => std_logic_vector(to_unsigned(107,8) ,
5509	 => std_logic_vector(to_unsigned(116,8) ,
5510	 => std_logic_vector(to_unsigned(118,8) ,
5511	 => std_logic_vector(to_unsigned(115,8) ,
5512	 => std_logic_vector(to_unsigned(114,8) ,
5513	 => std_logic_vector(to_unsigned(114,8) ,
5514	 => std_logic_vector(to_unsigned(108,8) ,
5515	 => std_logic_vector(to_unsigned(107,8) ,
5516	 => std_logic_vector(to_unsigned(111,8) ,
5517	 => std_logic_vector(to_unsigned(107,8) ,
5518	 => std_logic_vector(to_unsigned(99,8) ,
5519	 => std_logic_vector(to_unsigned(104,8) ,
5520	 => std_logic_vector(to_unsigned(112,8) ,
5521	 => std_logic_vector(to_unsigned(103,8) ,
5522	 => std_logic_vector(to_unsigned(92,8) ,
5523	 => std_logic_vector(to_unsigned(92,8) ,
5524	 => std_logic_vector(to_unsigned(99,8) ,
5525	 => std_logic_vector(to_unsigned(105,8) ,
5526	 => std_logic_vector(to_unsigned(99,8) ,
5527	 => std_logic_vector(to_unsigned(86,8) ,
5528	 => std_logic_vector(to_unsigned(84,8) ,
5529	 => std_logic_vector(to_unsigned(86,8) ,
5530	 => std_logic_vector(to_unsigned(85,8) ,
5531	 => std_logic_vector(to_unsigned(88,8) ,
5532	 => std_logic_vector(to_unsigned(82,8) ,
5533	 => std_logic_vector(to_unsigned(81,8) ,
5534	 => std_logic_vector(to_unsigned(79,8) ,
5535	 => std_logic_vector(to_unsigned(77,8) ,
5536	 => std_logic_vector(to_unsigned(77,8) ,
5537	 => std_logic_vector(to_unsigned(80,8) ,
5538	 => std_logic_vector(to_unsigned(77,8) ,
5539	 => std_logic_vector(to_unsigned(74,8) ,
5540	 => std_logic_vector(to_unsigned(78,8) ,
5541	 => std_logic_vector(to_unsigned(73,8) ,
5542	 => std_logic_vector(to_unsigned(73,8) ,
5543	 => std_logic_vector(to_unsigned(72,8) ,
5544	 => std_logic_vector(to_unsigned(72,8) ,
5545	 => std_logic_vector(to_unsigned(74,8) ,
5546	 => std_logic_vector(to_unsigned(76,8) ,
5547	 => std_logic_vector(to_unsigned(70,8) ,
5548	 => std_logic_vector(to_unsigned(72,8) ,
5549	 => std_logic_vector(to_unsigned(72,8) ,
5550	 => std_logic_vector(to_unsigned(72,8) ,
5551	 => std_logic_vector(to_unsigned(74,8) ,
5552	 => std_logic_vector(to_unsigned(76,8) ,
5553	 => std_logic_vector(to_unsigned(74,8) ,
5554	 => std_logic_vector(to_unsigned(78,8) ,
5555	 => std_logic_vector(to_unsigned(76,8) ,
5556	 => std_logic_vector(to_unsigned(78,8) ,
5557	 => std_logic_vector(to_unsigned(85,8) ,
5558	 => std_logic_vector(to_unsigned(82,8) ,
5559	 => std_logic_vector(to_unsigned(84,8) ,
5560	 => std_logic_vector(to_unsigned(85,8) ,
5561	 => std_logic_vector(to_unsigned(85,8) ,
5562	 => std_logic_vector(to_unsigned(85,8) ,
5563	 => std_logic_vector(to_unsigned(82,8) ,
5564	 => std_logic_vector(to_unsigned(82,8) ,
5565	 => std_logic_vector(to_unsigned(90,8) ,
5566	 => std_logic_vector(to_unsigned(92,8) ,
5567	 => std_logic_vector(to_unsigned(90,8) ,
5568	 => std_logic_vector(to_unsigned(91,8) ,
5569	 => std_logic_vector(to_unsigned(95,8) ,
5570	 => std_logic_vector(to_unsigned(93,8) ,
5571	 => std_logic_vector(to_unsigned(91,8) ,
5572	 => std_logic_vector(to_unsigned(92,8) ,
5573	 => std_logic_vector(to_unsigned(92,8) ,
5574	 => std_logic_vector(to_unsigned(90,8) ,
5575	 => std_logic_vector(to_unsigned(87,8) ,
5576	 => std_logic_vector(to_unsigned(90,8) ,
5577	 => std_logic_vector(to_unsigned(88,8) ,
5578	 => std_logic_vector(to_unsigned(86,8) ,
5579	 => std_logic_vector(to_unsigned(86,8) ,
5580	 => std_logic_vector(to_unsigned(81,8) ,
5581	 => std_logic_vector(to_unsigned(91,8) ,
5582	 => std_logic_vector(to_unsigned(93,8) ,
5583	 => std_logic_vector(to_unsigned(97,8) ,
5584	 => std_logic_vector(to_unsigned(97,8) ,
5585	 => std_logic_vector(to_unsigned(91,8) ,
5586	 => std_logic_vector(to_unsigned(93,8) ,
5587	 => std_logic_vector(to_unsigned(92,8) ,
5588	 => std_logic_vector(to_unsigned(95,8) ,
5589	 => std_logic_vector(to_unsigned(90,8) ,
5590	 => std_logic_vector(to_unsigned(91,8) ,
5591	 => std_logic_vector(to_unsigned(91,8) ,
5592	 => std_logic_vector(to_unsigned(90,8) ,
5593	 => std_logic_vector(to_unsigned(87,8) ,
5594	 => std_logic_vector(to_unsigned(92,8) ,
5595	 => std_logic_vector(to_unsigned(95,8) ,
5596	 => std_logic_vector(to_unsigned(90,8) ,
5597	 => std_logic_vector(to_unsigned(90,8) ,
5598	 => std_logic_vector(to_unsigned(88,8) ,
5599	 => std_logic_vector(to_unsigned(87,8) ,
5600	 => std_logic_vector(to_unsigned(91,8) ,
5601	 => std_logic_vector(to_unsigned(85,8) ,
5602	 => std_logic_vector(to_unsigned(86,8) ,
5603	 => std_logic_vector(to_unsigned(82,8) ,
5604	 => std_logic_vector(to_unsigned(81,8) ,
5605	 => std_logic_vector(to_unsigned(84,8) ,
5606	 => std_logic_vector(to_unsigned(84,8) ,
5607	 => std_logic_vector(to_unsigned(82,8) ,
5608	 => std_logic_vector(to_unsigned(82,8) ,
5609	 => std_logic_vector(to_unsigned(80,8) ,
5610	 => std_logic_vector(to_unsigned(78,8) ,
5611	 => std_logic_vector(to_unsigned(79,8) ,
5612	 => std_logic_vector(to_unsigned(78,8) ,
5613	 => std_logic_vector(to_unsigned(74,8) ,
5614	 => std_logic_vector(to_unsigned(79,8) ,
5615	 => std_logic_vector(to_unsigned(77,8) ,
5616	 => std_logic_vector(to_unsigned(71,8) ,
5617	 => std_logic_vector(to_unsigned(73,8) ,
5618	 => std_logic_vector(to_unsigned(71,8) ,
5619	 => std_logic_vector(to_unsigned(71,8) ,
5620	 => std_logic_vector(to_unsigned(71,8) ,
5621	 => std_logic_vector(to_unsigned(76,8) ,
5622	 => std_logic_vector(to_unsigned(73,8) ,
5623	 => std_logic_vector(to_unsigned(71,8) ,
5624	 => std_logic_vector(to_unsigned(72,8) ,
5625	 => std_logic_vector(to_unsigned(72,8) ,
5626	 => std_logic_vector(to_unsigned(72,8) ,
5627	 => std_logic_vector(to_unsigned(77,8) ,
5628	 => std_logic_vector(to_unsigned(77,8) ,
5629	 => std_logic_vector(to_unsigned(79,8) ,
5630	 => std_logic_vector(to_unsigned(79,8) ,
5631	 => std_logic_vector(to_unsigned(79,8) ,
5632	 => std_logic_vector(to_unsigned(79,8) ,
5633	 => std_logic_vector(to_unsigned(66,8) ,
5634	 => std_logic_vector(to_unsigned(58,8) ,
5635	 => std_logic_vector(to_unsigned(77,8) ,
5636	 => std_logic_vector(to_unsigned(78,8) ,
5637	 => std_logic_vector(to_unsigned(78,8) ,
5638	 => std_logic_vector(to_unsigned(77,8) ,
5639	 => std_logic_vector(to_unsigned(79,8) ,
5640	 => std_logic_vector(to_unsigned(82,8) ,
5641	 => std_logic_vector(to_unsigned(81,8) ,
5642	 => std_logic_vector(to_unsigned(72,8) ,
5643	 => std_logic_vector(to_unsigned(74,8) ,
5644	 => std_logic_vector(to_unsigned(82,8) ,
5645	 => std_logic_vector(to_unsigned(81,8) ,
5646	 => std_logic_vector(to_unsigned(81,8) ,
5647	 => std_logic_vector(to_unsigned(86,8) ,
5648	 => std_logic_vector(to_unsigned(88,8) ,
5649	 => std_logic_vector(to_unsigned(79,8) ,
5650	 => std_logic_vector(to_unsigned(80,8) ,
5651	 => std_logic_vector(to_unsigned(88,8) ,
5652	 => std_logic_vector(to_unsigned(85,8) ,
5653	 => std_logic_vector(to_unsigned(84,8) ,
5654	 => std_logic_vector(to_unsigned(87,8) ,
5655	 => std_logic_vector(to_unsigned(87,8) ,
5656	 => std_logic_vector(to_unsigned(95,8) ,
5657	 => std_logic_vector(to_unsigned(86,8) ,
5658	 => std_logic_vector(to_unsigned(82,8) ,
5659	 => std_logic_vector(to_unsigned(86,8) ,
5660	 => std_logic_vector(to_unsigned(85,8) ,
5661	 => std_logic_vector(to_unsigned(86,8) ,
5662	 => std_logic_vector(to_unsigned(85,8) ,
5663	 => std_logic_vector(to_unsigned(79,8) ,
5664	 => std_logic_vector(to_unsigned(85,8) ,
5665	 => std_logic_vector(to_unsigned(80,8) ,
5666	 => std_logic_vector(to_unsigned(73,8) ,
5667	 => std_logic_vector(to_unsigned(73,8) ,
5668	 => std_logic_vector(to_unsigned(64,8) ,
5669	 => std_logic_vector(to_unsigned(53,8) ,
5670	 => std_logic_vector(to_unsigned(57,8) ,
5671	 => std_logic_vector(to_unsigned(61,8) ,
5672	 => std_logic_vector(to_unsigned(65,8) ,
5673	 => std_logic_vector(to_unsigned(77,8) ,
5674	 => std_logic_vector(to_unsigned(82,8) ,
5675	 => std_logic_vector(to_unsigned(80,8) ,
5676	 => std_logic_vector(to_unsigned(68,8) ,
5677	 => std_logic_vector(to_unsigned(61,8) ,
5678	 => std_logic_vector(to_unsigned(63,8) ,
5679	 => std_logic_vector(to_unsigned(22,8) ,
5680	 => std_logic_vector(to_unsigned(0,8) ,
5681	 => std_logic_vector(to_unsigned(0,8) ,
5682	 => std_logic_vector(to_unsigned(3,8) ,
5683	 => std_logic_vector(to_unsigned(63,8) ,
5684	 => std_logic_vector(to_unsigned(86,8) ,
5685	 => std_logic_vector(to_unsigned(77,8) ,
5686	 => std_logic_vector(to_unsigned(80,8) ,
5687	 => std_logic_vector(to_unsigned(82,8) ,
5688	 => std_logic_vector(to_unsigned(81,8) ,
5689	 => std_logic_vector(to_unsigned(82,8) ,
5690	 => std_logic_vector(to_unsigned(90,8) ,
5691	 => std_logic_vector(to_unsigned(99,8) ,
5692	 => std_logic_vector(to_unsigned(114,8) ,
5693	 => std_logic_vector(to_unsigned(95,8) ,
5694	 => std_logic_vector(to_unsigned(87,8) ,
5695	 => std_logic_vector(to_unsigned(101,8) ,
5696	 => std_logic_vector(to_unsigned(95,8) ,
5697	 => std_logic_vector(to_unsigned(90,8) ,
5698	 => std_logic_vector(to_unsigned(86,8) ,
5699	 => std_logic_vector(to_unsigned(85,8) ,
5700	 => std_logic_vector(to_unsigned(85,8) ,
5701	 => std_logic_vector(to_unsigned(81,8) ,
5702	 => std_logic_vector(to_unsigned(82,8) ,
5703	 => std_logic_vector(to_unsigned(82,8) ,
5704	 => std_logic_vector(to_unsigned(85,8) ,
5705	 => std_logic_vector(to_unsigned(88,8) ,
5706	 => std_logic_vector(to_unsigned(84,8) ,
5707	 => std_logic_vector(to_unsigned(76,8) ,
5708	 => std_logic_vector(to_unsigned(72,8) ,
5709	 => std_logic_vector(to_unsigned(77,8) ,
5710	 => std_logic_vector(to_unsigned(79,8) ,
5711	 => std_logic_vector(to_unsigned(86,8) ,
5712	 => std_logic_vector(to_unsigned(93,8) ,
5713	 => std_logic_vector(to_unsigned(92,8) ,
5714	 => std_logic_vector(to_unsigned(95,8) ,
5715	 => std_logic_vector(to_unsigned(99,8) ,
5716	 => std_logic_vector(to_unsigned(104,8) ,
5717	 => std_logic_vector(to_unsigned(112,8) ,
5718	 => std_logic_vector(to_unsigned(108,8) ,
5719	 => std_logic_vector(to_unsigned(109,8) ,
5720	 => std_logic_vector(to_unsigned(118,8) ,
5721	 => std_logic_vector(to_unsigned(124,8) ,
5722	 => std_logic_vector(to_unsigned(127,8) ,
5723	 => std_logic_vector(to_unsigned(125,8) ,
5724	 => std_logic_vector(to_unsigned(127,8) ,
5725	 => std_logic_vector(to_unsigned(128,8) ,
5726	 => std_logic_vector(to_unsigned(127,8) ,
5727	 => std_logic_vector(to_unsigned(127,8) ,
5728	 => std_logic_vector(to_unsigned(127,8) ,
5729	 => std_logic_vector(to_unsigned(131,8) ,
5730	 => std_logic_vector(to_unsigned(130,8) ,
5731	 => std_logic_vector(to_unsigned(127,8) ,
5732	 => std_logic_vector(to_unsigned(133,8) ,
5733	 => std_logic_vector(to_unsigned(141,8) ,
5734	 => std_logic_vector(to_unsigned(141,8) ,
5735	 => std_logic_vector(to_unsigned(146,8) ,
5736	 => std_logic_vector(to_unsigned(142,8) ,
5737	 => std_logic_vector(to_unsigned(142,8) ,
5738	 => std_logic_vector(to_unsigned(149,8) ,
5739	 => std_logic_vector(to_unsigned(149,8) ,
5740	 => std_logic_vector(to_unsigned(146,8) ,
5741	 => std_logic_vector(to_unsigned(152,8) ,
5742	 => std_logic_vector(to_unsigned(154,8) ,
5743	 => std_logic_vector(to_unsigned(154,8) ,
5744	 => std_logic_vector(to_unsigned(152,8) ,
5745	 => std_logic_vector(to_unsigned(154,8) ,
5746	 => std_logic_vector(to_unsigned(159,8) ,
5747	 => std_logic_vector(to_unsigned(159,8) ,
5748	 => std_logic_vector(to_unsigned(157,8) ,
5749	 => std_logic_vector(to_unsigned(157,8) ,
5750	 => std_logic_vector(to_unsigned(157,8) ,
5751	 => std_logic_vector(to_unsigned(156,8) ,
5752	 => std_logic_vector(to_unsigned(152,8) ,
5753	 => std_logic_vector(to_unsigned(152,8) ,
5754	 => std_logic_vector(to_unsigned(161,8) ,
5755	 => std_logic_vector(to_unsigned(159,8) ,
5756	 => std_logic_vector(to_unsigned(157,8) ,
5757	 => std_logic_vector(to_unsigned(161,8) ,
5758	 => std_logic_vector(to_unsigned(157,8) ,
5759	 => std_logic_vector(to_unsigned(159,8) ,
5760	 => std_logic_vector(to_unsigned(163,8) ,
5761	 => std_logic_vector(to_unsigned(80,8) ,
5762	 => std_logic_vector(to_unsigned(86,8) ,
5763	 => std_logic_vector(to_unsigned(73,8) ,
5764	 => std_logic_vector(to_unsigned(68,8) ,
5765	 => std_logic_vector(to_unsigned(73,8) ,
5766	 => std_logic_vector(to_unsigned(74,8) ,
5767	 => std_logic_vector(to_unsigned(68,8) ,
5768	 => std_logic_vector(to_unsigned(70,8) ,
5769	 => std_logic_vector(to_unsigned(71,8) ,
5770	 => std_logic_vector(to_unsigned(68,8) ,
5771	 => std_logic_vector(to_unsigned(68,8) ,
5772	 => std_logic_vector(to_unsigned(69,8) ,
5773	 => std_logic_vector(to_unsigned(67,8) ,
5774	 => std_logic_vector(to_unsigned(72,8) ,
5775	 => std_logic_vector(to_unsigned(79,8) ,
5776	 => std_logic_vector(to_unsigned(72,8) ,
5777	 => std_logic_vector(to_unsigned(77,8) ,
5778	 => std_logic_vector(to_unsigned(70,8) ,
5779	 => std_logic_vector(to_unsigned(64,8) ,
5780	 => std_logic_vector(to_unsigned(70,8) ,
5781	 => std_logic_vector(to_unsigned(69,8) ,
5782	 => std_logic_vector(to_unsigned(65,8) ,
5783	 => std_logic_vector(to_unsigned(71,8) ,
5784	 => std_logic_vector(to_unsigned(77,8) ,
5785	 => std_logic_vector(to_unsigned(80,8) ,
5786	 => std_logic_vector(to_unsigned(73,8) ,
5787	 => std_logic_vector(to_unsigned(72,8) ,
5788	 => std_logic_vector(to_unsigned(71,8) ,
5789	 => std_logic_vector(to_unsigned(64,8) ,
5790	 => std_logic_vector(to_unsigned(65,8) ,
5791	 => std_logic_vector(to_unsigned(68,8) ,
5792	 => std_logic_vector(to_unsigned(70,8) ,
5793	 => std_logic_vector(to_unsigned(73,8) ,
5794	 => std_logic_vector(to_unsigned(74,8) ,
5795	 => std_logic_vector(to_unsigned(71,8) ,
5796	 => std_logic_vector(to_unsigned(70,8) ,
5797	 => std_logic_vector(to_unsigned(72,8) ,
5798	 => std_logic_vector(to_unsigned(76,8) ,
5799	 => std_logic_vector(to_unsigned(79,8) ,
5800	 => std_logic_vector(to_unsigned(76,8) ,
5801	 => std_logic_vector(to_unsigned(76,8) ,
5802	 => std_logic_vector(to_unsigned(80,8) ,
5803	 => std_logic_vector(to_unsigned(84,8) ,
5804	 => std_logic_vector(to_unsigned(85,8) ,
5805	 => std_logic_vector(to_unsigned(92,8) ,
5806	 => std_logic_vector(to_unsigned(95,8) ,
5807	 => std_logic_vector(to_unsigned(88,8) ,
5808	 => std_logic_vector(to_unsigned(90,8) ,
5809	 => std_logic_vector(to_unsigned(97,8) ,
5810	 => std_logic_vector(to_unsigned(100,8) ,
5811	 => std_logic_vector(to_unsigned(95,8) ,
5812	 => std_logic_vector(to_unsigned(99,8) ,
5813	 => std_logic_vector(to_unsigned(104,8) ,
5814	 => std_logic_vector(to_unsigned(108,8) ,
5815	 => std_logic_vector(to_unsigned(114,8) ,
5816	 => std_logic_vector(to_unsigned(114,8) ,
5817	 => std_logic_vector(to_unsigned(108,8) ,
5818	 => std_logic_vector(to_unsigned(114,8) ,
5819	 => std_logic_vector(to_unsigned(107,8) ,
5820	 => std_logic_vector(to_unsigned(103,8) ,
5821	 => std_logic_vector(to_unsigned(108,8) ,
5822	 => std_logic_vector(to_unsigned(100,8) ,
5823	 => std_logic_vector(to_unsigned(95,8) ,
5824	 => std_logic_vector(to_unsigned(97,8) ,
5825	 => std_logic_vector(to_unsigned(103,8) ,
5826	 => std_logic_vector(to_unsigned(109,8) ,
5827	 => std_logic_vector(to_unsigned(105,8) ,
5828	 => std_logic_vector(to_unsigned(111,8) ,
5829	 => std_logic_vector(to_unsigned(116,8) ,
5830	 => std_logic_vector(to_unsigned(111,8) ,
5831	 => std_logic_vector(to_unsigned(108,8) ,
5832	 => std_logic_vector(to_unsigned(109,8) ,
5833	 => std_logic_vector(to_unsigned(107,8) ,
5834	 => std_logic_vector(to_unsigned(105,8) ,
5835	 => std_logic_vector(to_unsigned(109,8) ,
5836	 => std_logic_vector(to_unsigned(115,8) ,
5837	 => std_logic_vector(to_unsigned(107,8) ,
5838	 => std_logic_vector(to_unsigned(101,8) ,
5839	 => std_logic_vector(to_unsigned(104,8) ,
5840	 => std_logic_vector(to_unsigned(104,8) ,
5841	 => std_logic_vector(to_unsigned(97,8) ,
5842	 => std_logic_vector(to_unsigned(97,8) ,
5843	 => std_logic_vector(to_unsigned(99,8) ,
5844	 => std_logic_vector(to_unsigned(96,8) ,
5845	 => std_logic_vector(to_unsigned(100,8) ,
5846	 => std_logic_vector(to_unsigned(100,8) ,
5847	 => std_logic_vector(to_unsigned(92,8) ,
5848	 => std_logic_vector(to_unsigned(90,8) ,
5849	 => std_logic_vector(to_unsigned(86,8) ,
5850	 => std_logic_vector(to_unsigned(79,8) ,
5851	 => std_logic_vector(to_unsigned(81,8) ,
5852	 => std_logic_vector(to_unsigned(84,8) ,
5853	 => std_logic_vector(to_unsigned(84,8) ,
5854	 => std_logic_vector(to_unsigned(81,8) ,
5855	 => std_logic_vector(to_unsigned(80,8) ,
5856	 => std_logic_vector(to_unsigned(81,8) ,
5857	 => std_logic_vector(to_unsigned(78,8) ,
5858	 => std_logic_vector(to_unsigned(77,8) ,
5859	 => std_logic_vector(to_unsigned(77,8) ,
5860	 => std_logic_vector(to_unsigned(78,8) ,
5861	 => std_logic_vector(to_unsigned(76,8) ,
5862	 => std_logic_vector(to_unsigned(73,8) ,
5863	 => std_logic_vector(to_unsigned(72,8) ,
5864	 => std_logic_vector(to_unsigned(78,8) ,
5865	 => std_logic_vector(to_unsigned(76,8) ,
5866	 => std_logic_vector(to_unsigned(72,8) ,
5867	 => std_logic_vector(to_unsigned(72,8) ,
5868	 => std_logic_vector(to_unsigned(73,8) ,
5869	 => std_logic_vector(to_unsigned(69,8) ,
5870	 => std_logic_vector(to_unsigned(67,8) ,
5871	 => std_logic_vector(to_unsigned(71,8) ,
5872	 => std_logic_vector(to_unsigned(74,8) ,
5873	 => std_logic_vector(to_unsigned(74,8) ,
5874	 => std_logic_vector(to_unsigned(77,8) ,
5875	 => std_logic_vector(to_unsigned(80,8) ,
5876	 => std_logic_vector(to_unsigned(79,8) ,
5877	 => std_logic_vector(to_unsigned(80,8) ,
5878	 => std_logic_vector(to_unsigned(84,8) ,
5879	 => std_logic_vector(to_unsigned(87,8) ,
5880	 => std_logic_vector(to_unsigned(90,8) ,
5881	 => std_logic_vector(to_unsigned(86,8) ,
5882	 => std_logic_vector(to_unsigned(88,8) ,
5883	 => std_logic_vector(to_unsigned(92,8) ,
5884	 => std_logic_vector(to_unsigned(93,8) ,
5885	 => std_logic_vector(to_unsigned(95,8) ,
5886	 => std_logic_vector(to_unsigned(92,8) ,
5887	 => std_logic_vector(to_unsigned(88,8) ,
5888	 => std_logic_vector(to_unsigned(87,8) ,
5889	 => std_logic_vector(to_unsigned(90,8) ,
5890	 => std_logic_vector(to_unsigned(90,8) ,
5891	 => std_logic_vector(to_unsigned(88,8) ,
5892	 => std_logic_vector(to_unsigned(88,8) ,
5893	 => std_logic_vector(to_unsigned(87,8) ,
5894	 => std_logic_vector(to_unsigned(86,8) ,
5895	 => std_logic_vector(to_unsigned(86,8) ,
5896	 => std_logic_vector(to_unsigned(88,8) ,
5897	 => std_logic_vector(to_unsigned(88,8) ,
5898	 => std_logic_vector(to_unsigned(85,8) ,
5899	 => std_logic_vector(to_unsigned(90,8) ,
5900	 => std_logic_vector(to_unsigned(91,8) ,
5901	 => std_logic_vector(to_unsigned(91,8) ,
5902	 => std_logic_vector(to_unsigned(90,8) ,
5903	 => std_logic_vector(to_unsigned(93,8) ,
5904	 => std_logic_vector(to_unsigned(97,8) ,
5905	 => std_logic_vector(to_unsigned(95,8) ,
5906	 => std_logic_vector(to_unsigned(95,8) ,
5907	 => std_logic_vector(to_unsigned(95,8) ,
5908	 => std_logic_vector(to_unsigned(92,8) ,
5909	 => std_logic_vector(to_unsigned(87,8) ,
5910	 => std_logic_vector(to_unsigned(88,8) ,
5911	 => std_logic_vector(to_unsigned(82,8) ,
5912	 => std_logic_vector(to_unsigned(88,8) ,
5913	 => std_logic_vector(to_unsigned(92,8) ,
5914	 => std_logic_vector(to_unsigned(88,8) ,
5915	 => std_logic_vector(to_unsigned(87,8) ,
5916	 => std_logic_vector(to_unsigned(90,8) ,
5917	 => std_logic_vector(to_unsigned(91,8) ,
5918	 => std_logic_vector(to_unsigned(92,8) ,
5919	 => std_logic_vector(to_unsigned(88,8) ,
5920	 => std_logic_vector(to_unsigned(91,8) ,
5921	 => std_logic_vector(to_unsigned(88,8) ,
5922	 => std_logic_vector(to_unsigned(86,8) ,
5923	 => std_logic_vector(to_unsigned(81,8) ,
5924	 => std_logic_vector(to_unsigned(80,8) ,
5925	 => std_logic_vector(to_unsigned(84,8) ,
5926	 => std_logic_vector(to_unsigned(84,8) ,
5927	 => std_logic_vector(to_unsigned(80,8) ,
5928	 => std_logic_vector(to_unsigned(79,8) ,
5929	 => std_logic_vector(to_unsigned(84,8) ,
5930	 => std_logic_vector(to_unsigned(79,8) ,
5931	 => std_logic_vector(to_unsigned(71,8) ,
5932	 => std_logic_vector(to_unsigned(74,8) ,
5933	 => std_logic_vector(to_unsigned(80,8) ,
5934	 => std_logic_vector(to_unsigned(79,8) ,
5935	 => std_logic_vector(to_unsigned(78,8) ,
5936	 => std_logic_vector(to_unsigned(77,8) ,
5937	 => std_logic_vector(to_unsigned(79,8) ,
5938	 => std_logic_vector(to_unsigned(72,8) ,
5939	 => std_logic_vector(to_unsigned(76,8) ,
5940	 => std_logic_vector(to_unsigned(77,8) ,
5941	 => std_logic_vector(to_unsigned(70,8) ,
5942	 => std_logic_vector(to_unsigned(74,8) ,
5943	 => std_logic_vector(to_unsigned(74,8) ,
5944	 => std_logic_vector(to_unsigned(74,8) ,
5945	 => std_logic_vector(to_unsigned(72,8) ,
5946	 => std_logic_vector(to_unsigned(78,8) ,
5947	 => std_logic_vector(to_unsigned(79,8) ,
5948	 => std_logic_vector(to_unsigned(77,8) ,
5949	 => std_logic_vector(to_unsigned(78,8) ,
5950	 => std_logic_vector(to_unsigned(80,8) ,
5951	 => std_logic_vector(to_unsigned(79,8) ,
5952	 => std_logic_vector(to_unsigned(77,8) ,
5953	 => std_logic_vector(to_unsigned(62,8) ,
5954	 => std_logic_vector(to_unsigned(57,8) ,
5955	 => std_logic_vector(to_unsigned(72,8) ,
5956	 => std_logic_vector(to_unsigned(79,8) ,
5957	 => std_logic_vector(to_unsigned(81,8) ,
5958	 => std_logic_vector(to_unsigned(77,8) ,
5959	 => std_logic_vector(to_unsigned(81,8) ,
5960	 => std_logic_vector(to_unsigned(86,8) ,
5961	 => std_logic_vector(to_unsigned(86,8) ,
5962	 => std_logic_vector(to_unsigned(87,8) ,
5963	 => std_logic_vector(to_unsigned(81,8) ,
5964	 => std_logic_vector(to_unsigned(80,8) ,
5965	 => std_logic_vector(to_unsigned(85,8) ,
5966	 => std_logic_vector(to_unsigned(90,8) ,
5967	 => std_logic_vector(to_unsigned(93,8) ,
5968	 => std_logic_vector(to_unsigned(90,8) ,
5969	 => std_logic_vector(to_unsigned(85,8) ,
5970	 => std_logic_vector(to_unsigned(86,8) ,
5971	 => std_logic_vector(to_unsigned(82,8) ,
5972	 => std_logic_vector(to_unsigned(86,8) ,
5973	 => std_logic_vector(to_unsigned(87,8) ,
5974	 => std_logic_vector(to_unsigned(81,8) ,
5975	 => std_logic_vector(to_unsigned(76,8) ,
5976	 => std_logic_vector(to_unsigned(84,8) ,
5977	 => std_logic_vector(to_unsigned(78,8) ,
5978	 => std_logic_vector(to_unsigned(72,8) ,
5979	 => std_logic_vector(to_unsigned(78,8) ,
5980	 => std_logic_vector(to_unsigned(74,8) ,
5981	 => std_logic_vector(to_unsigned(74,8) ,
5982	 => std_logic_vector(to_unsigned(73,8) ,
5983	 => std_logic_vector(to_unsigned(66,8) ,
5984	 => std_logic_vector(to_unsigned(68,8) ,
5985	 => std_logic_vector(to_unsigned(63,8) ,
5986	 => std_logic_vector(to_unsigned(60,8) ,
5987	 => std_logic_vector(to_unsigned(67,8) ,
5988	 => std_logic_vector(to_unsigned(64,8) ,
5989	 => std_logic_vector(to_unsigned(50,8) ,
5990	 => std_logic_vector(to_unsigned(52,8) ,
5991	 => std_logic_vector(to_unsigned(61,8) ,
5992	 => std_logic_vector(to_unsigned(64,8) ,
5993	 => std_logic_vector(to_unsigned(69,8) ,
5994	 => std_logic_vector(to_unsigned(68,8) ,
5995	 => std_logic_vector(to_unsigned(68,8) ,
5996	 => std_logic_vector(to_unsigned(70,8) ,
5997	 => std_logic_vector(to_unsigned(65,8) ,
5998	 => std_logic_vector(to_unsigned(59,8) ,
5999	 => std_logic_vector(to_unsigned(45,8) ,
6000	 => std_logic_vector(to_unsigned(2,8) ,
6001	 => std_logic_vector(to_unsigned(0,8) ,
6002	 => std_logic_vector(to_unsigned(1,8) ,
6003	 => std_logic_vector(to_unsigned(39,8) ,
6004	 => std_logic_vector(to_unsigned(90,8) ,
6005	 => std_logic_vector(to_unsigned(72,8) ,
6006	 => std_logic_vector(to_unsigned(76,8) ,
6007	 => std_logic_vector(to_unsigned(80,8) ,
6008	 => std_logic_vector(to_unsigned(81,8) ,
6009	 => std_logic_vector(to_unsigned(81,8) ,
6010	 => std_logic_vector(to_unsigned(87,8) ,
6011	 => std_logic_vector(to_unsigned(92,8) ,
6012	 => std_logic_vector(to_unsigned(92,8) ,
6013	 => std_logic_vector(to_unsigned(88,8) ,
6014	 => std_logic_vector(to_unsigned(92,8) ,
6015	 => std_logic_vector(to_unsigned(91,8) ,
6016	 => std_logic_vector(to_unsigned(84,8) ,
6017	 => std_logic_vector(to_unsigned(81,8) ,
6018	 => std_logic_vector(to_unsigned(78,8) ,
6019	 => std_logic_vector(to_unsigned(80,8) ,
6020	 => std_logic_vector(to_unsigned(79,8) ,
6021	 => std_logic_vector(to_unsigned(69,8) ,
6022	 => std_logic_vector(to_unsigned(67,8) ,
6023	 => std_logic_vector(to_unsigned(76,8) ,
6024	 => std_logic_vector(to_unsigned(81,8) ,
6025	 => std_logic_vector(to_unsigned(82,8) ,
6026	 => std_logic_vector(to_unsigned(79,8) ,
6027	 => std_logic_vector(to_unsigned(67,8) ,
6028	 => std_logic_vector(to_unsigned(69,8) ,
6029	 => std_logic_vector(to_unsigned(79,8) ,
6030	 => std_logic_vector(to_unsigned(82,8) ,
6031	 => std_logic_vector(to_unsigned(96,8) ,
6032	 => std_logic_vector(to_unsigned(95,8) ,
6033	 => std_logic_vector(to_unsigned(91,8) ,
6034	 => std_logic_vector(to_unsigned(103,8) ,
6035	 => std_logic_vector(to_unsigned(107,8) ,
6036	 => std_logic_vector(to_unsigned(104,8) ,
6037	 => std_logic_vector(to_unsigned(105,8) ,
6038	 => std_logic_vector(to_unsigned(105,8) ,
6039	 => std_logic_vector(to_unsigned(115,8) ,
6040	 => std_logic_vector(to_unsigned(118,8) ,
6041	 => std_logic_vector(to_unsigned(118,8) ,
6042	 => std_logic_vector(to_unsigned(122,8) ,
6043	 => std_logic_vector(to_unsigned(128,8) ,
6044	 => std_logic_vector(to_unsigned(119,8) ,
6045	 => std_logic_vector(to_unsigned(124,8) ,
6046	 => std_logic_vector(to_unsigned(130,8) ,
6047	 => std_logic_vector(to_unsigned(127,8) ,
6048	 => std_logic_vector(to_unsigned(122,8) ,
6049	 => std_logic_vector(to_unsigned(125,8) ,
6050	 => std_logic_vector(to_unsigned(127,8) ,
6051	 => std_logic_vector(to_unsigned(127,8) ,
6052	 => std_logic_vector(to_unsigned(131,8) ,
6053	 => std_logic_vector(to_unsigned(133,8) ,
6054	 => std_logic_vector(to_unsigned(130,8) ,
6055	 => std_logic_vector(to_unsigned(136,8) ,
6056	 => std_logic_vector(to_unsigned(136,8) ,
6057	 => std_logic_vector(to_unsigned(136,8) ,
6058	 => std_logic_vector(to_unsigned(144,8) ,
6059	 => std_logic_vector(to_unsigned(147,8) ,
6060	 => std_logic_vector(to_unsigned(144,8) ,
6061	 => std_logic_vector(to_unsigned(146,8) ,
6062	 => std_logic_vector(to_unsigned(149,8) ,
6063	 => std_logic_vector(to_unsigned(152,8) ,
6064	 => std_logic_vector(to_unsigned(154,8) ,
6065	 => std_logic_vector(to_unsigned(156,8) ,
6066	 => std_logic_vector(to_unsigned(157,8) ,
6067	 => std_logic_vector(to_unsigned(156,8) ,
6068	 => std_logic_vector(to_unsigned(156,8) ,
6069	 => std_logic_vector(to_unsigned(159,8) ,
6070	 => std_logic_vector(to_unsigned(156,8) ,
6071	 => std_logic_vector(to_unsigned(154,8) ,
6072	 => std_logic_vector(to_unsigned(147,8) ,
6073	 => std_logic_vector(to_unsigned(149,8) ,
6074	 => std_logic_vector(to_unsigned(154,8) ,
6075	 => std_logic_vector(to_unsigned(156,8) ,
6076	 => std_logic_vector(to_unsigned(157,8) ,
6077	 => std_logic_vector(to_unsigned(159,8) ,
6078	 => std_logic_vector(to_unsigned(156,8) ,
6079	 => std_logic_vector(to_unsigned(159,8) ,
6080	 => std_logic_vector(to_unsigned(163,8) ,
6081	 => std_logic_vector(to_unsigned(85,8) ,
6082	 => std_logic_vector(to_unsigned(82,8) ,
6083	 => std_logic_vector(to_unsigned(78,8) ,
6084	 => std_logic_vector(to_unsigned(76,8) ,
6085	 => std_logic_vector(to_unsigned(79,8) ,
6086	 => std_logic_vector(to_unsigned(74,8) ,
6087	 => std_logic_vector(to_unsigned(73,8) ,
6088	 => std_logic_vector(to_unsigned(74,8) ,
6089	 => std_logic_vector(to_unsigned(72,8) ,
6090	 => std_logic_vector(to_unsigned(71,8) ,
6091	 => std_logic_vector(to_unsigned(69,8) ,
6092	 => std_logic_vector(to_unsigned(70,8) ,
6093	 => std_logic_vector(to_unsigned(74,8) ,
6094	 => std_logic_vector(to_unsigned(77,8) ,
6095	 => std_logic_vector(to_unsigned(74,8) ,
6096	 => std_logic_vector(to_unsigned(72,8) ,
6097	 => std_logic_vector(to_unsigned(76,8) ,
6098	 => std_logic_vector(to_unsigned(76,8) ,
6099	 => std_logic_vector(to_unsigned(70,8) ,
6100	 => std_logic_vector(to_unsigned(71,8) ,
6101	 => std_logic_vector(to_unsigned(73,8) ,
6102	 => std_logic_vector(to_unsigned(69,8) ,
6103	 => std_logic_vector(to_unsigned(70,8) ,
6104	 => std_logic_vector(to_unsigned(72,8) ,
6105	 => std_logic_vector(to_unsigned(73,8) ,
6106	 => std_logic_vector(to_unsigned(70,8) ,
6107	 => std_logic_vector(to_unsigned(71,8) ,
6108	 => std_logic_vector(to_unsigned(71,8) ,
6109	 => std_logic_vector(to_unsigned(69,8) ,
6110	 => std_logic_vector(to_unsigned(66,8) ,
6111	 => std_logic_vector(to_unsigned(69,8) ,
6112	 => std_logic_vector(to_unsigned(74,8) ,
6113	 => std_logic_vector(to_unsigned(73,8) ,
6114	 => std_logic_vector(to_unsigned(76,8) ,
6115	 => std_logic_vector(to_unsigned(76,8) ,
6116	 => std_logic_vector(to_unsigned(71,8) ,
6117	 => std_logic_vector(to_unsigned(78,8) ,
6118	 => std_logic_vector(to_unsigned(81,8) ,
6119	 => std_logic_vector(to_unsigned(84,8) ,
6120	 => std_logic_vector(to_unsigned(85,8) ,
6121	 => std_logic_vector(to_unsigned(82,8) ,
6122	 => std_logic_vector(to_unsigned(81,8) ,
6123	 => std_logic_vector(to_unsigned(88,8) ,
6124	 => std_logic_vector(to_unsigned(91,8) ,
6125	 => std_logic_vector(to_unsigned(92,8) ,
6126	 => std_logic_vector(to_unsigned(91,8) ,
6127	 => std_logic_vector(to_unsigned(92,8) ,
6128	 => std_logic_vector(to_unsigned(95,8) ,
6129	 => std_logic_vector(to_unsigned(99,8) ,
6130	 => std_logic_vector(to_unsigned(96,8) ,
6131	 => std_logic_vector(to_unsigned(90,8) ,
6132	 => std_logic_vector(to_unsigned(100,8) ,
6133	 => std_logic_vector(to_unsigned(103,8) ,
6134	 => std_logic_vector(to_unsigned(107,8) ,
6135	 => std_logic_vector(to_unsigned(114,8) ,
6136	 => std_logic_vector(to_unsigned(115,8) ,
6137	 => std_logic_vector(to_unsigned(115,8) ,
6138	 => std_logic_vector(to_unsigned(121,8) ,
6139	 => std_logic_vector(to_unsigned(111,8) ,
6140	 => std_logic_vector(to_unsigned(104,8) ,
6141	 => std_logic_vector(to_unsigned(107,8) ,
6142	 => std_logic_vector(to_unsigned(104,8) ,
6143	 => std_logic_vector(to_unsigned(103,8) ,
6144	 => std_logic_vector(to_unsigned(104,8) ,
6145	 => std_logic_vector(to_unsigned(107,8) ,
6146	 => std_logic_vector(to_unsigned(108,8) ,
6147	 => std_logic_vector(to_unsigned(107,8) ,
6148	 => std_logic_vector(to_unsigned(109,8) ,
6149	 => std_logic_vector(to_unsigned(109,8) ,
6150	 => std_logic_vector(to_unsigned(107,8) ,
6151	 => std_logic_vector(to_unsigned(107,8) ,
6152	 => std_logic_vector(to_unsigned(107,8) ,
6153	 => std_logic_vector(to_unsigned(109,8) ,
6154	 => std_logic_vector(to_unsigned(109,8) ,
6155	 => std_logic_vector(to_unsigned(104,8) ,
6156	 => std_logic_vector(to_unsigned(105,8) ,
6157	 => std_logic_vector(to_unsigned(105,8) ,
6158	 => std_logic_vector(to_unsigned(105,8) ,
6159	 => std_logic_vector(to_unsigned(105,8) ,
6160	 => std_logic_vector(to_unsigned(99,8) ,
6161	 => std_logic_vector(to_unsigned(96,8) ,
6162	 => std_logic_vector(to_unsigned(100,8) ,
6163	 => std_logic_vector(to_unsigned(100,8) ,
6164	 => std_logic_vector(to_unsigned(96,8) ,
6165	 => std_logic_vector(to_unsigned(96,8) ,
6166	 => std_logic_vector(to_unsigned(97,8) ,
6167	 => std_logic_vector(to_unsigned(99,8) ,
6168	 => std_logic_vector(to_unsigned(97,8) ,
6169	 => std_logic_vector(to_unsigned(92,8) ,
6170	 => std_logic_vector(to_unsigned(87,8) ,
6171	 => std_logic_vector(to_unsigned(85,8) ,
6172	 => std_logic_vector(to_unsigned(87,8) ,
6173	 => std_logic_vector(to_unsigned(86,8) ,
6174	 => std_logic_vector(to_unsigned(85,8) ,
6175	 => std_logic_vector(to_unsigned(84,8) ,
6176	 => std_logic_vector(to_unsigned(81,8) ,
6177	 => std_logic_vector(to_unsigned(77,8) ,
6178	 => std_logic_vector(to_unsigned(82,8) ,
6179	 => std_logic_vector(to_unsigned(81,8) ,
6180	 => std_logic_vector(to_unsigned(80,8) ,
6181	 => std_logic_vector(to_unsigned(84,8) ,
6182	 => std_logic_vector(to_unsigned(77,8) ,
6183	 => std_logic_vector(to_unsigned(79,8) ,
6184	 => std_logic_vector(to_unsigned(78,8) ,
6185	 => std_logic_vector(to_unsigned(72,8) ,
6186	 => std_logic_vector(to_unsigned(70,8) ,
6187	 => std_logic_vector(to_unsigned(71,8) ,
6188	 => std_logic_vector(to_unsigned(70,8) ,
6189	 => std_logic_vector(to_unsigned(70,8) ,
6190	 => std_logic_vector(to_unsigned(73,8) ,
6191	 => std_logic_vector(to_unsigned(72,8) ,
6192	 => std_logic_vector(to_unsigned(71,8) ,
6193	 => std_logic_vector(to_unsigned(77,8) ,
6194	 => std_logic_vector(to_unsigned(79,8) ,
6195	 => std_logic_vector(to_unsigned(80,8) ,
6196	 => std_logic_vector(to_unsigned(81,8) ,
6197	 => std_logic_vector(to_unsigned(82,8) ,
6198	 => std_logic_vector(to_unsigned(84,8) ,
6199	 => std_logic_vector(to_unsigned(88,8) ,
6200	 => std_logic_vector(to_unsigned(90,8) ,
6201	 => std_logic_vector(to_unsigned(93,8) ,
6202	 => std_logic_vector(to_unsigned(92,8) ,
6203	 => std_logic_vector(to_unsigned(90,8) ,
6204	 => std_logic_vector(to_unsigned(101,8) ,
6205	 => std_logic_vector(to_unsigned(99,8) ,
6206	 => std_logic_vector(to_unsigned(90,8) ,
6207	 => std_logic_vector(to_unsigned(90,8) ,
6208	 => std_logic_vector(to_unsigned(88,8) ,
6209	 => std_logic_vector(to_unsigned(91,8) ,
6210	 => std_logic_vector(to_unsigned(92,8) ,
6211	 => std_logic_vector(to_unsigned(91,8) ,
6212	 => std_logic_vector(to_unsigned(87,8) ,
6213	 => std_logic_vector(to_unsigned(88,8) ,
6214	 => std_logic_vector(to_unsigned(88,8) ,
6215	 => std_logic_vector(to_unsigned(86,8) ,
6216	 => std_logic_vector(to_unsigned(86,8) ,
6217	 => std_logic_vector(to_unsigned(87,8) ,
6218	 => std_logic_vector(to_unsigned(82,8) ,
6219	 => std_logic_vector(to_unsigned(90,8) ,
6220	 => std_logic_vector(to_unsigned(93,8) ,
6221	 => std_logic_vector(to_unsigned(92,8) ,
6222	 => std_logic_vector(to_unsigned(88,8) ,
6223	 => std_logic_vector(to_unsigned(90,8) ,
6224	 => std_logic_vector(to_unsigned(93,8) ,
6225	 => std_logic_vector(to_unsigned(93,8) ,
6226	 => std_logic_vector(to_unsigned(96,8) ,
6227	 => std_logic_vector(to_unsigned(96,8) ,
6228	 => std_logic_vector(to_unsigned(88,8) ,
6229	 => std_logic_vector(to_unsigned(87,8) ,
6230	 => std_logic_vector(to_unsigned(90,8) ,
6231	 => std_logic_vector(to_unsigned(86,8) ,
6232	 => std_logic_vector(to_unsigned(90,8) ,
6233	 => std_logic_vector(to_unsigned(93,8) ,
6234	 => std_logic_vector(to_unsigned(90,8) ,
6235	 => std_logic_vector(to_unsigned(85,8) ,
6236	 => std_logic_vector(to_unsigned(85,8) ,
6237	 => std_logic_vector(to_unsigned(87,8) ,
6238	 => std_logic_vector(to_unsigned(90,8) ,
6239	 => std_logic_vector(to_unsigned(88,8) ,
6240	 => std_logic_vector(to_unsigned(85,8) ,
6241	 => std_logic_vector(to_unsigned(90,8) ,
6242	 => std_logic_vector(to_unsigned(90,8) ,
6243	 => std_logic_vector(to_unsigned(86,8) ,
6244	 => std_logic_vector(to_unsigned(85,8) ,
6245	 => std_logic_vector(to_unsigned(81,8) ,
6246	 => std_logic_vector(to_unsigned(78,8) ,
6247	 => std_logic_vector(to_unsigned(78,8) ,
6248	 => std_logic_vector(to_unsigned(80,8) ,
6249	 => std_logic_vector(to_unsigned(81,8) ,
6250	 => std_logic_vector(to_unsigned(79,8) ,
6251	 => std_logic_vector(to_unsigned(79,8) ,
6252	 => std_logic_vector(to_unsigned(79,8) ,
6253	 => std_logic_vector(to_unsigned(82,8) ,
6254	 => std_logic_vector(to_unsigned(81,8) ,
6255	 => std_logic_vector(to_unsigned(80,8) ,
6256	 => std_logic_vector(to_unsigned(79,8) ,
6257	 => std_logic_vector(to_unsigned(79,8) ,
6258	 => std_logic_vector(to_unsigned(76,8) ,
6259	 => std_logic_vector(to_unsigned(77,8) ,
6260	 => std_logic_vector(to_unsigned(79,8) ,
6261	 => std_logic_vector(to_unsigned(76,8) ,
6262	 => std_logic_vector(to_unsigned(81,8) ,
6263	 => std_logic_vector(to_unsigned(79,8) ,
6264	 => std_logic_vector(to_unsigned(73,8) ,
6265	 => std_logic_vector(to_unsigned(76,8) ,
6266	 => std_logic_vector(to_unsigned(78,8) ,
6267	 => std_logic_vector(to_unsigned(80,8) ,
6268	 => std_logic_vector(to_unsigned(77,8) ,
6269	 => std_logic_vector(to_unsigned(85,8) ,
6270	 => std_logic_vector(to_unsigned(84,8) ,
6271	 => std_logic_vector(to_unsigned(80,8) ,
6272	 => std_logic_vector(to_unsigned(85,8) ,
6273	 => std_logic_vector(to_unsigned(68,8) ,
6274	 => std_logic_vector(to_unsigned(68,8) ,
6275	 => std_logic_vector(to_unsigned(77,8) ,
6276	 => std_logic_vector(to_unsigned(86,8) ,
6277	 => std_logic_vector(to_unsigned(85,8) ,
6278	 => std_logic_vector(to_unsigned(79,8) ,
6279	 => std_logic_vector(to_unsigned(81,8) ,
6280	 => std_logic_vector(to_unsigned(86,8) ,
6281	 => std_logic_vector(to_unsigned(78,8) ,
6282	 => std_logic_vector(to_unsigned(78,8) ,
6283	 => std_logic_vector(to_unsigned(82,8) ,
6284	 => std_logic_vector(to_unsigned(81,8) ,
6285	 => std_logic_vector(to_unsigned(77,8) ,
6286	 => std_logic_vector(to_unsigned(74,8) ,
6287	 => std_logic_vector(to_unsigned(88,8) ,
6288	 => std_logic_vector(to_unsigned(91,8) ,
6289	 => std_logic_vector(to_unsigned(74,8) ,
6290	 => std_logic_vector(to_unsigned(74,8) ,
6291	 => std_logic_vector(to_unsigned(72,8) ,
6292	 => std_logic_vector(to_unsigned(77,8) ,
6293	 => std_logic_vector(to_unsigned(74,8) ,
6294	 => std_logic_vector(to_unsigned(74,8) ,
6295	 => std_logic_vector(to_unsigned(71,8) ,
6296	 => std_logic_vector(to_unsigned(71,8) ,
6297	 => std_logic_vector(to_unsigned(76,8) ,
6298	 => std_logic_vector(to_unsigned(73,8) ,
6299	 => std_logic_vector(to_unsigned(71,8) ,
6300	 => std_logic_vector(to_unsigned(66,8) ,
6301	 => std_logic_vector(to_unsigned(64,8) ,
6302	 => std_logic_vector(to_unsigned(61,8) ,
6303	 => std_logic_vector(to_unsigned(60,8) ,
6304	 => std_logic_vector(to_unsigned(64,8) ,
6305	 => std_logic_vector(to_unsigned(61,8) ,
6306	 => std_logic_vector(to_unsigned(62,8) ,
6307	 => std_logic_vector(to_unsigned(68,8) ,
6308	 => std_logic_vector(to_unsigned(63,8) ,
6309	 => std_logic_vector(to_unsigned(60,8) ,
6310	 => std_logic_vector(to_unsigned(59,8) ,
6311	 => std_logic_vector(to_unsigned(60,8) ,
6312	 => std_logic_vector(to_unsigned(59,8) ,
6313	 => std_logic_vector(to_unsigned(66,8) ,
6314	 => std_logic_vector(to_unsigned(64,8) ,
6315	 => std_logic_vector(to_unsigned(60,8) ,
6316	 => std_logic_vector(to_unsigned(59,8) ,
6317	 => std_logic_vector(to_unsigned(59,8) ,
6318	 => std_logic_vector(to_unsigned(58,8) ,
6319	 => std_logic_vector(to_unsigned(54,8) ,
6320	 => std_logic_vector(to_unsigned(4,8) ,
6321	 => std_logic_vector(to_unsigned(0,8) ,
6322	 => std_logic_vector(to_unsigned(0,8) ,
6323	 => std_logic_vector(to_unsigned(18,8) ,
6324	 => std_logic_vector(to_unsigned(81,8) ,
6325	 => std_logic_vector(to_unsigned(71,8) ,
6326	 => std_logic_vector(to_unsigned(80,8) ,
6327	 => std_logic_vector(to_unsigned(81,8) ,
6328	 => std_logic_vector(to_unsigned(74,8) ,
6329	 => std_logic_vector(to_unsigned(72,8) ,
6330	 => std_logic_vector(to_unsigned(76,8) ,
6331	 => std_logic_vector(to_unsigned(88,8) ,
6332	 => std_logic_vector(to_unsigned(90,8) ,
6333	 => std_logic_vector(to_unsigned(87,8) ,
6334	 => std_logic_vector(to_unsigned(91,8) ,
6335	 => std_logic_vector(to_unsigned(90,8) ,
6336	 => std_logic_vector(to_unsigned(87,8) ,
6337	 => std_logic_vector(to_unsigned(80,8) ,
6338	 => std_logic_vector(to_unsigned(77,8) ,
6339	 => std_logic_vector(to_unsigned(74,8) ,
6340	 => std_logic_vector(to_unsigned(76,8) ,
6341	 => std_logic_vector(to_unsigned(73,8) ,
6342	 => std_logic_vector(to_unsigned(71,8) ,
6343	 => std_logic_vector(to_unsigned(79,8) ,
6344	 => std_logic_vector(to_unsigned(78,8) ,
6345	 => std_logic_vector(to_unsigned(80,8) ,
6346	 => std_logic_vector(to_unsigned(81,8) ,
6347	 => std_logic_vector(to_unsigned(73,8) ,
6348	 => std_logic_vector(to_unsigned(73,8) ,
6349	 => std_logic_vector(to_unsigned(81,8) ,
6350	 => std_logic_vector(to_unsigned(97,8) ,
6351	 => std_logic_vector(to_unsigned(97,8) ,
6352	 => std_logic_vector(to_unsigned(88,8) ,
6353	 => std_logic_vector(to_unsigned(95,8) ,
6354	 => std_logic_vector(to_unsigned(97,8) ,
6355	 => std_logic_vector(to_unsigned(99,8) ,
6356	 => std_logic_vector(to_unsigned(97,8) ,
6357	 => std_logic_vector(to_unsigned(96,8) ,
6358	 => std_logic_vector(to_unsigned(97,8) ,
6359	 => std_logic_vector(to_unsigned(105,8) ,
6360	 => std_logic_vector(to_unsigned(109,8) ,
6361	 => std_logic_vector(to_unsigned(116,8) ,
6362	 => std_logic_vector(to_unsigned(115,8) ,
6363	 => std_logic_vector(to_unsigned(118,8) ,
6364	 => std_logic_vector(to_unsigned(122,8) ,
6365	 => std_logic_vector(to_unsigned(125,8) ,
6366	 => std_logic_vector(to_unsigned(128,8) ,
6367	 => std_logic_vector(to_unsigned(121,8) ,
6368	 => std_logic_vector(to_unsigned(124,8) ,
6369	 => std_logic_vector(to_unsigned(133,8) ,
6370	 => std_logic_vector(to_unsigned(128,8) ,
6371	 => std_logic_vector(to_unsigned(124,8) ,
6372	 => std_logic_vector(to_unsigned(128,8) ,
6373	 => std_logic_vector(to_unsigned(131,8) ,
6374	 => std_logic_vector(to_unsigned(125,8) ,
6375	 => std_logic_vector(to_unsigned(133,8) ,
6376	 => std_logic_vector(to_unsigned(134,8) ,
6377	 => std_logic_vector(to_unsigned(136,8) ,
6378	 => std_logic_vector(to_unsigned(144,8) ,
6379	 => std_logic_vector(to_unsigned(144,8) ,
6380	 => std_logic_vector(to_unsigned(141,8) ,
6381	 => std_logic_vector(to_unsigned(144,8) ,
6382	 => std_logic_vector(to_unsigned(147,8) ,
6383	 => std_logic_vector(to_unsigned(152,8) ,
6384	 => std_logic_vector(to_unsigned(152,8) ,
6385	 => std_logic_vector(to_unsigned(154,8) ,
6386	 => std_logic_vector(to_unsigned(156,8) ,
6387	 => std_logic_vector(to_unsigned(154,8) ,
6388	 => std_logic_vector(to_unsigned(154,8) ,
6389	 => std_logic_vector(to_unsigned(159,8) ,
6390	 => std_logic_vector(to_unsigned(154,8) ,
6391	 => std_logic_vector(to_unsigned(152,8) ,
6392	 => std_logic_vector(to_unsigned(154,8) ,
6393	 => std_logic_vector(to_unsigned(159,8) ,
6394	 => std_logic_vector(to_unsigned(152,8) ,
6395	 => std_logic_vector(to_unsigned(151,8) ,
6396	 => std_logic_vector(to_unsigned(152,8) ,
6397	 => std_logic_vector(to_unsigned(152,8) ,
6398	 => std_logic_vector(to_unsigned(156,8) ,
6399	 => std_logic_vector(to_unsigned(159,8) ,
6400	 => std_logic_vector(to_unsigned(159,8) ,
6401	 => std_logic_vector(to_unsigned(85,8) ,
6402	 => std_logic_vector(to_unsigned(77,8) ,
6403	 => std_logic_vector(to_unsigned(73,8) ,
6404	 => std_logic_vector(to_unsigned(79,8) ,
6405	 => std_logic_vector(to_unsigned(77,8) ,
6406	 => std_logic_vector(to_unsigned(74,8) ,
6407	 => std_logic_vector(to_unsigned(73,8) ,
6408	 => std_logic_vector(to_unsigned(77,8) ,
6409	 => std_logic_vector(to_unsigned(78,8) ,
6410	 => std_logic_vector(to_unsigned(76,8) ,
6411	 => std_logic_vector(to_unsigned(70,8) ,
6412	 => std_logic_vector(to_unsigned(72,8) ,
6413	 => std_logic_vector(to_unsigned(76,8) ,
6414	 => std_logic_vector(to_unsigned(72,8) ,
6415	 => std_logic_vector(to_unsigned(65,8) ,
6416	 => std_logic_vector(to_unsigned(74,8) ,
6417	 => std_logic_vector(to_unsigned(74,8) ,
6418	 => std_logic_vector(to_unsigned(74,8) ,
6419	 => std_logic_vector(to_unsigned(76,8) ,
6420	 => std_logic_vector(to_unsigned(74,8) ,
6421	 => std_logic_vector(to_unsigned(72,8) ,
6422	 => std_logic_vector(to_unsigned(71,8) ,
6423	 => std_logic_vector(to_unsigned(72,8) ,
6424	 => std_logic_vector(to_unsigned(69,8) ,
6425	 => std_logic_vector(to_unsigned(67,8) ,
6426	 => std_logic_vector(to_unsigned(72,8) ,
6427	 => std_logic_vector(to_unsigned(72,8) ,
6428	 => std_logic_vector(to_unsigned(77,8) ,
6429	 => std_logic_vector(to_unsigned(77,8) ,
6430	 => std_logic_vector(to_unsigned(68,8) ,
6431	 => std_logic_vector(to_unsigned(70,8) ,
6432	 => std_logic_vector(to_unsigned(77,8) ,
6433	 => std_logic_vector(to_unsigned(73,8) ,
6434	 => std_logic_vector(to_unsigned(76,8) ,
6435	 => std_logic_vector(to_unsigned(79,8) ,
6436	 => std_logic_vector(to_unsigned(76,8) ,
6437	 => std_logic_vector(to_unsigned(78,8) ,
6438	 => std_logic_vector(to_unsigned(79,8) ,
6439	 => std_logic_vector(to_unsigned(84,8) ,
6440	 => std_logic_vector(to_unsigned(86,8) ,
6441	 => std_logic_vector(to_unsigned(85,8) ,
6442	 => std_logic_vector(to_unsigned(82,8) ,
6443	 => std_logic_vector(to_unsigned(88,8) ,
6444	 => std_logic_vector(to_unsigned(91,8) ,
6445	 => std_logic_vector(to_unsigned(90,8) ,
6446	 => std_logic_vector(to_unsigned(91,8) ,
6447	 => std_logic_vector(to_unsigned(95,8) ,
6448	 => std_logic_vector(to_unsigned(97,8) ,
6449	 => std_logic_vector(to_unsigned(96,8) ,
6450	 => std_logic_vector(to_unsigned(97,8) ,
6451	 => std_logic_vector(to_unsigned(99,8) ,
6452	 => std_logic_vector(to_unsigned(103,8) ,
6453	 => std_logic_vector(to_unsigned(105,8) ,
6454	 => std_logic_vector(to_unsigned(108,8) ,
6455	 => std_logic_vector(to_unsigned(112,8) ,
6456	 => std_logic_vector(to_unsigned(112,8) ,
6457	 => std_logic_vector(to_unsigned(109,8) ,
6458	 => std_logic_vector(to_unsigned(109,8) ,
6459	 => std_logic_vector(to_unsigned(107,8) ,
6460	 => std_logic_vector(to_unsigned(104,8) ,
6461	 => std_logic_vector(to_unsigned(101,8) ,
6462	 => std_logic_vector(to_unsigned(99,8) ,
6463	 => std_logic_vector(to_unsigned(103,8) ,
6464	 => std_logic_vector(to_unsigned(104,8) ,
6465	 => std_logic_vector(to_unsigned(107,8) ,
6466	 => std_logic_vector(to_unsigned(111,8) ,
6467	 => std_logic_vector(to_unsigned(109,8) ,
6468	 => std_logic_vector(to_unsigned(109,8) ,
6469	 => std_logic_vector(to_unsigned(105,8) ,
6470	 => std_logic_vector(to_unsigned(103,8) ,
6471	 => std_logic_vector(to_unsigned(111,8) ,
6472	 => std_logic_vector(to_unsigned(111,8) ,
6473	 => std_logic_vector(to_unsigned(109,8) ,
6474	 => std_logic_vector(to_unsigned(111,8) ,
6475	 => std_logic_vector(to_unsigned(105,8) ,
6476	 => std_logic_vector(to_unsigned(103,8) ,
6477	 => std_logic_vector(to_unsigned(109,8) ,
6478	 => std_logic_vector(to_unsigned(107,8) ,
6479	 => std_logic_vector(to_unsigned(103,8) ,
6480	 => std_logic_vector(to_unsigned(96,8) ,
6481	 => std_logic_vector(to_unsigned(95,8) ,
6482	 => std_logic_vector(to_unsigned(99,8) ,
6483	 => std_logic_vector(to_unsigned(97,8) ,
6484	 => std_logic_vector(to_unsigned(93,8) ,
6485	 => std_logic_vector(to_unsigned(93,8) ,
6486	 => std_logic_vector(to_unsigned(96,8) ,
6487	 => std_logic_vector(to_unsigned(96,8) ,
6488	 => std_logic_vector(to_unsigned(101,8) ,
6489	 => std_logic_vector(to_unsigned(105,8) ,
6490	 => std_logic_vector(to_unsigned(104,8) ,
6491	 => std_logic_vector(to_unsigned(95,8) ,
6492	 => std_logic_vector(to_unsigned(90,8) ,
6493	 => std_logic_vector(to_unsigned(85,8) ,
6494	 => std_logic_vector(to_unsigned(85,8) ,
6495	 => std_logic_vector(to_unsigned(90,8) ,
6496	 => std_logic_vector(to_unsigned(86,8) ,
6497	 => std_logic_vector(to_unsigned(86,8) ,
6498	 => std_logic_vector(to_unsigned(85,8) ,
6499	 => std_logic_vector(to_unsigned(82,8) ,
6500	 => std_logic_vector(to_unsigned(79,8) ,
6501	 => std_logic_vector(to_unsigned(79,8) ,
6502	 => std_logic_vector(to_unsigned(82,8) ,
6503	 => std_logic_vector(to_unsigned(80,8) ,
6504	 => std_logic_vector(to_unsigned(68,8) ,
6505	 => std_logic_vector(to_unsigned(69,8) ,
6506	 => std_logic_vector(to_unsigned(71,8) ,
6507	 => std_logic_vector(to_unsigned(72,8) ,
6508	 => std_logic_vector(to_unsigned(74,8) ,
6509	 => std_logic_vector(to_unsigned(72,8) ,
6510	 => std_logic_vector(to_unsigned(69,8) ,
6511	 => std_logic_vector(to_unsigned(72,8) ,
6512	 => std_logic_vector(to_unsigned(69,8) ,
6513	 => std_logic_vector(to_unsigned(78,8) ,
6514	 => std_logic_vector(to_unsigned(86,8) ,
6515	 => std_logic_vector(to_unsigned(84,8) ,
6516	 => std_logic_vector(to_unsigned(77,8) ,
6517	 => std_logic_vector(to_unsigned(80,8) ,
6518	 => std_logic_vector(to_unsigned(87,8) ,
6519	 => std_logic_vector(to_unsigned(88,8) ,
6520	 => std_logic_vector(to_unsigned(86,8) ,
6521	 => std_logic_vector(to_unsigned(87,8) ,
6522	 => std_logic_vector(to_unsigned(87,8) ,
6523	 => std_logic_vector(to_unsigned(88,8) ,
6524	 => std_logic_vector(to_unsigned(96,8) ,
6525	 => std_logic_vector(to_unsigned(96,8) ,
6526	 => std_logic_vector(to_unsigned(91,8) ,
6527	 => std_logic_vector(to_unsigned(91,8) ,
6528	 => std_logic_vector(to_unsigned(95,8) ,
6529	 => std_logic_vector(to_unsigned(96,8) ,
6530	 => std_logic_vector(to_unsigned(92,8) ,
6531	 => std_logic_vector(to_unsigned(92,8) ,
6532	 => std_logic_vector(to_unsigned(87,8) ,
6533	 => std_logic_vector(to_unsigned(86,8) ,
6534	 => std_logic_vector(to_unsigned(86,8) ,
6535	 => std_logic_vector(to_unsigned(86,8) ,
6536	 => std_logic_vector(to_unsigned(87,8) ,
6537	 => std_logic_vector(to_unsigned(84,8) ,
6538	 => std_logic_vector(to_unsigned(84,8) ,
6539	 => std_logic_vector(to_unsigned(90,8) ,
6540	 => std_logic_vector(to_unsigned(90,8) ,
6541	 => std_logic_vector(to_unsigned(91,8) ,
6542	 => std_logic_vector(to_unsigned(95,8) ,
6543	 => std_logic_vector(to_unsigned(93,8) ,
6544	 => std_logic_vector(to_unsigned(90,8) ,
6545	 => std_logic_vector(to_unsigned(96,8) ,
6546	 => std_logic_vector(to_unsigned(99,8) ,
6547	 => std_logic_vector(to_unsigned(88,8) ,
6548	 => std_logic_vector(to_unsigned(87,8) ,
6549	 => std_logic_vector(to_unsigned(90,8) ,
6550	 => std_logic_vector(to_unsigned(87,8) ,
6551	 => std_logic_vector(to_unsigned(91,8) ,
6552	 => std_logic_vector(to_unsigned(88,8) ,
6553	 => std_logic_vector(to_unsigned(87,8) ,
6554	 => std_logic_vector(to_unsigned(88,8) ,
6555	 => std_logic_vector(to_unsigned(88,8) ,
6556	 => std_logic_vector(to_unsigned(87,8) ,
6557	 => std_logic_vector(to_unsigned(87,8) ,
6558	 => std_logic_vector(to_unsigned(88,8) ,
6559	 => std_logic_vector(to_unsigned(87,8) ,
6560	 => std_logic_vector(to_unsigned(82,8) ,
6561	 => std_logic_vector(to_unsigned(87,8) ,
6562	 => std_logic_vector(to_unsigned(90,8) ,
6563	 => std_logic_vector(to_unsigned(86,8) ,
6564	 => std_logic_vector(to_unsigned(87,8) ,
6565	 => std_logic_vector(to_unsigned(88,8) ,
6566	 => std_logic_vector(to_unsigned(87,8) ,
6567	 => std_logic_vector(to_unsigned(86,8) ,
6568	 => std_logic_vector(to_unsigned(84,8) ,
6569	 => std_logic_vector(to_unsigned(86,8) ,
6570	 => std_logic_vector(to_unsigned(82,8) ,
6571	 => std_logic_vector(to_unsigned(87,8) ,
6572	 => std_logic_vector(to_unsigned(90,8) ,
6573	 => std_logic_vector(to_unsigned(84,8) ,
6574	 => std_logic_vector(to_unsigned(84,8) ,
6575	 => std_logic_vector(to_unsigned(88,8) ,
6576	 => std_logic_vector(to_unsigned(81,8) ,
6577	 => std_logic_vector(to_unsigned(82,8) ,
6578	 => std_logic_vector(to_unsigned(78,8) ,
6579	 => std_logic_vector(to_unsigned(73,8) ,
6580	 => std_logic_vector(to_unsigned(74,8) ,
6581	 => std_logic_vector(to_unsigned(77,8) ,
6582	 => std_logic_vector(to_unsigned(84,8) ,
6583	 => std_logic_vector(to_unsigned(82,8) ,
6584	 => std_logic_vector(to_unsigned(78,8) ,
6585	 => std_logic_vector(to_unsigned(80,8) ,
6586	 => std_logic_vector(to_unsigned(78,8) ,
6587	 => std_logic_vector(to_unsigned(86,8) ,
6588	 => std_logic_vector(to_unsigned(90,8) ,
6589	 => std_logic_vector(to_unsigned(82,8) ,
6590	 => std_logic_vector(to_unsigned(87,8) ,
6591	 => std_logic_vector(to_unsigned(87,8) ,
6592	 => std_logic_vector(to_unsigned(72,8) ,
6593	 => std_logic_vector(to_unsigned(64,8) ,
6594	 => std_logic_vector(to_unsigned(62,8) ,
6595	 => std_logic_vector(to_unsigned(64,8) ,
6596	 => std_logic_vector(to_unsigned(76,8) ,
6597	 => std_logic_vector(to_unsigned(73,8) ,
6598	 => std_logic_vector(to_unsigned(74,8) ,
6599	 => std_logic_vector(to_unsigned(77,8) ,
6600	 => std_logic_vector(to_unsigned(80,8) ,
6601	 => std_logic_vector(to_unsigned(66,8) ,
6602	 => std_logic_vector(to_unsigned(57,8) ,
6603	 => std_logic_vector(to_unsigned(61,8) ,
6604	 => std_logic_vector(to_unsigned(63,8) ,
6605	 => std_logic_vector(to_unsigned(63,8) ,
6606	 => std_logic_vector(to_unsigned(65,8) ,
6607	 => std_logic_vector(to_unsigned(74,8) ,
6608	 => std_logic_vector(to_unsigned(73,8) ,
6609	 => std_logic_vector(to_unsigned(63,8) ,
6610	 => std_logic_vector(to_unsigned(66,8) ,
6611	 => std_logic_vector(to_unsigned(69,8) ,
6612	 => std_logic_vector(to_unsigned(65,8) ,
6613	 => std_logic_vector(to_unsigned(66,8) ,
6614	 => std_logic_vector(to_unsigned(69,8) ,
6615	 => std_logic_vector(to_unsigned(69,8) ,
6616	 => std_logic_vector(to_unsigned(71,8) ,
6617	 => std_logic_vector(to_unsigned(71,8) ,
6618	 => std_logic_vector(to_unsigned(71,8) ,
6619	 => std_logic_vector(to_unsigned(69,8) ,
6620	 => std_logic_vector(to_unsigned(65,8) ,
6621	 => std_logic_vector(to_unsigned(60,8) ,
6622	 => std_logic_vector(to_unsigned(56,8) ,
6623	 => std_logic_vector(to_unsigned(62,8) ,
6624	 => std_logic_vector(to_unsigned(65,8) ,
6625	 => std_logic_vector(to_unsigned(68,8) ,
6626	 => std_logic_vector(to_unsigned(67,8) ,
6627	 => std_logic_vector(to_unsigned(65,8) ,
6628	 => std_logic_vector(to_unsigned(58,8) ,
6629	 => std_logic_vector(to_unsigned(62,8) ,
6630	 => std_logic_vector(to_unsigned(66,8) ,
6631	 => std_logic_vector(to_unsigned(68,8) ,
6632	 => std_logic_vector(to_unsigned(57,8) ,
6633	 => std_logic_vector(to_unsigned(54,8) ,
6634	 => std_logic_vector(to_unsigned(57,8) ,
6635	 => std_logic_vector(to_unsigned(51,8) ,
6636	 => std_logic_vector(to_unsigned(46,8) ,
6637	 => std_logic_vector(to_unsigned(49,8) ,
6638	 => std_logic_vector(to_unsigned(49,8) ,
6639	 => std_logic_vector(to_unsigned(52,8) ,
6640	 => std_logic_vector(to_unsigned(7,8) ,
6641	 => std_logic_vector(to_unsigned(0,8) ,
6642	 => std_logic_vector(to_unsigned(0,8) ,
6643	 => std_logic_vector(to_unsigned(11,8) ,
6644	 => std_logic_vector(to_unsigned(81,8) ,
6645	 => std_logic_vector(to_unsigned(72,8) ,
6646	 => std_logic_vector(to_unsigned(72,8) ,
6647	 => std_logic_vector(to_unsigned(73,8) ,
6648	 => std_logic_vector(to_unsigned(74,8) ,
6649	 => std_logic_vector(to_unsigned(84,8) ,
6650	 => std_logic_vector(to_unsigned(81,8) ,
6651	 => std_logic_vector(to_unsigned(84,8) ,
6652	 => std_logic_vector(to_unsigned(88,8) ,
6653	 => std_logic_vector(to_unsigned(85,8) ,
6654	 => std_logic_vector(to_unsigned(88,8) ,
6655	 => std_logic_vector(to_unsigned(86,8) ,
6656	 => std_logic_vector(to_unsigned(84,8) ,
6657	 => std_logic_vector(to_unsigned(78,8) ,
6658	 => std_logic_vector(to_unsigned(80,8) ,
6659	 => std_logic_vector(to_unsigned(86,8) ,
6660	 => std_logic_vector(to_unsigned(87,8) ,
6661	 => std_logic_vector(to_unsigned(86,8) ,
6662	 => std_logic_vector(to_unsigned(84,8) ,
6663	 => std_logic_vector(to_unsigned(82,8) ,
6664	 => std_logic_vector(to_unsigned(79,8) ,
6665	 => std_logic_vector(to_unsigned(84,8) ,
6666	 => std_logic_vector(to_unsigned(85,8) ,
6667	 => std_logic_vector(to_unsigned(82,8) ,
6668	 => std_logic_vector(to_unsigned(93,8) ,
6669	 => std_logic_vector(to_unsigned(95,8) ,
6670	 => std_logic_vector(to_unsigned(99,8) ,
6671	 => std_logic_vector(to_unsigned(96,8) ,
6672	 => std_logic_vector(to_unsigned(93,8) ,
6673	 => std_logic_vector(to_unsigned(101,8) ,
6674	 => std_logic_vector(to_unsigned(91,8) ,
6675	 => std_logic_vector(to_unsigned(90,8) ,
6676	 => std_logic_vector(to_unsigned(96,8) ,
6677	 => std_logic_vector(to_unsigned(97,8) ,
6678	 => std_logic_vector(to_unsigned(95,8) ,
6679	 => std_logic_vector(to_unsigned(99,8) ,
6680	 => std_logic_vector(to_unsigned(107,8) ,
6681	 => std_logic_vector(to_unsigned(127,8) ,
6682	 => std_logic_vector(to_unsigned(127,8) ,
6683	 => std_logic_vector(to_unsigned(119,8) ,
6684	 => std_logic_vector(to_unsigned(121,8) ,
6685	 => std_logic_vector(to_unsigned(124,8) ,
6686	 => std_logic_vector(to_unsigned(128,8) ,
6687	 => std_logic_vector(to_unsigned(115,8) ,
6688	 => std_logic_vector(to_unsigned(111,8) ,
6689	 => std_logic_vector(to_unsigned(122,8) ,
6690	 => std_logic_vector(to_unsigned(133,8) ,
6691	 => std_logic_vector(to_unsigned(128,8) ,
6692	 => std_logic_vector(to_unsigned(122,8) ,
6693	 => std_logic_vector(to_unsigned(128,8) ,
6694	 => std_logic_vector(to_unsigned(128,8) ,
6695	 => std_logic_vector(to_unsigned(134,8) ,
6696	 => std_logic_vector(to_unsigned(138,8) ,
6697	 => std_logic_vector(to_unsigned(146,8) ,
6698	 => std_logic_vector(to_unsigned(147,8) ,
6699	 => std_logic_vector(to_unsigned(147,8) ,
6700	 => std_logic_vector(to_unsigned(147,8) ,
6701	 => std_logic_vector(to_unsigned(147,8) ,
6702	 => std_logic_vector(to_unsigned(147,8) ,
6703	 => std_logic_vector(to_unsigned(152,8) ,
6704	 => std_logic_vector(to_unsigned(152,8) ,
6705	 => std_logic_vector(to_unsigned(154,8) ,
6706	 => std_logic_vector(to_unsigned(152,8) ,
6707	 => std_logic_vector(to_unsigned(152,8) ,
6708	 => std_logic_vector(to_unsigned(151,8) ,
6709	 => std_logic_vector(to_unsigned(154,8) ,
6710	 => std_logic_vector(to_unsigned(157,8) ,
6711	 => std_logic_vector(to_unsigned(156,8) ,
6712	 => std_logic_vector(to_unsigned(154,8) ,
6713	 => std_logic_vector(to_unsigned(152,8) ,
6714	 => std_logic_vector(to_unsigned(156,8) ,
6715	 => std_logic_vector(to_unsigned(152,8) ,
6716	 => std_logic_vector(to_unsigned(152,8) ,
6717	 => std_logic_vector(to_unsigned(152,8) ,
6718	 => std_logic_vector(to_unsigned(154,8) ,
6719	 => std_logic_vector(to_unsigned(154,8) ,
6720	 => std_logic_vector(to_unsigned(152,8) ,
6721	 => std_logic_vector(to_unsigned(84,8) ,
6722	 => std_logic_vector(to_unsigned(74,8) ,
6723	 => std_logic_vector(to_unsigned(74,8) ,
6724	 => std_logic_vector(to_unsigned(80,8) ,
6725	 => std_logic_vector(to_unsigned(78,8) ,
6726	 => std_logic_vector(to_unsigned(72,8) ,
6727	 => std_logic_vector(to_unsigned(72,8) ,
6728	 => std_logic_vector(to_unsigned(71,8) ,
6729	 => std_logic_vector(to_unsigned(68,8) ,
6730	 => std_logic_vector(to_unsigned(72,8) ,
6731	 => std_logic_vector(to_unsigned(72,8) ,
6732	 => std_logic_vector(to_unsigned(71,8) ,
6733	 => std_logic_vector(to_unsigned(70,8) ,
6734	 => std_logic_vector(to_unsigned(72,8) ,
6735	 => std_logic_vector(to_unsigned(69,8) ,
6736	 => std_logic_vector(to_unsigned(68,8) ,
6737	 => std_logic_vector(to_unsigned(76,8) ,
6738	 => std_logic_vector(to_unsigned(76,8) ,
6739	 => std_logic_vector(to_unsigned(77,8) ,
6740	 => std_logic_vector(to_unsigned(76,8) ,
6741	 => std_logic_vector(to_unsigned(71,8) ,
6742	 => std_logic_vector(to_unsigned(70,8) ,
6743	 => std_logic_vector(to_unsigned(69,8) ,
6744	 => std_logic_vector(to_unsigned(70,8) ,
6745	 => std_logic_vector(to_unsigned(76,8) ,
6746	 => std_logic_vector(to_unsigned(74,8) ,
6747	 => std_logic_vector(to_unsigned(69,8) ,
6748	 => std_logic_vector(to_unsigned(73,8) ,
6749	 => std_logic_vector(to_unsigned(80,8) ,
6750	 => std_logic_vector(to_unsigned(74,8) ,
6751	 => std_logic_vector(to_unsigned(76,8) ,
6752	 => std_logic_vector(to_unsigned(72,8) ,
6753	 => std_logic_vector(to_unsigned(74,8) ,
6754	 => std_logic_vector(to_unsigned(74,8) ,
6755	 => std_logic_vector(to_unsigned(74,8) ,
6756	 => std_logic_vector(to_unsigned(78,8) ,
6757	 => std_logic_vector(to_unsigned(73,8) ,
6758	 => std_logic_vector(to_unsigned(77,8) ,
6759	 => std_logic_vector(to_unsigned(82,8) ,
6760	 => std_logic_vector(to_unsigned(81,8) ,
6761	 => std_logic_vector(to_unsigned(85,8) ,
6762	 => std_logic_vector(to_unsigned(87,8) ,
6763	 => std_logic_vector(to_unsigned(90,8) ,
6764	 => std_logic_vector(to_unsigned(86,8) ,
6765	 => std_logic_vector(to_unsigned(87,8) ,
6766	 => std_logic_vector(to_unsigned(91,8) ,
6767	 => std_logic_vector(to_unsigned(93,8) ,
6768	 => std_logic_vector(to_unsigned(92,8) ,
6769	 => std_logic_vector(to_unsigned(95,8) ,
6770	 => std_logic_vector(to_unsigned(101,8) ,
6771	 => std_logic_vector(to_unsigned(101,8) ,
6772	 => std_logic_vector(to_unsigned(100,8) ,
6773	 => std_logic_vector(to_unsigned(103,8) ,
6774	 => std_logic_vector(to_unsigned(101,8) ,
6775	 => std_logic_vector(to_unsigned(105,8) ,
6776	 => std_logic_vector(to_unsigned(103,8) ,
6777	 => std_logic_vector(to_unsigned(101,8) ,
6778	 => std_logic_vector(to_unsigned(104,8) ,
6779	 => std_logic_vector(to_unsigned(104,8) ,
6780	 => std_logic_vector(to_unsigned(100,8) ,
6781	 => std_logic_vector(to_unsigned(97,8) ,
6782	 => std_logic_vector(to_unsigned(96,8) ,
6783	 => std_logic_vector(to_unsigned(101,8) ,
6784	 => std_logic_vector(to_unsigned(103,8) ,
6785	 => std_logic_vector(to_unsigned(103,8) ,
6786	 => std_logic_vector(to_unsigned(109,8) ,
6787	 => std_logic_vector(to_unsigned(108,8) ,
6788	 => std_logic_vector(to_unsigned(105,8) ,
6789	 => std_logic_vector(to_unsigned(111,8) ,
6790	 => std_logic_vector(to_unsigned(108,8) ,
6791	 => std_logic_vector(to_unsigned(108,8) ,
6792	 => std_logic_vector(to_unsigned(108,8) ,
6793	 => std_logic_vector(to_unsigned(108,8) ,
6794	 => std_logic_vector(to_unsigned(114,8) ,
6795	 => std_logic_vector(to_unsigned(109,8) ,
6796	 => std_logic_vector(to_unsigned(105,8) ,
6797	 => std_logic_vector(to_unsigned(111,8) ,
6798	 => std_logic_vector(to_unsigned(109,8) ,
6799	 => std_logic_vector(to_unsigned(108,8) ,
6800	 => std_logic_vector(to_unsigned(101,8) ,
6801	 => std_logic_vector(to_unsigned(100,8) ,
6802	 => std_logic_vector(to_unsigned(93,8) ,
6803	 => std_logic_vector(to_unsigned(96,8) ,
6804	 => std_logic_vector(to_unsigned(96,8) ,
6805	 => std_logic_vector(to_unsigned(95,8) ,
6806	 => std_logic_vector(to_unsigned(92,8) ,
6807	 => std_logic_vector(to_unsigned(88,8) ,
6808	 => std_logic_vector(to_unsigned(93,8) ,
6809	 => std_logic_vector(to_unsigned(99,8) ,
6810	 => std_logic_vector(to_unsigned(101,8) ,
6811	 => std_logic_vector(to_unsigned(97,8) ,
6812	 => std_logic_vector(to_unsigned(91,8) ,
6813	 => std_logic_vector(to_unsigned(87,8) ,
6814	 => std_logic_vector(to_unsigned(86,8) ,
6815	 => std_logic_vector(to_unsigned(90,8) ,
6816	 => std_logic_vector(to_unsigned(86,8) ,
6817	 => std_logic_vector(to_unsigned(88,8) ,
6818	 => std_logic_vector(to_unsigned(84,8) ,
6819	 => std_logic_vector(to_unsigned(81,8) ,
6820	 => std_logic_vector(to_unsigned(79,8) ,
6821	 => std_logic_vector(to_unsigned(79,8) ,
6822	 => std_logic_vector(to_unsigned(84,8) ,
6823	 => std_logic_vector(to_unsigned(76,8) ,
6824	 => std_logic_vector(to_unsigned(73,8) ,
6825	 => std_logic_vector(to_unsigned(78,8) ,
6826	 => std_logic_vector(to_unsigned(74,8) ,
6827	 => std_logic_vector(to_unsigned(76,8) ,
6828	 => std_logic_vector(to_unsigned(78,8) ,
6829	 => std_logic_vector(to_unsigned(76,8) ,
6830	 => std_logic_vector(to_unsigned(68,8) ,
6831	 => std_logic_vector(to_unsigned(71,8) ,
6832	 => std_logic_vector(to_unsigned(74,8) ,
6833	 => std_logic_vector(to_unsigned(78,8) ,
6834	 => std_logic_vector(to_unsigned(82,8) ,
6835	 => std_logic_vector(to_unsigned(82,8) ,
6836	 => std_logic_vector(to_unsigned(81,8) ,
6837	 => std_logic_vector(to_unsigned(84,8) ,
6838	 => std_logic_vector(to_unsigned(86,8) ,
6839	 => std_logic_vector(to_unsigned(87,8) ,
6840	 => std_logic_vector(to_unsigned(90,8) ,
6841	 => std_logic_vector(to_unsigned(86,8) ,
6842	 => std_logic_vector(to_unsigned(87,8) ,
6843	 => std_logic_vector(to_unsigned(88,8) ,
6844	 => std_logic_vector(to_unsigned(96,8) ,
6845	 => std_logic_vector(to_unsigned(97,8) ,
6846	 => std_logic_vector(to_unsigned(93,8) ,
6847	 => std_logic_vector(to_unsigned(91,8) ,
6848	 => std_logic_vector(to_unsigned(95,8) ,
6849	 => std_logic_vector(to_unsigned(97,8) ,
6850	 => std_logic_vector(to_unsigned(92,8) ,
6851	 => std_logic_vector(to_unsigned(96,8) ,
6852	 => std_logic_vector(to_unsigned(99,8) ,
6853	 => std_logic_vector(to_unsigned(95,8) ,
6854	 => std_logic_vector(to_unsigned(90,8) ,
6855	 => std_logic_vector(to_unsigned(85,8) ,
6856	 => std_logic_vector(to_unsigned(88,8) ,
6857	 => std_logic_vector(to_unsigned(88,8) ,
6858	 => std_logic_vector(to_unsigned(92,8) ,
6859	 => std_logic_vector(to_unsigned(97,8) ,
6860	 => std_logic_vector(to_unsigned(96,8) ,
6861	 => std_logic_vector(to_unsigned(95,8) ,
6862	 => std_logic_vector(to_unsigned(95,8) ,
6863	 => std_logic_vector(to_unsigned(97,8) ,
6864	 => std_logic_vector(to_unsigned(104,8) ,
6865	 => std_logic_vector(to_unsigned(107,8) ,
6866	 => std_logic_vector(to_unsigned(101,8) ,
6867	 => std_logic_vector(to_unsigned(96,8) ,
6868	 => std_logic_vector(to_unsigned(97,8) ,
6869	 => std_logic_vector(to_unsigned(95,8) ,
6870	 => std_logic_vector(to_unsigned(91,8) ,
6871	 => std_logic_vector(to_unsigned(95,8) ,
6872	 => std_logic_vector(to_unsigned(97,8) ,
6873	 => std_logic_vector(to_unsigned(93,8) ,
6874	 => std_logic_vector(to_unsigned(92,8) ,
6875	 => std_logic_vector(to_unsigned(97,8) ,
6876	 => std_logic_vector(to_unsigned(101,8) ,
6877	 => std_logic_vector(to_unsigned(99,8) ,
6878	 => std_logic_vector(to_unsigned(96,8) ,
6879	 => std_logic_vector(to_unsigned(97,8) ,
6880	 => std_logic_vector(to_unsigned(101,8) ,
6881	 => std_logic_vector(to_unsigned(100,8) ,
6882	 => std_logic_vector(to_unsigned(90,8) ,
6883	 => std_logic_vector(to_unsigned(90,8) ,
6884	 => std_logic_vector(to_unsigned(92,8) ,
6885	 => std_logic_vector(to_unsigned(92,8) ,
6886	 => std_logic_vector(to_unsigned(93,8) ,
6887	 => std_logic_vector(to_unsigned(93,8) ,
6888	 => std_logic_vector(to_unsigned(90,8) ,
6889	 => std_logic_vector(to_unsigned(93,8) ,
6890	 => std_logic_vector(to_unsigned(92,8) ,
6891	 => std_logic_vector(to_unsigned(91,8) ,
6892	 => std_logic_vector(to_unsigned(87,8) ,
6893	 => std_logic_vector(to_unsigned(86,8) ,
6894	 => std_logic_vector(to_unsigned(90,8) ,
6895	 => std_logic_vector(to_unsigned(90,8) ,
6896	 => std_logic_vector(to_unsigned(82,8) ,
6897	 => std_logic_vector(to_unsigned(88,8) ,
6898	 => std_logic_vector(to_unsigned(85,8) ,
6899	 => std_logic_vector(to_unsigned(84,8) ,
6900	 => std_logic_vector(to_unsigned(84,8) ,
6901	 => std_logic_vector(to_unsigned(82,8) ,
6902	 => std_logic_vector(to_unsigned(80,8) ,
6903	 => std_logic_vector(to_unsigned(78,8) ,
6904	 => std_logic_vector(to_unsigned(84,8) ,
6905	 => std_logic_vector(to_unsigned(85,8) ,
6906	 => std_logic_vector(to_unsigned(81,8) ,
6907	 => std_logic_vector(to_unsigned(79,8) ,
6908	 => std_logic_vector(to_unsigned(88,8) ,
6909	 => std_logic_vector(to_unsigned(84,8) ,
6910	 => std_logic_vector(to_unsigned(84,8) ,
6911	 => std_logic_vector(to_unsigned(81,8) ,
6912	 => std_logic_vector(to_unsigned(63,8) ,
6913	 => std_logic_vector(to_unsigned(53,8) ,
6914	 => std_logic_vector(to_unsigned(59,8) ,
6915	 => std_logic_vector(to_unsigned(56,8) ,
6916	 => std_logic_vector(to_unsigned(60,8) ,
6917	 => std_logic_vector(to_unsigned(65,8) ,
6918	 => std_logic_vector(to_unsigned(59,8) ,
6919	 => std_logic_vector(to_unsigned(62,8) ,
6920	 => std_logic_vector(to_unsigned(68,8) ,
6921	 => std_logic_vector(to_unsigned(62,8) ,
6922	 => std_logic_vector(to_unsigned(59,8) ,
6923	 => std_logic_vector(to_unsigned(67,8) ,
6924	 => std_logic_vector(to_unsigned(66,8) ,
6925	 => std_logic_vector(to_unsigned(61,8) ,
6926	 => std_logic_vector(to_unsigned(64,8) ,
6927	 => std_logic_vector(to_unsigned(66,8) ,
6928	 => std_logic_vector(to_unsigned(65,8) ,
6929	 => std_logic_vector(to_unsigned(70,8) ,
6930	 => std_logic_vector(to_unsigned(71,8) ,
6931	 => std_logic_vector(to_unsigned(68,8) ,
6932	 => std_logic_vector(to_unsigned(61,8) ,
6933	 => std_logic_vector(to_unsigned(68,8) ,
6934	 => std_logic_vector(to_unsigned(67,8) ,
6935	 => std_logic_vector(to_unsigned(61,8) ,
6936	 => std_logic_vector(to_unsigned(69,8) ,
6937	 => std_logic_vector(to_unsigned(68,8) ,
6938	 => std_logic_vector(to_unsigned(69,8) ,
6939	 => std_logic_vector(to_unsigned(63,8) ,
6940	 => std_logic_vector(to_unsigned(67,8) ,
6941	 => std_logic_vector(to_unsigned(70,8) ,
6942	 => std_logic_vector(to_unsigned(67,8) ,
6943	 => std_logic_vector(to_unsigned(64,8) ,
6944	 => std_logic_vector(to_unsigned(65,8) ,
6945	 => std_logic_vector(to_unsigned(70,8) ,
6946	 => std_logic_vector(to_unsigned(66,8) ,
6947	 => std_logic_vector(to_unsigned(65,8) ,
6948	 => std_logic_vector(to_unsigned(61,8) ,
6949	 => std_logic_vector(to_unsigned(58,8) ,
6950	 => std_logic_vector(to_unsigned(58,8) ,
6951	 => std_logic_vector(to_unsigned(64,8) ,
6952	 => std_logic_vector(to_unsigned(58,8) ,
6953	 => std_logic_vector(to_unsigned(55,8) ,
6954	 => std_logic_vector(to_unsigned(58,8) ,
6955	 => std_logic_vector(to_unsigned(55,8) ,
6956	 => std_logic_vector(to_unsigned(53,8) ,
6957	 => std_logic_vector(to_unsigned(60,8) ,
6958	 => std_logic_vector(to_unsigned(57,8) ,
6959	 => std_logic_vector(to_unsigned(66,8) ,
6960	 => std_logic_vector(to_unsigned(20,8) ,
6961	 => std_logic_vector(to_unsigned(1,8) ,
6962	 => std_logic_vector(to_unsigned(0,8) ,
6963	 => std_logic_vector(to_unsigned(4,8) ,
6964	 => std_logic_vector(to_unsigned(62,8) ,
6965	 => std_logic_vector(to_unsigned(77,8) ,
6966	 => std_logic_vector(to_unsigned(71,8) ,
6967	 => std_logic_vector(to_unsigned(74,8) ,
6968	 => std_logic_vector(to_unsigned(79,8) ,
6969	 => std_logic_vector(to_unsigned(88,8) ,
6970	 => std_logic_vector(to_unsigned(82,8) ,
6971	 => std_logic_vector(to_unsigned(84,8) ,
6972	 => std_logic_vector(to_unsigned(86,8) ,
6973	 => std_logic_vector(to_unsigned(85,8) ,
6974	 => std_logic_vector(to_unsigned(87,8) ,
6975	 => std_logic_vector(to_unsigned(84,8) ,
6976	 => std_logic_vector(to_unsigned(78,8) ,
6977	 => std_logic_vector(to_unsigned(74,8) ,
6978	 => std_logic_vector(to_unsigned(81,8) ,
6979	 => std_logic_vector(to_unsigned(101,8) ,
6980	 => std_logic_vector(to_unsigned(103,8) ,
6981	 => std_logic_vector(to_unsigned(95,8) ,
6982	 => std_logic_vector(to_unsigned(92,8) ,
6983	 => std_logic_vector(to_unsigned(85,8) ,
6984	 => std_logic_vector(to_unsigned(82,8) ,
6985	 => std_logic_vector(to_unsigned(92,8) ,
6986	 => std_logic_vector(to_unsigned(95,8) ,
6987	 => std_logic_vector(to_unsigned(88,8) ,
6988	 => std_logic_vector(to_unsigned(96,8) ,
6989	 => std_logic_vector(to_unsigned(88,8) ,
6990	 => std_logic_vector(to_unsigned(88,8) ,
6991	 => std_logic_vector(to_unsigned(92,8) ,
6992	 => std_logic_vector(to_unsigned(95,8) ,
6993	 => std_logic_vector(to_unsigned(92,8) ,
6994	 => std_logic_vector(to_unsigned(90,8) ,
6995	 => std_logic_vector(to_unsigned(95,8) ,
6996	 => std_logic_vector(to_unsigned(93,8) ,
6997	 => std_logic_vector(to_unsigned(100,8) ,
6998	 => std_logic_vector(to_unsigned(100,8) ,
6999	 => std_logic_vector(to_unsigned(101,8) ,
7000	 => std_logic_vector(to_unsigned(112,8) ,
7001	 => std_logic_vector(to_unsigned(131,8) ,
7002	 => std_logic_vector(to_unsigned(130,8) ,
7003	 => std_logic_vector(to_unsigned(125,8) ,
7004	 => std_logic_vector(to_unsigned(112,8) ,
7005	 => std_logic_vector(to_unsigned(107,8) ,
7006	 => std_logic_vector(to_unsigned(114,8) ,
7007	 => std_logic_vector(to_unsigned(115,8) ,
7008	 => std_logic_vector(to_unsigned(114,8) ,
7009	 => std_logic_vector(to_unsigned(121,8) ,
7010	 => std_logic_vector(to_unsigned(128,8) ,
7011	 => std_logic_vector(to_unsigned(128,8) ,
7012	 => std_logic_vector(to_unsigned(124,8) ,
7013	 => std_logic_vector(to_unsigned(121,8) ,
7014	 => std_logic_vector(to_unsigned(131,8) ,
7015	 => std_logic_vector(to_unsigned(139,8) ,
7016	 => std_logic_vector(to_unsigned(136,8) ,
7017	 => std_logic_vector(to_unsigned(136,8) ,
7018	 => std_logic_vector(to_unsigned(142,8) ,
7019	 => std_logic_vector(to_unsigned(146,8) ,
7020	 => std_logic_vector(to_unsigned(146,8) ,
7021	 => std_logic_vector(to_unsigned(146,8) ,
7022	 => std_logic_vector(to_unsigned(146,8) ,
7023	 => std_logic_vector(to_unsigned(147,8) ,
7024	 => std_logic_vector(to_unsigned(147,8) ,
7025	 => std_logic_vector(to_unsigned(149,8) ,
7026	 => std_logic_vector(to_unsigned(147,8) ,
7027	 => std_logic_vector(to_unsigned(151,8) ,
7028	 => std_logic_vector(to_unsigned(149,8) ,
7029	 => std_logic_vector(to_unsigned(149,8) ,
7030	 => std_logic_vector(to_unsigned(154,8) ,
7031	 => std_logic_vector(to_unsigned(151,8) ,
7032	 => std_logic_vector(to_unsigned(147,8) ,
7033	 => std_logic_vector(to_unsigned(144,8) ,
7034	 => std_logic_vector(to_unsigned(151,8) ,
7035	 => std_logic_vector(to_unsigned(149,8) ,
7036	 => std_logic_vector(to_unsigned(152,8) ,
7037	 => std_logic_vector(to_unsigned(154,8) ,
7038	 => std_logic_vector(to_unsigned(151,8) ,
7039	 => std_logic_vector(to_unsigned(151,8) ,
7040	 => std_logic_vector(to_unsigned(152,8) ,
7041	 => std_logic_vector(to_unsigned(81,8) ,
7042	 => std_logic_vector(to_unsigned(77,8) ,
7043	 => std_logic_vector(to_unsigned(77,8) ,
7044	 => std_logic_vector(to_unsigned(82,8) ,
7045	 => std_logic_vector(to_unsigned(81,8) ,
7046	 => std_logic_vector(to_unsigned(72,8) ,
7047	 => std_logic_vector(to_unsigned(67,8) ,
7048	 => std_logic_vector(to_unsigned(69,8) ,
7049	 => std_logic_vector(to_unsigned(71,8) ,
7050	 => std_logic_vector(to_unsigned(73,8) ,
7051	 => std_logic_vector(to_unsigned(70,8) ,
7052	 => std_logic_vector(to_unsigned(72,8) ,
7053	 => std_logic_vector(to_unsigned(72,8) ,
7054	 => std_logic_vector(to_unsigned(72,8) ,
7055	 => std_logic_vector(to_unsigned(79,8) ,
7056	 => std_logic_vector(to_unsigned(72,8) ,
7057	 => std_logic_vector(to_unsigned(74,8) ,
7058	 => std_logic_vector(to_unsigned(71,8) ,
7059	 => std_logic_vector(to_unsigned(73,8) ,
7060	 => std_logic_vector(to_unsigned(72,8) ,
7061	 => std_logic_vector(to_unsigned(69,8) ,
7062	 => std_logic_vector(to_unsigned(74,8) ,
7063	 => std_logic_vector(to_unsigned(68,8) ,
7064	 => std_logic_vector(to_unsigned(68,8) ,
7065	 => std_logic_vector(to_unsigned(74,8) ,
7066	 => std_logic_vector(to_unsigned(77,8) ,
7067	 => std_logic_vector(to_unsigned(76,8) ,
7068	 => std_logic_vector(to_unsigned(72,8) ,
7069	 => std_logic_vector(to_unsigned(73,8) ,
7070	 => std_logic_vector(to_unsigned(73,8) ,
7071	 => std_logic_vector(to_unsigned(78,8) ,
7072	 => std_logic_vector(to_unsigned(70,8) ,
7073	 => std_logic_vector(to_unsigned(69,8) ,
7074	 => std_logic_vector(to_unsigned(73,8) ,
7075	 => std_logic_vector(to_unsigned(74,8) ,
7076	 => std_logic_vector(to_unsigned(77,8) ,
7077	 => std_logic_vector(to_unsigned(73,8) ,
7078	 => std_logic_vector(to_unsigned(76,8) ,
7079	 => std_logic_vector(to_unsigned(78,8) ,
7080	 => std_logic_vector(to_unsigned(79,8) ,
7081	 => std_logic_vector(to_unsigned(86,8) ,
7082	 => std_logic_vector(to_unsigned(87,8) ,
7083	 => std_logic_vector(to_unsigned(87,8) ,
7084	 => std_logic_vector(to_unsigned(88,8) ,
7085	 => std_logic_vector(to_unsigned(91,8) ,
7086	 => std_logic_vector(to_unsigned(88,8) ,
7087	 => std_logic_vector(to_unsigned(91,8) ,
7088	 => std_logic_vector(to_unsigned(92,8) ,
7089	 => std_logic_vector(to_unsigned(95,8) ,
7090	 => std_logic_vector(to_unsigned(99,8) ,
7091	 => std_logic_vector(to_unsigned(97,8) ,
7092	 => std_logic_vector(to_unsigned(96,8) ,
7093	 => std_logic_vector(to_unsigned(101,8) ,
7094	 => std_logic_vector(to_unsigned(104,8) ,
7095	 => std_logic_vector(to_unsigned(103,8) ,
7096	 => std_logic_vector(to_unsigned(104,8) ,
7097	 => std_logic_vector(to_unsigned(107,8) ,
7098	 => std_logic_vector(to_unsigned(104,8) ,
7099	 => std_logic_vector(to_unsigned(100,8) ,
7100	 => std_logic_vector(to_unsigned(101,8) ,
7101	 => std_logic_vector(to_unsigned(103,8) ,
7102	 => std_logic_vector(to_unsigned(99,8) ,
7103	 => std_logic_vector(to_unsigned(103,8) ,
7104	 => std_logic_vector(to_unsigned(105,8) ,
7105	 => std_logic_vector(to_unsigned(105,8) ,
7106	 => std_logic_vector(to_unsigned(109,8) ,
7107	 => std_logic_vector(to_unsigned(107,8) ,
7108	 => std_logic_vector(to_unsigned(107,8) ,
7109	 => std_logic_vector(to_unsigned(114,8) ,
7110	 => std_logic_vector(to_unsigned(112,8) ,
7111	 => std_logic_vector(to_unsigned(105,8) ,
7112	 => std_logic_vector(to_unsigned(107,8) ,
7113	 => std_logic_vector(to_unsigned(112,8) ,
7114	 => std_logic_vector(to_unsigned(112,8) ,
7115	 => std_logic_vector(to_unsigned(107,8) ,
7116	 => std_logic_vector(to_unsigned(107,8) ,
7117	 => std_logic_vector(to_unsigned(109,8) ,
7118	 => std_logic_vector(to_unsigned(107,8) ,
7119	 => std_logic_vector(to_unsigned(108,8) ,
7120	 => std_logic_vector(to_unsigned(105,8) ,
7121	 => std_logic_vector(to_unsigned(103,8) ,
7122	 => std_logic_vector(to_unsigned(99,8) ,
7123	 => std_logic_vector(to_unsigned(100,8) ,
7124	 => std_logic_vector(to_unsigned(100,8) ,
7125	 => std_logic_vector(to_unsigned(97,8) ,
7126	 => std_logic_vector(to_unsigned(92,8) ,
7127	 => std_logic_vector(to_unsigned(90,8) ,
7128	 => std_logic_vector(to_unsigned(91,8) ,
7129	 => std_logic_vector(to_unsigned(91,8) ,
7130	 => std_logic_vector(to_unsigned(93,8) ,
7131	 => std_logic_vector(to_unsigned(99,8) ,
7132	 => std_logic_vector(to_unsigned(96,8) ,
7133	 => std_logic_vector(to_unsigned(91,8) ,
7134	 => std_logic_vector(to_unsigned(90,8) ,
7135	 => std_logic_vector(to_unsigned(87,8) ,
7136	 => std_logic_vector(to_unsigned(85,8) ,
7137	 => std_logic_vector(to_unsigned(88,8) ,
7138	 => std_logic_vector(to_unsigned(85,8) ,
7139	 => std_logic_vector(to_unsigned(84,8) ,
7140	 => std_logic_vector(to_unsigned(85,8) ,
7141	 => std_logic_vector(to_unsigned(85,8) ,
7142	 => std_logic_vector(to_unsigned(80,8) ,
7143	 => std_logic_vector(to_unsigned(79,8) ,
7144	 => std_logic_vector(to_unsigned(85,8) ,
7145	 => std_logic_vector(to_unsigned(77,8) ,
7146	 => std_logic_vector(to_unsigned(79,8) ,
7147	 => std_logic_vector(to_unsigned(77,8) ,
7148	 => std_logic_vector(to_unsigned(74,8) ,
7149	 => std_logic_vector(to_unsigned(77,8) ,
7150	 => std_logic_vector(to_unsigned(76,8) ,
7151	 => std_logic_vector(to_unsigned(78,8) ,
7152	 => std_logic_vector(to_unsigned(78,8) ,
7153	 => std_logic_vector(to_unsigned(74,8) ,
7154	 => std_logic_vector(to_unsigned(78,8) ,
7155	 => std_logic_vector(to_unsigned(82,8) ,
7156	 => std_logic_vector(to_unsigned(86,8) ,
7157	 => std_logic_vector(to_unsigned(84,8) ,
7158	 => std_logic_vector(to_unsigned(85,8) ,
7159	 => std_logic_vector(to_unsigned(90,8) ,
7160	 => std_logic_vector(to_unsigned(97,8) ,
7161	 => std_logic_vector(to_unsigned(99,8) ,
7162	 => std_logic_vector(to_unsigned(96,8) ,
7163	 => std_logic_vector(to_unsigned(90,8) ,
7164	 => std_logic_vector(to_unsigned(95,8) ,
7165	 => std_logic_vector(to_unsigned(96,8) ,
7166	 => std_logic_vector(to_unsigned(97,8) ,
7167	 => std_logic_vector(to_unsigned(95,8) ,
7168	 => std_logic_vector(to_unsigned(95,8) ,
7169	 => std_logic_vector(to_unsigned(97,8) ,
7170	 => std_logic_vector(to_unsigned(99,8) ,
7171	 => std_logic_vector(to_unsigned(104,8) ,
7172	 => std_logic_vector(to_unsigned(104,8) ,
7173	 => std_logic_vector(to_unsigned(100,8) ,
7174	 => std_logic_vector(to_unsigned(96,8) ,
7175	 => std_logic_vector(to_unsigned(88,8) ,
7176	 => std_logic_vector(to_unsigned(92,8) ,
7177	 => std_logic_vector(to_unsigned(95,8) ,
7178	 => std_logic_vector(to_unsigned(96,8) ,
7179	 => std_logic_vector(to_unsigned(99,8) ,
7180	 => std_logic_vector(to_unsigned(97,8) ,
7181	 => std_logic_vector(to_unsigned(99,8) ,
7182	 => std_logic_vector(to_unsigned(99,8) ,
7183	 => std_logic_vector(to_unsigned(103,8) ,
7184	 => std_logic_vector(to_unsigned(114,8) ,
7185	 => std_logic_vector(to_unsigned(114,8) ,
7186	 => std_logic_vector(to_unsigned(112,8) ,
7187	 => std_logic_vector(to_unsigned(107,8) ,
7188	 => std_logic_vector(to_unsigned(103,8) ,
7189	 => std_logic_vector(to_unsigned(101,8) ,
7190	 => std_logic_vector(to_unsigned(103,8) ,
7191	 => std_logic_vector(to_unsigned(107,8) ,
7192	 => std_logic_vector(to_unsigned(105,8) ,
7193	 => std_logic_vector(to_unsigned(104,8) ,
7194	 => std_logic_vector(to_unsigned(104,8) ,
7195	 => std_logic_vector(to_unsigned(105,8) ,
7196	 => std_logic_vector(to_unsigned(105,8) ,
7197	 => std_logic_vector(to_unsigned(104,8) ,
7198	 => std_logic_vector(to_unsigned(104,8) ,
7199	 => std_logic_vector(to_unsigned(107,8) ,
7200	 => std_logic_vector(to_unsigned(108,8) ,
7201	 => std_logic_vector(to_unsigned(109,8) ,
7202	 => std_logic_vector(to_unsigned(100,8) ,
7203	 => std_logic_vector(to_unsigned(95,8) ,
7204	 => std_logic_vector(to_unsigned(93,8) ,
7205	 => std_logic_vector(to_unsigned(95,8) ,
7206	 => std_logic_vector(to_unsigned(95,8) ,
7207	 => std_logic_vector(to_unsigned(96,8) ,
7208	 => std_logic_vector(to_unsigned(95,8) ,
7209	 => std_logic_vector(to_unsigned(93,8) ,
7210	 => std_logic_vector(to_unsigned(92,8) ,
7211	 => std_logic_vector(to_unsigned(91,8) ,
7212	 => std_logic_vector(to_unsigned(88,8) ,
7213	 => std_logic_vector(to_unsigned(91,8) ,
7214	 => std_logic_vector(to_unsigned(87,8) ,
7215	 => std_logic_vector(to_unsigned(84,8) ,
7216	 => std_logic_vector(to_unsigned(84,8) ,
7217	 => std_logic_vector(to_unsigned(90,8) ,
7218	 => std_logic_vector(to_unsigned(88,8) ,
7219	 => std_logic_vector(to_unsigned(87,8) ,
7220	 => std_logic_vector(to_unsigned(86,8) ,
7221	 => std_logic_vector(to_unsigned(78,8) ,
7222	 => std_logic_vector(to_unsigned(73,8) ,
7223	 => std_logic_vector(to_unsigned(70,8) ,
7224	 => std_logic_vector(to_unsigned(66,8) ,
7225	 => std_logic_vector(to_unsigned(68,8) ,
7226	 => std_logic_vector(to_unsigned(71,8) ,
7227	 => std_logic_vector(to_unsigned(72,8) ,
7228	 => std_logic_vector(to_unsigned(76,8) ,
7229	 => std_logic_vector(to_unsigned(77,8) ,
7230	 => std_logic_vector(to_unsigned(69,8) ,
7231	 => std_logic_vector(to_unsigned(67,8) ,
7232	 => std_logic_vector(to_unsigned(69,8) ,
7233	 => std_logic_vector(to_unsigned(67,8) ,
7234	 => std_logic_vector(to_unsigned(68,8) ,
7235	 => std_logic_vector(to_unsigned(59,8) ,
7236	 => std_logic_vector(to_unsigned(57,8) ,
7237	 => std_logic_vector(to_unsigned(66,8) ,
7238	 => std_logic_vector(to_unsigned(57,8) ,
7239	 => std_logic_vector(to_unsigned(64,8) ,
7240	 => std_logic_vector(to_unsigned(73,8) ,
7241	 => std_logic_vector(to_unsigned(68,8) ,
7242	 => std_logic_vector(to_unsigned(64,8) ,
7243	 => std_logic_vector(to_unsigned(73,8) ,
7244	 => std_logic_vector(to_unsigned(77,8) ,
7245	 => std_logic_vector(to_unsigned(69,8) ,
7246	 => std_logic_vector(to_unsigned(65,8) ,
7247	 => std_logic_vector(to_unsigned(62,8) ,
7248	 => std_logic_vector(to_unsigned(69,8) ,
7249	 => std_logic_vector(to_unsigned(72,8) ,
7250	 => std_logic_vector(to_unsigned(64,8) ,
7251	 => std_logic_vector(to_unsigned(67,8) ,
7252	 => std_logic_vector(to_unsigned(64,8) ,
7253	 => std_logic_vector(to_unsigned(64,8) ,
7254	 => std_logic_vector(to_unsigned(70,8) ,
7255	 => std_logic_vector(to_unsigned(68,8) ,
7256	 => std_logic_vector(to_unsigned(68,8) ,
7257	 => std_logic_vector(to_unsigned(68,8) ,
7258	 => std_logic_vector(to_unsigned(71,8) ,
7259	 => std_logic_vector(to_unsigned(66,8) ,
7260	 => std_logic_vector(to_unsigned(65,8) ,
7261	 => std_logic_vector(to_unsigned(68,8) ,
7262	 => std_logic_vector(to_unsigned(68,8) ,
7263	 => std_logic_vector(to_unsigned(65,8) ,
7264	 => std_logic_vector(to_unsigned(66,8) ,
7265	 => std_logic_vector(to_unsigned(69,8) ,
7266	 => std_logic_vector(to_unsigned(69,8) ,
7267	 => std_logic_vector(to_unsigned(67,8) ,
7268	 => std_logic_vector(to_unsigned(62,8) ,
7269	 => std_logic_vector(to_unsigned(59,8) ,
7270	 => std_logic_vector(to_unsigned(58,8) ,
7271	 => std_logic_vector(to_unsigned(55,8) ,
7272	 => std_logic_vector(to_unsigned(56,8) ,
7273	 => std_logic_vector(to_unsigned(60,8) ,
7274	 => std_logic_vector(to_unsigned(63,8) ,
7275	 => std_logic_vector(to_unsigned(65,8) ,
7276	 => std_logic_vector(to_unsigned(62,8) ,
7277	 => std_logic_vector(to_unsigned(60,8) ,
7278	 => std_logic_vector(to_unsigned(57,8) ,
7279	 => std_logic_vector(to_unsigned(63,8) ,
7280	 => std_logic_vector(to_unsigned(36,8) ,
7281	 => std_logic_vector(to_unsigned(1,8) ,
7282	 => std_logic_vector(to_unsigned(0,8) ,
7283	 => std_logic_vector(to_unsigned(1,8) ,
7284	 => std_logic_vector(to_unsigned(35,8) ,
7285	 => std_logic_vector(to_unsigned(87,8) ,
7286	 => std_logic_vector(to_unsigned(72,8) ,
7287	 => std_logic_vector(to_unsigned(71,8) ,
7288	 => std_logic_vector(to_unsigned(76,8) ,
7289	 => std_logic_vector(to_unsigned(81,8) ,
7290	 => std_logic_vector(to_unsigned(80,8) ,
7291	 => std_logic_vector(to_unsigned(84,8) ,
7292	 => std_logic_vector(to_unsigned(85,8) ,
7293	 => std_logic_vector(to_unsigned(81,8) ,
7294	 => std_logic_vector(to_unsigned(79,8) ,
7295	 => std_logic_vector(to_unsigned(73,8) ,
7296	 => std_logic_vector(to_unsigned(70,8) ,
7297	 => std_logic_vector(to_unsigned(74,8) ,
7298	 => std_logic_vector(to_unsigned(80,8) ,
7299	 => std_logic_vector(to_unsigned(99,8) ,
7300	 => std_logic_vector(to_unsigned(100,8) ,
7301	 => std_logic_vector(to_unsigned(96,8) ,
7302	 => std_logic_vector(to_unsigned(96,8) ,
7303	 => std_logic_vector(to_unsigned(90,8) ,
7304	 => std_logic_vector(to_unsigned(79,8) ,
7305	 => std_logic_vector(to_unsigned(86,8) ,
7306	 => std_logic_vector(to_unsigned(92,8) ,
7307	 => std_logic_vector(to_unsigned(90,8) ,
7308	 => std_logic_vector(to_unsigned(85,8) ,
7309	 => std_logic_vector(to_unsigned(85,8) ,
7310	 => std_logic_vector(to_unsigned(90,8) ,
7311	 => std_logic_vector(to_unsigned(85,8) ,
7312	 => std_logic_vector(to_unsigned(90,8) ,
7313	 => std_logic_vector(to_unsigned(93,8) ,
7314	 => std_logic_vector(to_unsigned(91,8) ,
7315	 => std_logic_vector(to_unsigned(96,8) ,
7316	 => std_logic_vector(to_unsigned(93,8) ,
7317	 => std_logic_vector(to_unsigned(97,8) ,
7318	 => std_logic_vector(to_unsigned(100,8) ,
7319	 => std_logic_vector(to_unsigned(100,8) ,
7320	 => std_logic_vector(to_unsigned(99,8) ,
7321	 => std_logic_vector(to_unsigned(109,8) ,
7322	 => std_logic_vector(to_unsigned(111,8) ,
7323	 => std_logic_vector(to_unsigned(114,8) ,
7324	 => std_logic_vector(to_unsigned(104,8) ,
7325	 => std_logic_vector(to_unsigned(101,8) ,
7326	 => std_logic_vector(to_unsigned(105,8) ,
7327	 => std_logic_vector(to_unsigned(105,8) ,
7328	 => std_logic_vector(to_unsigned(111,8) ,
7329	 => std_logic_vector(to_unsigned(121,8) ,
7330	 => std_logic_vector(to_unsigned(118,8) ,
7331	 => std_logic_vector(to_unsigned(116,8) ,
7332	 => std_logic_vector(to_unsigned(125,8) ,
7333	 => std_logic_vector(to_unsigned(122,8) ,
7334	 => std_logic_vector(to_unsigned(128,8) ,
7335	 => std_logic_vector(to_unsigned(139,8) ,
7336	 => std_logic_vector(to_unsigned(136,8) ,
7337	 => std_logic_vector(to_unsigned(131,8) ,
7338	 => std_logic_vector(to_unsigned(136,8) ,
7339	 => std_logic_vector(to_unsigned(141,8) ,
7340	 => std_logic_vector(to_unsigned(136,8) ,
7341	 => std_logic_vector(to_unsigned(141,8) ,
7342	 => std_logic_vector(to_unsigned(144,8) ,
7343	 => std_logic_vector(to_unsigned(149,8) ,
7344	 => std_logic_vector(to_unsigned(149,8) ,
7345	 => std_logic_vector(to_unsigned(149,8) ,
7346	 => std_logic_vector(to_unsigned(142,8) ,
7347	 => std_logic_vector(to_unsigned(144,8) ,
7348	 => std_logic_vector(to_unsigned(146,8) ,
7349	 => std_logic_vector(to_unsigned(146,8) ,
7350	 => std_logic_vector(to_unsigned(147,8) ,
7351	 => std_logic_vector(to_unsigned(144,8) ,
7352	 => std_logic_vector(to_unsigned(144,8) ,
7353	 => std_logic_vector(to_unsigned(152,8) ,
7354	 => std_logic_vector(to_unsigned(151,8) ,
7355	 => std_logic_vector(to_unsigned(144,8) ,
7356	 => std_logic_vector(to_unsigned(149,8) ,
7357	 => std_logic_vector(to_unsigned(154,8) ,
7358	 => std_logic_vector(to_unsigned(152,8) ,
7359	 => std_logic_vector(to_unsigned(147,8) ,
7360	 => std_logic_vector(to_unsigned(149,8) ,
7361	 => std_logic_vector(to_unsigned(79,8) ,
7362	 => std_logic_vector(to_unsigned(80,8) ,
7363	 => std_logic_vector(to_unsigned(81,8) ,
7364	 => std_logic_vector(to_unsigned(81,8) ,
7365	 => std_logic_vector(to_unsigned(77,8) ,
7366	 => std_logic_vector(to_unsigned(74,8) ,
7367	 => std_logic_vector(to_unsigned(70,8) ,
7368	 => std_logic_vector(to_unsigned(79,8) ,
7369	 => std_logic_vector(to_unsigned(86,8) ,
7370	 => std_logic_vector(to_unsigned(79,8) ,
7371	 => std_logic_vector(to_unsigned(66,8) ,
7372	 => std_logic_vector(to_unsigned(71,8) ,
7373	 => std_logic_vector(to_unsigned(78,8) ,
7374	 => std_logic_vector(to_unsigned(73,8) ,
7375	 => std_logic_vector(to_unsigned(72,8) ,
7376	 => std_logic_vector(to_unsigned(74,8) ,
7377	 => std_logic_vector(to_unsigned(69,8) ,
7378	 => std_logic_vector(to_unsigned(72,8) ,
7379	 => std_logic_vector(to_unsigned(73,8) ,
7380	 => std_logic_vector(to_unsigned(71,8) ,
7381	 => std_logic_vector(to_unsigned(72,8) ,
7382	 => std_logic_vector(to_unsigned(77,8) ,
7383	 => std_logic_vector(to_unsigned(67,8) ,
7384	 => std_logic_vector(to_unsigned(67,8) ,
7385	 => std_logic_vector(to_unsigned(73,8) ,
7386	 => std_logic_vector(to_unsigned(74,8) ,
7387	 => std_logic_vector(to_unsigned(76,8) ,
7388	 => std_logic_vector(to_unsigned(71,8) ,
7389	 => std_logic_vector(to_unsigned(71,8) ,
7390	 => std_logic_vector(to_unsigned(71,8) ,
7391	 => std_logic_vector(to_unsigned(76,8) ,
7392	 => std_logic_vector(to_unsigned(76,8) ,
7393	 => std_logic_vector(to_unsigned(72,8) ,
7394	 => std_logic_vector(to_unsigned(76,8) ,
7395	 => std_logic_vector(to_unsigned(78,8) ,
7396	 => std_logic_vector(to_unsigned(77,8) ,
7397	 => std_logic_vector(to_unsigned(77,8) ,
7398	 => std_logic_vector(to_unsigned(78,8) ,
7399	 => std_logic_vector(to_unsigned(79,8) ,
7400	 => std_logic_vector(to_unsigned(79,8) ,
7401	 => std_logic_vector(to_unsigned(80,8) ,
7402	 => std_logic_vector(to_unsigned(81,8) ,
7403	 => std_logic_vector(to_unsigned(90,8) ,
7404	 => std_logic_vector(to_unsigned(92,8) ,
7405	 => std_logic_vector(to_unsigned(93,8) ,
7406	 => std_logic_vector(to_unsigned(90,8) ,
7407	 => std_logic_vector(to_unsigned(92,8) ,
7408	 => std_logic_vector(to_unsigned(97,8) ,
7409	 => std_logic_vector(to_unsigned(97,8) ,
7410	 => std_logic_vector(to_unsigned(95,8) ,
7411	 => std_logic_vector(to_unsigned(96,8) ,
7412	 => std_logic_vector(to_unsigned(96,8) ,
7413	 => std_logic_vector(to_unsigned(99,8) ,
7414	 => std_logic_vector(to_unsigned(100,8) ,
7415	 => std_logic_vector(to_unsigned(95,8) ,
7416	 => std_logic_vector(to_unsigned(99,8) ,
7417	 => std_logic_vector(to_unsigned(105,8) ,
7418	 => std_logic_vector(to_unsigned(103,8) ,
7419	 => std_logic_vector(to_unsigned(96,8) ,
7420	 => std_logic_vector(to_unsigned(97,8) ,
7421	 => std_logic_vector(to_unsigned(103,8) ,
7422	 => std_logic_vector(to_unsigned(99,8) ,
7423	 => std_logic_vector(to_unsigned(99,8) ,
7424	 => std_logic_vector(to_unsigned(107,8) ,
7425	 => std_logic_vector(to_unsigned(100,8) ,
7426	 => std_logic_vector(to_unsigned(104,8) ,
7427	 => std_logic_vector(to_unsigned(111,8) ,
7428	 => std_logic_vector(to_unsigned(111,8) ,
7429	 => std_logic_vector(to_unsigned(112,8) ,
7430	 => std_logic_vector(to_unsigned(109,8) ,
7431	 => std_logic_vector(to_unsigned(107,8) ,
7432	 => std_logic_vector(to_unsigned(112,8) ,
7433	 => std_logic_vector(to_unsigned(114,8) ,
7434	 => std_logic_vector(to_unsigned(112,8) ,
7435	 => std_logic_vector(to_unsigned(103,8) ,
7436	 => std_logic_vector(to_unsigned(105,8) ,
7437	 => std_logic_vector(to_unsigned(107,8) ,
7438	 => std_logic_vector(to_unsigned(103,8) ,
7439	 => std_logic_vector(to_unsigned(107,8) ,
7440	 => std_logic_vector(to_unsigned(104,8) ,
7441	 => std_logic_vector(to_unsigned(100,8) ,
7442	 => std_logic_vector(to_unsigned(100,8) ,
7443	 => std_logic_vector(to_unsigned(103,8) ,
7444	 => std_logic_vector(to_unsigned(103,8) ,
7445	 => std_logic_vector(to_unsigned(101,8) ,
7446	 => std_logic_vector(to_unsigned(97,8) ,
7447	 => std_logic_vector(to_unsigned(100,8) ,
7448	 => std_logic_vector(to_unsigned(103,8) ,
7449	 => std_logic_vector(to_unsigned(97,8) ,
7450	 => std_logic_vector(to_unsigned(93,8) ,
7451	 => std_logic_vector(to_unsigned(100,8) ,
7452	 => std_logic_vector(to_unsigned(103,8) ,
7453	 => std_logic_vector(to_unsigned(96,8) ,
7454	 => std_logic_vector(to_unsigned(93,8) ,
7455	 => std_logic_vector(to_unsigned(96,8) ,
7456	 => std_logic_vector(to_unsigned(93,8) ,
7457	 => std_logic_vector(to_unsigned(92,8) ,
7458	 => std_logic_vector(to_unsigned(92,8) ,
7459	 => std_logic_vector(to_unsigned(88,8) ,
7460	 => std_logic_vector(to_unsigned(86,8) ,
7461	 => std_logic_vector(to_unsigned(84,8) ,
7462	 => std_logic_vector(to_unsigned(78,8) ,
7463	 => std_logic_vector(to_unsigned(82,8) ,
7464	 => std_logic_vector(to_unsigned(81,8) ,
7465	 => std_logic_vector(to_unsigned(76,8) ,
7466	 => std_logic_vector(to_unsigned(79,8) ,
7467	 => std_logic_vector(to_unsigned(74,8) ,
7468	 => std_logic_vector(to_unsigned(78,8) ,
7469	 => std_logic_vector(to_unsigned(76,8) ,
7470	 => std_logic_vector(to_unsigned(76,8) ,
7471	 => std_logic_vector(to_unsigned(77,8) ,
7472	 => std_logic_vector(to_unsigned(77,8) ,
7473	 => std_logic_vector(to_unsigned(76,8) ,
7474	 => std_logic_vector(to_unsigned(80,8) ,
7475	 => std_logic_vector(to_unsigned(85,8) ,
7476	 => std_logic_vector(to_unsigned(90,8) ,
7477	 => std_logic_vector(to_unsigned(90,8) ,
7478	 => std_logic_vector(to_unsigned(87,8) ,
7479	 => std_logic_vector(to_unsigned(91,8) ,
7480	 => std_logic_vector(to_unsigned(97,8) ,
7481	 => std_logic_vector(to_unsigned(95,8) ,
7482	 => std_logic_vector(to_unsigned(97,8) ,
7483	 => std_logic_vector(to_unsigned(97,8) ,
7484	 => std_logic_vector(to_unsigned(95,8) ,
7485	 => std_logic_vector(to_unsigned(93,8) ,
7486	 => std_logic_vector(to_unsigned(95,8) ,
7487	 => std_logic_vector(to_unsigned(95,8) ,
7488	 => std_logic_vector(to_unsigned(95,8) ,
7489	 => std_logic_vector(to_unsigned(99,8) ,
7490	 => std_logic_vector(to_unsigned(104,8) ,
7491	 => std_logic_vector(to_unsigned(107,8) ,
7492	 => std_logic_vector(to_unsigned(104,8) ,
7493	 => std_logic_vector(to_unsigned(104,8) ,
7494	 => std_logic_vector(to_unsigned(103,8) ,
7495	 => std_logic_vector(to_unsigned(99,8) ,
7496	 => std_logic_vector(to_unsigned(96,8) ,
7497	 => std_logic_vector(to_unsigned(99,8) ,
7498	 => std_logic_vector(to_unsigned(99,8) ,
7499	 => std_logic_vector(to_unsigned(101,8) ,
7500	 => std_logic_vector(to_unsigned(100,8) ,
7501	 => std_logic_vector(to_unsigned(105,8) ,
7502	 => std_logic_vector(to_unsigned(112,8) ,
7503	 => std_logic_vector(to_unsigned(114,8) ,
7504	 => std_logic_vector(to_unsigned(116,8) ,
7505	 => std_logic_vector(to_unsigned(119,8) ,
7506	 => std_logic_vector(to_unsigned(119,8) ,
7507	 => std_logic_vector(to_unsigned(115,8) ,
7508	 => std_logic_vector(to_unsigned(105,8) ,
7509	 => std_logic_vector(to_unsigned(105,8) ,
7510	 => std_logic_vector(to_unsigned(111,8) ,
7511	 => std_logic_vector(to_unsigned(109,8) ,
7512	 => std_logic_vector(to_unsigned(101,8) ,
7513	 => std_logic_vector(to_unsigned(105,8) ,
7514	 => std_logic_vector(to_unsigned(109,8) ,
7515	 => std_logic_vector(to_unsigned(107,8) ,
7516	 => std_logic_vector(to_unsigned(104,8) ,
7517	 => std_logic_vector(to_unsigned(107,8) ,
7518	 => std_logic_vector(to_unsigned(111,8) ,
7519	 => std_logic_vector(to_unsigned(109,8) ,
7520	 => std_logic_vector(to_unsigned(104,8) ,
7521	 => std_logic_vector(to_unsigned(105,8) ,
7522	 => std_logic_vector(to_unsigned(101,8) ,
7523	 => std_logic_vector(to_unsigned(99,8) ,
7524	 => std_logic_vector(to_unsigned(96,8) ,
7525	 => std_logic_vector(to_unsigned(95,8) ,
7526	 => std_logic_vector(to_unsigned(97,8) ,
7527	 => std_logic_vector(to_unsigned(99,8) ,
7528	 => std_logic_vector(to_unsigned(99,8) ,
7529	 => std_logic_vector(to_unsigned(96,8) ,
7530	 => std_logic_vector(to_unsigned(96,8) ,
7531	 => std_logic_vector(to_unsigned(90,8) ,
7532	 => std_logic_vector(to_unsigned(78,8) ,
7533	 => std_logic_vector(to_unsigned(77,8) ,
7534	 => std_logic_vector(to_unsigned(72,8) ,
7535	 => std_logic_vector(to_unsigned(73,8) ,
7536	 => std_logic_vector(to_unsigned(81,8) ,
7537	 => std_logic_vector(to_unsigned(87,8) ,
7538	 => std_logic_vector(to_unsigned(81,8) ,
7539	 => std_logic_vector(to_unsigned(67,8) ,
7540	 => std_logic_vector(to_unsigned(66,8) ,
7541	 => std_logic_vector(to_unsigned(68,8) ,
7542	 => std_logic_vector(to_unsigned(74,8) ,
7543	 => std_logic_vector(to_unsigned(71,8) ,
7544	 => std_logic_vector(to_unsigned(60,8) ,
7545	 => std_logic_vector(to_unsigned(64,8) ,
7546	 => std_logic_vector(to_unsigned(68,8) ,
7547	 => std_logic_vector(to_unsigned(74,8) ,
7548	 => std_logic_vector(to_unsigned(81,8) ,
7549	 => std_logic_vector(to_unsigned(76,8) ,
7550	 => std_logic_vector(to_unsigned(72,8) ,
7551	 => std_logic_vector(to_unsigned(69,8) ,
7552	 => std_logic_vector(to_unsigned(66,8) ,
7553	 => std_logic_vector(to_unsigned(67,8) ,
7554	 => std_logic_vector(to_unsigned(68,8) ,
7555	 => std_logic_vector(to_unsigned(65,8) ,
7556	 => std_logic_vector(to_unsigned(63,8) ,
7557	 => std_logic_vector(to_unsigned(63,8) ,
7558	 => std_logic_vector(to_unsigned(70,8) ,
7559	 => std_logic_vector(to_unsigned(66,8) ,
7560	 => std_logic_vector(to_unsigned(66,8) ,
7561	 => std_logic_vector(to_unsigned(71,8) ,
7562	 => std_logic_vector(to_unsigned(66,8) ,
7563	 => std_logic_vector(to_unsigned(67,8) ,
7564	 => std_logic_vector(to_unsigned(68,8) ,
7565	 => std_logic_vector(to_unsigned(63,8) ,
7566	 => std_logic_vector(to_unsigned(68,8) ,
7567	 => std_logic_vector(to_unsigned(69,8) ,
7568	 => std_logic_vector(to_unsigned(73,8) ,
7569	 => std_logic_vector(to_unsigned(71,8) ,
7570	 => std_logic_vector(to_unsigned(64,8) ,
7571	 => std_logic_vector(to_unsigned(70,8) ,
7572	 => std_logic_vector(to_unsigned(68,8) ,
7573	 => std_logic_vector(to_unsigned(64,8) ,
7574	 => std_logic_vector(to_unsigned(64,8) ,
7575	 => std_logic_vector(to_unsigned(63,8) ,
7576	 => std_logic_vector(to_unsigned(70,8) ,
7577	 => std_logic_vector(to_unsigned(67,8) ,
7578	 => std_logic_vector(to_unsigned(68,8) ,
7579	 => std_logic_vector(to_unsigned(74,8) ,
7580	 => std_logic_vector(to_unsigned(68,8) ,
7581	 => std_logic_vector(to_unsigned(66,8) ,
7582	 => std_logic_vector(to_unsigned(68,8) ,
7583	 => std_logic_vector(to_unsigned(71,8) ,
7584	 => std_logic_vector(to_unsigned(72,8) ,
7585	 => std_logic_vector(to_unsigned(70,8) ,
7586	 => std_logic_vector(to_unsigned(64,8) ,
7587	 => std_logic_vector(to_unsigned(65,8) ,
7588	 => std_logic_vector(to_unsigned(63,8) ,
7589	 => std_logic_vector(to_unsigned(63,8) ,
7590	 => std_logic_vector(to_unsigned(59,8) ,
7591	 => std_logic_vector(to_unsigned(53,8) ,
7592	 => std_logic_vector(to_unsigned(56,8) ,
7593	 => std_logic_vector(to_unsigned(59,8) ,
7594	 => std_logic_vector(to_unsigned(56,8) ,
7595	 => std_logic_vector(to_unsigned(55,8) ,
7596	 => std_logic_vector(to_unsigned(56,8) ,
7597	 => std_logic_vector(to_unsigned(53,8) ,
7598	 => std_logic_vector(to_unsigned(52,8) ,
7599	 => std_logic_vector(to_unsigned(51,8) ,
7600	 => std_logic_vector(to_unsigned(39,8) ,
7601	 => std_logic_vector(to_unsigned(3,8) ,
7602	 => std_logic_vector(to_unsigned(0,8) ,
7603	 => std_logic_vector(to_unsigned(0,8) ,
7604	 => std_logic_vector(to_unsigned(18,8) ,
7605	 => std_logic_vector(to_unsigned(79,8) ,
7606	 => std_logic_vector(to_unsigned(65,8) ,
7607	 => std_logic_vector(to_unsigned(71,8) ,
7608	 => std_logic_vector(to_unsigned(81,8) ,
7609	 => std_logic_vector(to_unsigned(79,8) ,
7610	 => std_logic_vector(to_unsigned(78,8) ,
7611	 => std_logic_vector(to_unsigned(85,8) ,
7612	 => std_logic_vector(to_unsigned(90,8) ,
7613	 => std_logic_vector(to_unsigned(82,8) ,
7614	 => std_logic_vector(to_unsigned(73,8) ,
7615	 => std_logic_vector(to_unsigned(69,8) ,
7616	 => std_logic_vector(to_unsigned(69,8) ,
7617	 => std_logic_vector(to_unsigned(73,8) ,
7618	 => std_logic_vector(to_unsigned(80,8) ,
7619	 => std_logic_vector(to_unsigned(95,8) ,
7620	 => std_logic_vector(to_unsigned(99,8) ,
7621	 => std_logic_vector(to_unsigned(99,8) ,
7622	 => std_logic_vector(to_unsigned(101,8) ,
7623	 => std_logic_vector(to_unsigned(96,8) ,
7624	 => std_logic_vector(to_unsigned(85,8) ,
7625	 => std_logic_vector(to_unsigned(82,8) ,
7626	 => std_logic_vector(to_unsigned(82,8) ,
7627	 => std_logic_vector(to_unsigned(93,8) ,
7628	 => std_logic_vector(to_unsigned(101,8) ,
7629	 => std_logic_vector(to_unsigned(87,8) ,
7630	 => std_logic_vector(to_unsigned(87,8) ,
7631	 => std_logic_vector(to_unsigned(82,8) ,
7632	 => std_logic_vector(to_unsigned(92,8) ,
7633	 => std_logic_vector(to_unsigned(97,8) ,
7634	 => std_logic_vector(to_unsigned(91,8) ,
7635	 => std_logic_vector(to_unsigned(97,8) ,
7636	 => std_logic_vector(to_unsigned(95,8) ,
7637	 => std_logic_vector(to_unsigned(99,8) ,
7638	 => std_logic_vector(to_unsigned(103,8) ,
7639	 => std_logic_vector(to_unsigned(107,8) ,
7640	 => std_logic_vector(to_unsigned(99,8) ,
7641	 => std_logic_vector(to_unsigned(104,8) ,
7642	 => std_logic_vector(to_unsigned(105,8) ,
7643	 => std_logic_vector(to_unsigned(108,8) ,
7644	 => std_logic_vector(to_unsigned(107,8) ,
7645	 => std_logic_vector(to_unsigned(109,8) ,
7646	 => std_logic_vector(to_unsigned(114,8) ,
7647	 => std_logic_vector(to_unsigned(108,8) ,
7648	 => std_logic_vector(to_unsigned(107,8) ,
7649	 => std_logic_vector(to_unsigned(111,8) ,
7650	 => std_logic_vector(to_unsigned(114,8) ,
7651	 => std_logic_vector(to_unsigned(111,8) ,
7652	 => std_logic_vector(to_unsigned(111,8) ,
7653	 => std_logic_vector(to_unsigned(115,8) ,
7654	 => std_logic_vector(to_unsigned(118,8) ,
7655	 => std_logic_vector(to_unsigned(128,8) ,
7656	 => std_logic_vector(to_unsigned(131,8) ,
7657	 => std_logic_vector(to_unsigned(133,8) ,
7658	 => std_logic_vector(to_unsigned(134,8) ,
7659	 => std_logic_vector(to_unsigned(138,8) ,
7660	 => std_logic_vector(to_unsigned(136,8) ,
7661	 => std_logic_vector(to_unsigned(141,8) ,
7662	 => std_logic_vector(to_unsigned(141,8) ,
7663	 => std_logic_vector(to_unsigned(141,8) ,
7664	 => std_logic_vector(to_unsigned(146,8) ,
7665	 => std_logic_vector(to_unsigned(151,8) ,
7666	 => std_logic_vector(to_unsigned(144,8) ,
7667	 => std_logic_vector(to_unsigned(142,8) ,
7668	 => std_logic_vector(to_unsigned(146,8) ,
7669	 => std_logic_vector(to_unsigned(144,8) ,
7670	 => std_logic_vector(to_unsigned(146,8) ,
7671	 => std_logic_vector(to_unsigned(149,8) ,
7672	 => std_logic_vector(to_unsigned(142,8) ,
7673	 => std_logic_vector(to_unsigned(147,8) ,
7674	 => std_logic_vector(to_unsigned(154,8) ,
7675	 => std_logic_vector(to_unsigned(147,8) ,
7676	 => std_logic_vector(to_unsigned(151,8) ,
7677	 => std_logic_vector(to_unsigned(156,8) ,
7678	 => std_logic_vector(to_unsigned(151,8) ,
7679	 => std_logic_vector(to_unsigned(149,8) ,
7680	 => std_logic_vector(to_unsigned(151,8) ,
7681	 => std_logic_vector(to_unsigned(84,8) ,
7682	 => std_logic_vector(to_unsigned(77,8) ,
7683	 => std_logic_vector(to_unsigned(77,8) ,
7684	 => std_logic_vector(to_unsigned(78,8) ,
7685	 => std_logic_vector(to_unsigned(73,8) ,
7686	 => std_logic_vector(to_unsigned(73,8) ,
7687	 => std_logic_vector(to_unsigned(77,8) ,
7688	 => std_logic_vector(to_unsigned(73,8) ,
7689	 => std_logic_vector(to_unsigned(72,8) ,
7690	 => std_logic_vector(to_unsigned(77,8) ,
7691	 => std_logic_vector(to_unsigned(73,8) ,
7692	 => std_logic_vector(to_unsigned(73,8) ,
7693	 => std_logic_vector(to_unsigned(74,8) ,
7694	 => std_logic_vector(to_unsigned(70,8) ,
7695	 => std_logic_vector(to_unsigned(70,8) ,
7696	 => std_logic_vector(to_unsigned(69,8) ,
7697	 => std_logic_vector(to_unsigned(69,8) ,
7698	 => std_logic_vector(to_unsigned(76,8) ,
7699	 => std_logic_vector(to_unsigned(74,8) ,
7700	 => std_logic_vector(to_unsigned(72,8) ,
7701	 => std_logic_vector(to_unsigned(70,8) ,
7702	 => std_logic_vector(to_unsigned(70,8) ,
7703	 => std_logic_vector(to_unsigned(69,8) ,
7704	 => std_logic_vector(to_unsigned(72,8) ,
7705	 => std_logic_vector(to_unsigned(77,8) ,
7706	 => std_logic_vector(to_unsigned(77,8) ,
7707	 => std_logic_vector(to_unsigned(74,8) ,
7708	 => std_logic_vector(to_unsigned(72,8) ,
7709	 => std_logic_vector(to_unsigned(76,8) ,
7710	 => std_logic_vector(to_unsigned(77,8) ,
7711	 => std_logic_vector(to_unsigned(73,8) ,
7712	 => std_logic_vector(to_unsigned(76,8) ,
7713	 => std_logic_vector(to_unsigned(74,8) ,
7714	 => std_logic_vector(to_unsigned(74,8) ,
7715	 => std_logic_vector(to_unsigned(78,8) ,
7716	 => std_logic_vector(to_unsigned(82,8) ,
7717	 => std_logic_vector(to_unsigned(80,8) ,
7718	 => std_logic_vector(to_unsigned(84,8) ,
7719	 => std_logic_vector(to_unsigned(82,8) ,
7720	 => std_logic_vector(to_unsigned(80,8) ,
7721	 => std_logic_vector(to_unsigned(81,8) ,
7722	 => std_logic_vector(to_unsigned(82,8) ,
7723	 => std_logic_vector(to_unsigned(86,8) ,
7724	 => std_logic_vector(to_unsigned(85,8) ,
7725	 => std_logic_vector(to_unsigned(91,8) ,
7726	 => std_logic_vector(to_unsigned(97,8) ,
7727	 => std_logic_vector(to_unsigned(99,8) ,
7728	 => std_logic_vector(to_unsigned(96,8) ,
7729	 => std_logic_vector(to_unsigned(97,8) ,
7730	 => std_logic_vector(to_unsigned(99,8) ,
7731	 => std_logic_vector(to_unsigned(100,8) ,
7732	 => std_logic_vector(to_unsigned(100,8) ,
7733	 => std_logic_vector(to_unsigned(99,8) ,
7734	 => std_logic_vector(to_unsigned(95,8) ,
7735	 => std_logic_vector(to_unsigned(92,8) ,
7736	 => std_logic_vector(to_unsigned(97,8) ,
7737	 => std_logic_vector(to_unsigned(104,8) ,
7738	 => std_logic_vector(to_unsigned(107,8) ,
7739	 => std_logic_vector(to_unsigned(100,8) ,
7740	 => std_logic_vector(to_unsigned(93,8) ,
7741	 => std_logic_vector(to_unsigned(101,8) ,
7742	 => std_logic_vector(to_unsigned(100,8) ,
7743	 => std_logic_vector(to_unsigned(100,8) ,
7744	 => std_logic_vector(to_unsigned(109,8) ,
7745	 => std_logic_vector(to_unsigned(103,8) ,
7746	 => std_logic_vector(to_unsigned(103,8) ,
7747	 => std_logic_vector(to_unsigned(112,8) ,
7748	 => std_logic_vector(to_unsigned(114,8) ,
7749	 => std_logic_vector(to_unsigned(114,8) ,
7750	 => std_logic_vector(to_unsigned(112,8) ,
7751	 => std_logic_vector(to_unsigned(116,8) ,
7752	 => std_logic_vector(to_unsigned(118,8) ,
7753	 => std_logic_vector(to_unsigned(115,8) ,
7754	 => std_logic_vector(to_unsigned(114,8) ,
7755	 => std_logic_vector(to_unsigned(112,8) ,
7756	 => std_logic_vector(to_unsigned(109,8) ,
7757	 => std_logic_vector(to_unsigned(109,8) ,
7758	 => std_logic_vector(to_unsigned(105,8) ,
7759	 => std_logic_vector(to_unsigned(109,8) ,
7760	 => std_logic_vector(to_unsigned(111,8) ,
7761	 => std_logic_vector(to_unsigned(108,8) ,
7762	 => std_logic_vector(to_unsigned(101,8) ,
7763	 => std_logic_vector(to_unsigned(104,8) ,
7764	 => std_logic_vector(to_unsigned(105,8) ,
7765	 => std_logic_vector(to_unsigned(105,8) ,
7766	 => std_logic_vector(to_unsigned(101,8) ,
7767	 => std_logic_vector(to_unsigned(103,8) ,
7768	 => std_logic_vector(to_unsigned(105,8) ,
7769	 => std_logic_vector(to_unsigned(101,8) ,
7770	 => std_logic_vector(to_unsigned(99,8) ,
7771	 => std_logic_vector(to_unsigned(103,8) ,
7772	 => std_logic_vector(to_unsigned(107,8) ,
7773	 => std_logic_vector(to_unsigned(103,8) ,
7774	 => std_logic_vector(to_unsigned(100,8) ,
7775	 => std_logic_vector(to_unsigned(97,8) ,
7776	 => std_logic_vector(to_unsigned(96,8) ,
7777	 => std_logic_vector(to_unsigned(93,8) ,
7778	 => std_logic_vector(to_unsigned(95,8) ,
7779	 => std_logic_vector(to_unsigned(92,8) ,
7780	 => std_logic_vector(to_unsigned(86,8) ,
7781	 => std_logic_vector(to_unsigned(80,8) ,
7782	 => std_logic_vector(to_unsigned(76,8) ,
7783	 => std_logic_vector(to_unsigned(79,8) ,
7784	 => std_logic_vector(to_unsigned(79,8) ,
7785	 => std_logic_vector(to_unsigned(81,8) ,
7786	 => std_logic_vector(to_unsigned(78,8) ,
7787	 => std_logic_vector(to_unsigned(77,8) ,
7788	 => std_logic_vector(to_unsigned(79,8) ,
7789	 => std_logic_vector(to_unsigned(74,8) ,
7790	 => std_logic_vector(to_unsigned(74,8) ,
7791	 => std_logic_vector(to_unsigned(80,8) ,
7792	 => std_logic_vector(to_unsigned(77,8) ,
7793	 => std_logic_vector(to_unsigned(76,8) ,
7794	 => std_logic_vector(to_unsigned(78,8) ,
7795	 => std_logic_vector(to_unsigned(85,8) ,
7796	 => std_logic_vector(to_unsigned(91,8) ,
7797	 => std_logic_vector(to_unsigned(92,8) ,
7798	 => std_logic_vector(to_unsigned(92,8) ,
7799	 => std_logic_vector(to_unsigned(91,8) ,
7800	 => std_logic_vector(to_unsigned(99,8) ,
7801	 => std_logic_vector(to_unsigned(97,8) ,
7802	 => std_logic_vector(to_unsigned(95,8) ,
7803	 => std_logic_vector(to_unsigned(96,8) ,
7804	 => std_logic_vector(to_unsigned(95,8) ,
7805	 => std_logic_vector(to_unsigned(93,8) ,
7806	 => std_logic_vector(to_unsigned(99,8) ,
7807	 => std_logic_vector(to_unsigned(104,8) ,
7808	 => std_logic_vector(to_unsigned(101,8) ,
7809	 => std_logic_vector(to_unsigned(104,8) ,
7810	 => std_logic_vector(to_unsigned(109,8) ,
7811	 => std_logic_vector(to_unsigned(111,8) ,
7812	 => std_logic_vector(to_unsigned(111,8) ,
7813	 => std_logic_vector(to_unsigned(109,8) ,
7814	 => std_logic_vector(to_unsigned(114,8) ,
7815	 => std_logic_vector(to_unsigned(107,8) ,
7816	 => std_logic_vector(to_unsigned(100,8) ,
7817	 => std_logic_vector(to_unsigned(103,8) ,
7818	 => std_logic_vector(to_unsigned(101,8) ,
7819	 => std_logic_vector(to_unsigned(104,8) ,
7820	 => std_logic_vector(to_unsigned(107,8) ,
7821	 => std_logic_vector(to_unsigned(111,8) ,
7822	 => std_logic_vector(to_unsigned(114,8) ,
7823	 => std_logic_vector(to_unsigned(112,8) ,
7824	 => std_logic_vector(to_unsigned(115,8) ,
7825	 => std_logic_vector(to_unsigned(115,8) ,
7826	 => std_logic_vector(to_unsigned(114,8) ,
7827	 => std_logic_vector(to_unsigned(112,8) ,
7828	 => std_logic_vector(to_unsigned(109,8) ,
7829	 => std_logic_vector(to_unsigned(111,8) ,
7830	 => std_logic_vector(to_unsigned(109,8) ,
7831	 => std_logic_vector(to_unsigned(107,8) ,
7832	 => std_logic_vector(to_unsigned(103,8) ,
7833	 => std_logic_vector(to_unsigned(104,8) ,
7834	 => std_logic_vector(to_unsigned(105,8) ,
7835	 => std_logic_vector(to_unsigned(104,8) ,
7836	 => std_logic_vector(to_unsigned(107,8) ,
7837	 => std_logic_vector(to_unsigned(105,8) ,
7838	 => std_logic_vector(to_unsigned(109,8) ,
7839	 => std_logic_vector(to_unsigned(109,8) ,
7840	 => std_logic_vector(to_unsigned(107,8) ,
7841	 => std_logic_vector(to_unsigned(97,8) ,
7842	 => std_logic_vector(to_unsigned(88,8) ,
7843	 => std_logic_vector(to_unsigned(93,8) ,
7844	 => std_logic_vector(to_unsigned(91,8) ,
7845	 => std_logic_vector(to_unsigned(87,8) ,
7846	 => std_logic_vector(to_unsigned(91,8) ,
7847	 => std_logic_vector(to_unsigned(96,8) ,
7848	 => std_logic_vector(to_unsigned(97,8) ,
7849	 => std_logic_vector(to_unsigned(95,8) ,
7850	 => std_logic_vector(to_unsigned(93,8) ,
7851	 => std_logic_vector(to_unsigned(84,8) ,
7852	 => std_logic_vector(to_unsigned(61,8) ,
7853	 => std_logic_vector(to_unsigned(63,8) ,
7854	 => std_logic_vector(to_unsigned(70,8) ,
7855	 => std_logic_vector(to_unsigned(71,8) ,
7856	 => std_logic_vector(to_unsigned(80,8) ,
7857	 => std_logic_vector(to_unsigned(92,8) ,
7858	 => std_logic_vector(to_unsigned(84,8) ,
7859	 => std_logic_vector(to_unsigned(65,8) ,
7860	 => std_logic_vector(to_unsigned(65,8) ,
7861	 => std_logic_vector(to_unsigned(66,8) ,
7862	 => std_logic_vector(to_unsigned(69,8) ,
7863	 => std_logic_vector(to_unsigned(74,8) ,
7864	 => std_logic_vector(to_unsigned(69,8) ,
7865	 => std_logic_vector(to_unsigned(67,8) ,
7866	 => std_logic_vector(to_unsigned(76,8) ,
7867	 => std_logic_vector(to_unsigned(82,8) ,
7868	 => std_logic_vector(to_unsigned(86,8) ,
7869	 => std_logic_vector(to_unsigned(81,8) ,
7870	 => std_logic_vector(to_unsigned(80,8) ,
7871	 => std_logic_vector(to_unsigned(67,8) ,
7872	 => std_logic_vector(to_unsigned(65,8) ,
7873	 => std_logic_vector(to_unsigned(64,8) ,
7874	 => std_logic_vector(to_unsigned(64,8) ,
7875	 => std_logic_vector(to_unsigned(66,8) ,
7876	 => std_logic_vector(to_unsigned(74,8) ,
7877	 => std_logic_vector(to_unsigned(72,8) ,
7878	 => std_logic_vector(to_unsigned(76,8) ,
7879	 => std_logic_vector(to_unsigned(66,8) ,
7880	 => std_logic_vector(to_unsigned(66,8) ,
7881	 => std_logic_vector(to_unsigned(71,8) ,
7882	 => std_logic_vector(to_unsigned(69,8) ,
7883	 => std_logic_vector(to_unsigned(66,8) ,
7884	 => std_logic_vector(to_unsigned(67,8) ,
7885	 => std_logic_vector(to_unsigned(63,8) ,
7886	 => std_logic_vector(to_unsigned(71,8) ,
7887	 => std_logic_vector(to_unsigned(79,8) ,
7888	 => std_logic_vector(to_unsigned(77,8) ,
7889	 => std_logic_vector(to_unsigned(77,8) ,
7890	 => std_logic_vector(to_unsigned(74,8) ,
7891	 => std_logic_vector(to_unsigned(73,8) ,
7892	 => std_logic_vector(to_unsigned(67,8) ,
7893	 => std_logic_vector(to_unsigned(66,8) ,
7894	 => std_logic_vector(to_unsigned(71,8) ,
7895	 => std_logic_vector(to_unsigned(68,8) ,
7896	 => std_logic_vector(to_unsigned(68,8) ,
7897	 => std_logic_vector(to_unsigned(69,8) ,
7898	 => std_logic_vector(to_unsigned(66,8) ,
7899	 => std_logic_vector(to_unsigned(66,8) ,
7900	 => std_logic_vector(to_unsigned(66,8) ,
7901	 => std_logic_vector(to_unsigned(71,8) ,
7902	 => std_logic_vector(to_unsigned(70,8) ,
7903	 => std_logic_vector(to_unsigned(73,8) ,
7904	 => std_logic_vector(to_unsigned(70,8) ,
7905	 => std_logic_vector(to_unsigned(63,8) ,
7906	 => std_logic_vector(to_unsigned(59,8) ,
7907	 => std_logic_vector(to_unsigned(65,8) ,
7908	 => std_logic_vector(to_unsigned(66,8) ,
7909	 => std_logic_vector(to_unsigned(64,8) ,
7910	 => std_logic_vector(to_unsigned(61,8) ,
7911	 => std_logic_vector(to_unsigned(58,8) ,
7912	 => std_logic_vector(to_unsigned(61,8) ,
7913	 => std_logic_vector(to_unsigned(63,8) ,
7914	 => std_logic_vector(to_unsigned(62,8) ,
7915	 => std_logic_vector(to_unsigned(59,8) ,
7916	 => std_logic_vector(to_unsigned(55,8) ,
7917	 => std_logic_vector(to_unsigned(51,8) ,
7918	 => std_logic_vector(to_unsigned(53,8) ,
7919	 => std_logic_vector(to_unsigned(53,8) ,
7920	 => std_logic_vector(to_unsigned(48,8) ,
7921	 => std_logic_vector(to_unsigned(7,8) ,
7922	 => std_logic_vector(to_unsigned(0,8) ,
7923	 => std_logic_vector(to_unsigned(0,8) ,
7924	 => std_logic_vector(to_unsigned(9,8) ,
7925	 => std_logic_vector(to_unsigned(74,8) ,
7926	 => std_logic_vector(to_unsigned(71,8) ,
7927	 => std_logic_vector(to_unsigned(69,8) ,
7928	 => std_logic_vector(to_unsigned(79,8) ,
7929	 => std_logic_vector(to_unsigned(81,8) ,
7930	 => std_logic_vector(to_unsigned(74,8) ,
7931	 => std_logic_vector(to_unsigned(80,8) ,
7932	 => std_logic_vector(to_unsigned(99,8) ,
7933	 => std_logic_vector(to_unsigned(93,8) ,
7934	 => std_logic_vector(to_unsigned(86,8) ,
7935	 => std_logic_vector(to_unsigned(85,8) ,
7936	 => std_logic_vector(to_unsigned(76,8) ,
7937	 => std_logic_vector(to_unsigned(72,8) ,
7938	 => std_logic_vector(to_unsigned(80,8) ,
7939	 => std_logic_vector(to_unsigned(97,8) ,
7940	 => std_logic_vector(to_unsigned(99,8) ,
7941	 => std_logic_vector(to_unsigned(92,8) ,
7942	 => std_logic_vector(to_unsigned(90,8) ,
7943	 => std_logic_vector(to_unsigned(84,8) ,
7944	 => std_logic_vector(to_unsigned(82,8) ,
7945	 => std_logic_vector(to_unsigned(81,8) ,
7946	 => std_logic_vector(to_unsigned(79,8) ,
7947	 => std_logic_vector(to_unsigned(91,8) ,
7948	 => std_logic_vector(to_unsigned(93,8) ,
7949	 => std_logic_vector(to_unsigned(79,8) ,
7950	 => std_logic_vector(to_unsigned(86,8) ,
7951	 => std_logic_vector(to_unsigned(84,8) ,
7952	 => std_logic_vector(to_unsigned(87,8) ,
7953	 => std_logic_vector(to_unsigned(91,8) ,
7954	 => std_logic_vector(to_unsigned(85,8) ,
7955	 => std_logic_vector(to_unsigned(93,8) ,
7956	 => std_logic_vector(to_unsigned(93,8) ,
7957	 => std_logic_vector(to_unsigned(95,8) ,
7958	 => std_logic_vector(to_unsigned(99,8) ,
7959	 => std_logic_vector(to_unsigned(101,8) ,
7960	 => std_logic_vector(to_unsigned(101,8) ,
7961	 => std_logic_vector(to_unsigned(105,8) ,
7962	 => std_logic_vector(to_unsigned(112,8) ,
7963	 => std_logic_vector(to_unsigned(108,8) ,
7964	 => std_logic_vector(to_unsigned(103,8) ,
7965	 => std_logic_vector(to_unsigned(107,8) ,
7966	 => std_logic_vector(to_unsigned(109,8) ,
7967	 => std_logic_vector(to_unsigned(107,8) ,
7968	 => std_logic_vector(to_unsigned(104,8) ,
7969	 => std_logic_vector(to_unsigned(104,8) ,
7970	 => std_logic_vector(to_unsigned(105,8) ,
7971	 => std_logic_vector(to_unsigned(108,8) ,
7972	 => std_logic_vector(to_unsigned(111,8) ,
7973	 => std_logic_vector(to_unsigned(108,8) ,
7974	 => std_logic_vector(to_unsigned(109,8) ,
7975	 => std_logic_vector(to_unsigned(115,8) ,
7976	 => std_logic_vector(to_unsigned(119,8) ,
7977	 => std_logic_vector(to_unsigned(127,8) ,
7978	 => std_logic_vector(to_unsigned(128,8) ,
7979	 => std_logic_vector(to_unsigned(133,8) ,
7980	 => std_logic_vector(to_unsigned(131,8) ,
7981	 => std_logic_vector(to_unsigned(131,8) ,
7982	 => std_logic_vector(to_unsigned(136,8) ,
7983	 => std_logic_vector(to_unsigned(141,8) ,
7984	 => std_logic_vector(to_unsigned(142,8) ,
7985	 => std_logic_vector(to_unsigned(141,8) ,
7986	 => std_logic_vector(to_unsigned(138,8) ,
7987	 => std_logic_vector(to_unsigned(139,8) ,
7988	 => std_logic_vector(to_unsigned(142,8) ,
7989	 => std_logic_vector(to_unsigned(141,8) ,
7990	 => std_logic_vector(to_unsigned(141,8) ,
7991	 => std_logic_vector(to_unsigned(147,8) ,
7992	 => std_logic_vector(to_unsigned(142,8) ,
7993	 => std_logic_vector(to_unsigned(142,8) ,
7994	 => std_logic_vector(to_unsigned(149,8) ,
7995	 => std_logic_vector(to_unsigned(144,8) ,
7996	 => std_logic_vector(to_unsigned(147,8) ,
7997	 => std_logic_vector(to_unsigned(152,8) ,
7998	 => std_logic_vector(to_unsigned(151,8) ,
7999	 => std_logic_vector(to_unsigned(152,8) ,
8000	 => std_logic_vector(to_unsigned(154,8) ,
8001	 => std_logic_vector(to_unsigned(81,8) ,
8002	 => std_logic_vector(to_unsigned(72,8) ,
8003	 => std_logic_vector(to_unsigned(68,8) ,
8004	 => std_logic_vector(to_unsigned(79,8) ,
8005	 => std_logic_vector(to_unsigned(76,8) ,
8006	 => std_logic_vector(to_unsigned(77,8) ,
8007	 => std_logic_vector(to_unsigned(74,8) ,
8008	 => std_logic_vector(to_unsigned(67,8) ,
8009	 => std_logic_vector(to_unsigned(70,8) ,
8010	 => std_logic_vector(to_unsigned(74,8) ,
8011	 => std_logic_vector(to_unsigned(78,8) ,
8012	 => std_logic_vector(to_unsigned(76,8) ,
8013	 => std_logic_vector(to_unsigned(69,8) ,
8014	 => std_logic_vector(to_unsigned(72,8) ,
8015	 => std_logic_vector(to_unsigned(71,8) ,
8016	 => std_logic_vector(to_unsigned(70,8) ,
8017	 => std_logic_vector(to_unsigned(73,8) ,
8018	 => std_logic_vector(to_unsigned(71,8) ,
8019	 => std_logic_vector(to_unsigned(72,8) ,
8020	 => std_logic_vector(to_unsigned(77,8) ,
8021	 => std_logic_vector(to_unsigned(72,8) ,
8022	 => std_logic_vector(to_unsigned(69,8) ,
8023	 => std_logic_vector(to_unsigned(74,8) ,
8024	 => std_logic_vector(to_unsigned(79,8) ,
8025	 => std_logic_vector(to_unsigned(76,8) ,
8026	 => std_logic_vector(to_unsigned(79,8) ,
8027	 => std_logic_vector(to_unsigned(81,8) ,
8028	 => std_logic_vector(to_unsigned(76,8) ,
8029	 => std_logic_vector(to_unsigned(78,8) ,
8030	 => std_logic_vector(to_unsigned(87,8) ,
8031	 => std_logic_vector(to_unsigned(80,8) ,
8032	 => std_logic_vector(to_unsigned(81,8) ,
8033	 => std_logic_vector(to_unsigned(85,8) ,
8034	 => std_logic_vector(to_unsigned(80,8) ,
8035	 => std_logic_vector(to_unsigned(80,8) ,
8036	 => std_logic_vector(to_unsigned(87,8) ,
8037	 => std_logic_vector(to_unsigned(85,8) ,
8038	 => std_logic_vector(to_unsigned(87,8) ,
8039	 => std_logic_vector(to_unsigned(86,8) ,
8040	 => std_logic_vector(to_unsigned(84,8) ,
8041	 => std_logic_vector(to_unsigned(90,8) ,
8042	 => std_logic_vector(to_unsigned(95,8) ,
8043	 => std_logic_vector(to_unsigned(95,8) ,
8044	 => std_logic_vector(to_unsigned(92,8) ,
8045	 => std_logic_vector(to_unsigned(92,8) ,
8046	 => std_logic_vector(to_unsigned(100,8) ,
8047	 => std_logic_vector(to_unsigned(99,8) ,
8048	 => std_logic_vector(to_unsigned(95,8) ,
8049	 => std_logic_vector(to_unsigned(97,8) ,
8050	 => std_logic_vector(to_unsigned(103,8) ,
8051	 => std_logic_vector(to_unsigned(104,8) ,
8052	 => std_logic_vector(to_unsigned(104,8) ,
8053	 => std_logic_vector(to_unsigned(103,8) ,
8054	 => std_logic_vector(to_unsigned(101,8) ,
8055	 => std_logic_vector(to_unsigned(104,8) ,
8056	 => std_logic_vector(to_unsigned(103,8) ,
8057	 => std_logic_vector(to_unsigned(104,8) ,
8058	 => std_logic_vector(to_unsigned(108,8) ,
8059	 => std_logic_vector(to_unsigned(99,8) ,
8060	 => std_logic_vector(to_unsigned(99,8) ,
8061	 => std_logic_vector(to_unsigned(111,8) ,
8062	 => std_logic_vector(to_unsigned(109,8) ,
8063	 => std_logic_vector(to_unsigned(103,8) ,
8064	 => std_logic_vector(to_unsigned(103,8) ,
8065	 => std_logic_vector(to_unsigned(105,8) ,
8066	 => std_logic_vector(to_unsigned(108,8) ,
8067	 => std_logic_vector(to_unsigned(111,8) ,
8068	 => std_logic_vector(to_unsigned(111,8) ,
8069	 => std_logic_vector(to_unsigned(112,8) ,
8070	 => std_logic_vector(to_unsigned(112,8) ,
8071	 => std_logic_vector(to_unsigned(118,8) ,
8072	 => std_logic_vector(to_unsigned(119,8) ,
8073	 => std_logic_vector(to_unsigned(114,8) ,
8074	 => std_logic_vector(to_unsigned(116,8) ,
8075	 => std_logic_vector(to_unsigned(118,8) ,
8076	 => std_logic_vector(to_unsigned(114,8) ,
8077	 => std_logic_vector(to_unsigned(114,8) ,
8078	 => std_logic_vector(to_unsigned(112,8) ,
8079	 => std_logic_vector(to_unsigned(112,8) ,
8080	 => std_logic_vector(to_unsigned(118,8) ,
8081	 => std_logic_vector(to_unsigned(115,8) ,
8082	 => std_logic_vector(to_unsigned(103,8) ,
8083	 => std_logic_vector(to_unsigned(104,8) ,
8084	 => std_logic_vector(to_unsigned(103,8) ,
8085	 => std_logic_vector(to_unsigned(111,8) ,
8086	 => std_logic_vector(to_unsigned(111,8) ,
8087	 => std_logic_vector(to_unsigned(104,8) ,
8088	 => std_logic_vector(to_unsigned(111,8) ,
8089	 => std_logic_vector(to_unsigned(109,8) ,
8090	 => std_logic_vector(to_unsigned(107,8) ,
8091	 => std_logic_vector(to_unsigned(104,8) ,
8092	 => std_logic_vector(to_unsigned(100,8) ,
8093	 => std_logic_vector(to_unsigned(103,8) ,
8094	 => std_logic_vector(to_unsigned(103,8) ,
8095	 => std_logic_vector(to_unsigned(99,8) ,
8096	 => std_logic_vector(to_unsigned(100,8) ,
8097	 => std_logic_vector(to_unsigned(99,8) ,
8098	 => std_logic_vector(to_unsigned(93,8) ,
8099	 => std_logic_vector(to_unsigned(95,8) ,
8100	 => std_logic_vector(to_unsigned(91,8) ,
8101	 => std_logic_vector(to_unsigned(85,8) ,
8102	 => std_logic_vector(to_unsigned(79,8) ,
8103	 => std_logic_vector(to_unsigned(82,8) ,
8104	 => std_logic_vector(to_unsigned(84,8) ,
8105	 => std_logic_vector(to_unsigned(80,8) ,
8106	 => std_logic_vector(to_unsigned(76,8) ,
8107	 => std_logic_vector(to_unsigned(78,8) ,
8108	 => std_logic_vector(to_unsigned(82,8) ,
8109	 => std_logic_vector(to_unsigned(85,8) ,
8110	 => std_logic_vector(to_unsigned(85,8) ,
8111	 => std_logic_vector(to_unsigned(85,8) ,
8112	 => std_logic_vector(to_unsigned(81,8) ,
8113	 => std_logic_vector(to_unsigned(84,8) ,
8114	 => std_logic_vector(to_unsigned(80,8) ,
8115	 => std_logic_vector(to_unsigned(90,8) ,
8116	 => std_logic_vector(to_unsigned(97,8) ,
8117	 => std_logic_vector(to_unsigned(93,8) ,
8118	 => std_logic_vector(to_unsigned(96,8) ,
8119	 => std_logic_vector(to_unsigned(100,8) ,
8120	 => std_logic_vector(to_unsigned(107,8) ,
8121	 => std_logic_vector(to_unsigned(109,8) ,
8122	 => std_logic_vector(to_unsigned(104,8) ,
8123	 => std_logic_vector(to_unsigned(99,8) ,
8124	 => std_logic_vector(to_unsigned(100,8) ,
8125	 => std_logic_vector(to_unsigned(105,8) ,
8126	 => std_logic_vector(to_unsigned(109,8) ,
8127	 => std_logic_vector(to_unsigned(114,8) ,
8128	 => std_logic_vector(to_unsigned(115,8) ,
8129	 => std_logic_vector(to_unsigned(109,8) ,
8130	 => std_logic_vector(to_unsigned(109,8) ,
8131	 => std_logic_vector(to_unsigned(115,8) ,
8132	 => std_logic_vector(to_unsigned(116,8) ,
8133	 => std_logic_vector(to_unsigned(111,8) ,
8134	 => std_logic_vector(to_unsigned(114,8) ,
8135	 => std_logic_vector(to_unsigned(109,8) ,
8136	 => std_logic_vector(to_unsigned(103,8) ,
8137	 => std_logic_vector(to_unsigned(105,8) ,
8138	 => std_logic_vector(to_unsigned(107,8) ,
8139	 => std_logic_vector(to_unsigned(111,8) ,
8140	 => std_logic_vector(to_unsigned(118,8) ,
8141	 => std_logic_vector(to_unsigned(119,8) ,
8142	 => std_logic_vector(to_unsigned(116,8) ,
8143	 => std_logic_vector(to_unsigned(116,8) ,
8144	 => std_logic_vector(to_unsigned(119,8) ,
8145	 => std_logic_vector(to_unsigned(115,8) ,
8146	 => std_logic_vector(to_unsigned(118,8) ,
8147	 => std_logic_vector(to_unsigned(111,8) ,
8148	 => std_logic_vector(to_unsigned(107,8) ,
8149	 => std_logic_vector(to_unsigned(112,8) ,
8150	 => std_logic_vector(to_unsigned(112,8) ,
8151	 => std_logic_vector(to_unsigned(109,8) ,
8152	 => std_logic_vector(to_unsigned(109,8) ,
8153	 => std_logic_vector(to_unsigned(107,8) ,
8154	 => std_logic_vector(to_unsigned(111,8) ,
8155	 => std_logic_vector(to_unsigned(108,8) ,
8156	 => std_logic_vector(to_unsigned(107,8) ,
8157	 => std_logic_vector(to_unsigned(111,8) ,
8158	 => std_logic_vector(to_unsigned(109,8) ,
8159	 => std_logic_vector(to_unsigned(107,8) ,
8160	 => std_logic_vector(to_unsigned(108,8) ,
8161	 => std_logic_vector(to_unsigned(99,8) ,
8162	 => std_logic_vector(to_unsigned(87,8) ,
8163	 => std_logic_vector(to_unsigned(88,8) ,
8164	 => std_logic_vector(to_unsigned(90,8) ,
8165	 => std_logic_vector(to_unsigned(85,8) ,
8166	 => std_logic_vector(to_unsigned(91,8) ,
8167	 => std_logic_vector(to_unsigned(91,8) ,
8168	 => std_logic_vector(to_unsigned(87,8) ,
8169	 => std_logic_vector(to_unsigned(92,8) ,
8170	 => std_logic_vector(to_unsigned(88,8) ,
8171	 => std_logic_vector(to_unsigned(76,8) ,
8172	 => std_logic_vector(to_unsigned(60,8) ,
8173	 => std_logic_vector(to_unsigned(60,8) ,
8174	 => std_logic_vector(to_unsigned(71,8) ,
8175	 => std_logic_vector(to_unsigned(73,8) ,
8176	 => std_logic_vector(to_unsigned(81,8) ,
8177	 => std_logic_vector(to_unsigned(87,8) ,
8178	 => std_logic_vector(to_unsigned(80,8) ,
8179	 => std_logic_vector(to_unsigned(80,8) ,
8180	 => std_logic_vector(to_unsigned(84,8) ,
8181	 => std_logic_vector(to_unsigned(76,8) ,
8182	 => std_logic_vector(to_unsigned(85,8) ,
8183	 => std_logic_vector(to_unsigned(85,8) ,
8184	 => std_logic_vector(to_unsigned(80,8) ,
8185	 => std_logic_vector(to_unsigned(80,8) ,
8186	 => std_logic_vector(to_unsigned(84,8) ,
8187	 => std_logic_vector(to_unsigned(82,8) ,
8188	 => std_logic_vector(to_unsigned(78,8) ,
8189	 => std_logic_vector(to_unsigned(78,8) ,
8190	 => std_logic_vector(to_unsigned(78,8) ,
8191	 => std_logic_vector(to_unsigned(73,8) ,
8192	 => std_logic_vector(to_unsigned(67,8) ,
8193	 => std_logic_vector(to_unsigned(65,8) ,
8194	 => std_logic_vector(to_unsigned(67,8) ,
8195	 => std_logic_vector(to_unsigned(69,8) ,
8196	 => std_logic_vector(to_unsigned(72,8) ,
8197	 => std_logic_vector(to_unsigned(77,8) ,
8198	 => std_logic_vector(to_unsigned(74,8) ,
8199	 => std_logic_vector(to_unsigned(74,8) ,
8200	 => std_logic_vector(to_unsigned(68,8) ,
8201	 => std_logic_vector(to_unsigned(66,8) ,
8202	 => std_logic_vector(to_unsigned(73,8) ,
8203	 => std_logic_vector(to_unsigned(70,8) ,
8204	 => std_logic_vector(to_unsigned(68,8) ,
8205	 => std_logic_vector(to_unsigned(77,8) ,
8206	 => std_logic_vector(to_unsigned(82,8) ,
8207	 => std_logic_vector(to_unsigned(85,8) ,
8208	 => std_logic_vector(to_unsigned(92,8) ,
8209	 => std_logic_vector(to_unsigned(84,8) ,
8210	 => std_logic_vector(to_unsigned(82,8) ,
8211	 => std_logic_vector(to_unsigned(84,8) ,
8212	 => std_logic_vector(to_unsigned(70,8) ,
8213	 => std_logic_vector(to_unsigned(69,8) ,
8214	 => std_logic_vector(to_unsigned(74,8) ,
8215	 => std_logic_vector(to_unsigned(70,8) ,
8216	 => std_logic_vector(to_unsigned(69,8) ,
8217	 => std_logic_vector(to_unsigned(74,8) ,
8218	 => std_logic_vector(to_unsigned(71,8) ,
8219	 => std_logic_vector(to_unsigned(68,8) ,
8220	 => std_logic_vector(to_unsigned(73,8) ,
8221	 => std_logic_vector(to_unsigned(78,8) ,
8222	 => std_logic_vector(to_unsigned(73,8) ,
8223	 => std_logic_vector(to_unsigned(74,8) ,
8224	 => std_logic_vector(to_unsigned(73,8) ,
8225	 => std_logic_vector(to_unsigned(63,8) ,
8226	 => std_logic_vector(to_unsigned(63,8) ,
8227	 => std_logic_vector(to_unsigned(69,8) ,
8228	 => std_logic_vector(to_unsigned(65,8) ,
8229	 => std_logic_vector(to_unsigned(59,8) ,
8230	 => std_logic_vector(to_unsigned(63,8) ,
8231	 => std_logic_vector(to_unsigned(62,8) ,
8232	 => std_logic_vector(to_unsigned(73,8) ,
8233	 => std_logic_vector(to_unsigned(79,8) ,
8234	 => std_logic_vector(to_unsigned(84,8) ,
8235	 => std_logic_vector(to_unsigned(74,8) ,
8236	 => std_logic_vector(to_unsigned(57,8) ,
8237	 => std_logic_vector(to_unsigned(55,8) ,
8238	 => std_logic_vector(to_unsigned(56,8) ,
8239	 => std_logic_vector(to_unsigned(53,8) ,
8240	 => std_logic_vector(to_unsigned(51,8) ,
8241	 => std_logic_vector(to_unsigned(13,8) ,
8242	 => std_logic_vector(to_unsigned(0,8) ,
8243	 => std_logic_vector(to_unsigned(0,8) ,
8244	 => std_logic_vector(to_unsigned(3,8) ,
8245	 => std_logic_vector(to_unsigned(61,8) ,
8246	 => std_logic_vector(to_unsigned(81,8) ,
8247	 => std_logic_vector(to_unsigned(69,8) ,
8248	 => std_logic_vector(to_unsigned(74,8) ,
8249	 => std_logic_vector(to_unsigned(76,8) ,
8250	 => std_logic_vector(to_unsigned(77,8) ,
8251	 => std_logic_vector(to_unsigned(91,8) ,
8252	 => std_logic_vector(to_unsigned(101,8) ,
8253	 => std_logic_vector(to_unsigned(96,8) ,
8254	 => std_logic_vector(to_unsigned(96,8) ,
8255	 => std_logic_vector(to_unsigned(95,8) ,
8256	 => std_logic_vector(to_unsigned(82,8) ,
8257	 => std_logic_vector(to_unsigned(84,8) ,
8258	 => std_logic_vector(to_unsigned(85,8) ,
8259	 => std_logic_vector(to_unsigned(82,8) ,
8260	 => std_logic_vector(to_unsigned(84,8) ,
8261	 => std_logic_vector(to_unsigned(82,8) ,
8262	 => std_logic_vector(to_unsigned(85,8) ,
8263	 => std_logic_vector(to_unsigned(70,8) ,
8264	 => std_logic_vector(to_unsigned(79,8) ,
8265	 => std_logic_vector(to_unsigned(82,8) ,
8266	 => std_logic_vector(to_unsigned(77,8) ,
8267	 => std_logic_vector(to_unsigned(77,8) ,
8268	 => std_logic_vector(to_unsigned(76,8) ,
8269	 => std_logic_vector(to_unsigned(79,8) ,
8270	 => std_logic_vector(to_unsigned(84,8) ,
8271	 => std_logic_vector(to_unsigned(84,8) ,
8272	 => std_logic_vector(to_unsigned(85,8) ,
8273	 => std_logic_vector(to_unsigned(87,8) ,
8274	 => std_logic_vector(to_unsigned(82,8) ,
8275	 => std_logic_vector(to_unsigned(84,8) ,
8276	 => std_logic_vector(to_unsigned(82,8) ,
8277	 => std_logic_vector(to_unsigned(88,8) ,
8278	 => std_logic_vector(to_unsigned(95,8) ,
8279	 => std_logic_vector(to_unsigned(95,8) ,
8280	 => std_logic_vector(to_unsigned(100,8) ,
8281	 => std_logic_vector(to_unsigned(100,8) ,
8282	 => std_logic_vector(to_unsigned(108,8) ,
8283	 => std_logic_vector(to_unsigned(104,8) ,
8284	 => std_logic_vector(to_unsigned(93,8) ,
8285	 => std_logic_vector(to_unsigned(101,8) ,
8286	 => std_logic_vector(to_unsigned(101,8) ,
8287	 => std_logic_vector(to_unsigned(100,8) ,
8288	 => std_logic_vector(to_unsigned(97,8) ,
8289	 => std_logic_vector(to_unsigned(99,8) ,
8290	 => std_logic_vector(to_unsigned(108,8) ,
8291	 => std_logic_vector(to_unsigned(114,8) ,
8292	 => std_logic_vector(to_unsigned(119,8) ,
8293	 => std_logic_vector(to_unsigned(116,8) ,
8294	 => std_logic_vector(to_unsigned(111,8) ,
8295	 => std_logic_vector(to_unsigned(111,8) ,
8296	 => std_logic_vector(to_unsigned(114,8) ,
8297	 => std_logic_vector(to_unsigned(116,8) ,
8298	 => std_logic_vector(to_unsigned(124,8) ,
8299	 => std_logic_vector(to_unsigned(127,8) ,
8300	 => std_logic_vector(to_unsigned(125,8) ,
8301	 => std_logic_vector(to_unsigned(121,8) ,
8302	 => std_logic_vector(to_unsigned(125,8) ,
8303	 => std_logic_vector(to_unsigned(133,8) ,
8304	 => std_logic_vector(to_unsigned(136,8) ,
8305	 => std_logic_vector(to_unsigned(141,8) ,
8306	 => std_logic_vector(to_unsigned(141,8) ,
8307	 => std_logic_vector(to_unsigned(139,8) ,
8308	 => std_logic_vector(to_unsigned(142,8) ,
8309	 => std_logic_vector(to_unsigned(147,8) ,
8310	 => std_logic_vector(to_unsigned(147,8) ,
8311	 => std_logic_vector(to_unsigned(146,8) ,
8312	 => std_logic_vector(to_unsigned(146,8) ,
8313	 => std_logic_vector(to_unsigned(149,8) ,
8314	 => std_logic_vector(to_unsigned(149,8) ,
8315	 => std_logic_vector(to_unsigned(147,8) ,
8316	 => std_logic_vector(to_unsigned(151,8) ,
8317	 => std_logic_vector(to_unsigned(152,8) ,
8318	 => std_logic_vector(to_unsigned(152,8) ,
8319	 => std_logic_vector(to_unsigned(152,8) ,
8320	 => std_logic_vector(to_unsigned(152,8) ,
8321	 => std_logic_vector(to_unsigned(86,8) ,
8322	 => std_logic_vector(to_unsigned(80,8) ,
8323	 => std_logic_vector(to_unsigned(73,8) ,
8324	 => std_logic_vector(to_unsigned(73,8) ,
8325	 => std_logic_vector(to_unsigned(77,8) ,
8326	 => std_logic_vector(to_unsigned(77,8) ,
8327	 => std_logic_vector(to_unsigned(72,8) ,
8328	 => std_logic_vector(to_unsigned(69,8) ,
8329	 => std_logic_vector(to_unsigned(72,8) ,
8330	 => std_logic_vector(to_unsigned(77,8) ,
8331	 => std_logic_vector(to_unsigned(79,8) ,
8332	 => std_logic_vector(to_unsigned(77,8) ,
8333	 => std_logic_vector(to_unsigned(73,8) ,
8334	 => std_logic_vector(to_unsigned(73,8) ,
8335	 => std_logic_vector(to_unsigned(70,8) ,
8336	 => std_logic_vector(to_unsigned(76,8) ,
8337	 => std_logic_vector(to_unsigned(81,8) ,
8338	 => std_logic_vector(to_unsigned(76,8) ,
8339	 => std_logic_vector(to_unsigned(73,8) ,
8340	 => std_logic_vector(to_unsigned(79,8) ,
8341	 => std_logic_vector(to_unsigned(80,8) ,
8342	 => std_logic_vector(to_unsigned(78,8) ,
8343	 => std_logic_vector(to_unsigned(81,8) ,
8344	 => std_logic_vector(to_unsigned(85,8) ,
8345	 => std_logic_vector(to_unsigned(81,8) ,
8346	 => std_logic_vector(to_unsigned(82,8) ,
8347	 => std_logic_vector(to_unsigned(86,8) ,
8348	 => std_logic_vector(to_unsigned(84,8) ,
8349	 => std_logic_vector(to_unsigned(79,8) ,
8350	 => std_logic_vector(to_unsigned(84,8) ,
8351	 => std_logic_vector(to_unsigned(84,8) ,
8352	 => std_logic_vector(to_unsigned(85,8) ,
8353	 => std_logic_vector(to_unsigned(87,8) ,
8354	 => std_logic_vector(to_unsigned(84,8) ,
8355	 => std_logic_vector(to_unsigned(82,8) ,
8356	 => std_logic_vector(to_unsigned(81,8) ,
8357	 => std_logic_vector(to_unsigned(85,8) ,
8358	 => std_logic_vector(to_unsigned(86,8) ,
8359	 => std_logic_vector(to_unsigned(85,8) ,
8360	 => std_logic_vector(to_unsigned(85,8) ,
8361	 => std_logic_vector(to_unsigned(87,8) ,
8362	 => std_logic_vector(to_unsigned(92,8) ,
8363	 => std_logic_vector(to_unsigned(99,8) ,
8364	 => std_logic_vector(to_unsigned(99,8) ,
8365	 => std_logic_vector(to_unsigned(95,8) ,
8366	 => std_logic_vector(to_unsigned(95,8) ,
8367	 => std_logic_vector(to_unsigned(93,8) ,
8368	 => std_logic_vector(to_unsigned(95,8) ,
8369	 => std_logic_vector(to_unsigned(101,8) ,
8370	 => std_logic_vector(to_unsigned(105,8) ,
8371	 => std_logic_vector(to_unsigned(101,8) ,
8372	 => std_logic_vector(to_unsigned(101,8) ,
8373	 => std_logic_vector(to_unsigned(100,8) ,
8374	 => std_logic_vector(to_unsigned(97,8) ,
8375	 => std_logic_vector(to_unsigned(107,8) ,
8376	 => std_logic_vector(to_unsigned(112,8) ,
8377	 => std_logic_vector(to_unsigned(107,8) ,
8378	 => std_logic_vector(to_unsigned(108,8) ,
8379	 => std_logic_vector(to_unsigned(100,8) ,
8380	 => std_logic_vector(to_unsigned(100,8) ,
8381	 => std_logic_vector(to_unsigned(112,8) ,
8382	 => std_logic_vector(to_unsigned(109,8) ,
8383	 => std_logic_vector(to_unsigned(107,8) ,
8384	 => std_logic_vector(to_unsigned(109,8) ,
8385	 => std_logic_vector(to_unsigned(107,8) ,
8386	 => std_logic_vector(to_unsigned(116,8) ,
8387	 => std_logic_vector(to_unsigned(119,8) ,
8388	 => std_logic_vector(to_unsigned(112,8) ,
8389	 => std_logic_vector(to_unsigned(116,8) ,
8390	 => std_logic_vector(to_unsigned(115,8) ,
8391	 => std_logic_vector(to_unsigned(118,8) ,
8392	 => std_logic_vector(to_unsigned(118,8) ,
8393	 => std_logic_vector(to_unsigned(116,8) ,
8394	 => std_logic_vector(to_unsigned(119,8) ,
8395	 => std_logic_vector(to_unsigned(115,8) ,
8396	 => std_logic_vector(to_unsigned(114,8) ,
8397	 => std_logic_vector(to_unsigned(114,8) ,
8398	 => std_logic_vector(to_unsigned(112,8) ,
8399	 => std_logic_vector(to_unsigned(111,8) ,
8400	 => std_logic_vector(to_unsigned(115,8) ,
8401	 => std_logic_vector(to_unsigned(114,8) ,
8402	 => std_logic_vector(to_unsigned(109,8) ,
8403	 => std_logic_vector(to_unsigned(109,8) ,
8404	 => std_logic_vector(to_unsigned(107,8) ,
8405	 => std_logic_vector(to_unsigned(114,8) ,
8406	 => std_logic_vector(to_unsigned(112,8) ,
8407	 => std_logic_vector(to_unsigned(103,8) ,
8408	 => std_logic_vector(to_unsigned(108,8) ,
8409	 => std_logic_vector(to_unsigned(104,8) ,
8410	 => std_logic_vector(to_unsigned(104,8) ,
8411	 => std_logic_vector(to_unsigned(105,8) ,
8412	 => std_logic_vector(to_unsigned(103,8) ,
8413	 => std_logic_vector(to_unsigned(101,8) ,
8414	 => std_logic_vector(to_unsigned(99,8) ,
8415	 => std_logic_vector(to_unsigned(103,8) ,
8416	 => std_logic_vector(to_unsigned(104,8) ,
8417	 => std_logic_vector(to_unsigned(99,8) ,
8418	 => std_logic_vector(to_unsigned(95,8) ,
8419	 => std_logic_vector(to_unsigned(92,8) ,
8420	 => std_logic_vector(to_unsigned(93,8) ,
8421	 => std_logic_vector(to_unsigned(90,8) ,
8422	 => std_logic_vector(to_unsigned(84,8) ,
8423	 => std_logic_vector(to_unsigned(82,8) ,
8424	 => std_logic_vector(to_unsigned(84,8) ,
8425	 => std_logic_vector(to_unsigned(81,8) ,
8426	 => std_logic_vector(to_unsigned(79,8) ,
8427	 => std_logic_vector(to_unsigned(82,8) ,
8428	 => std_logic_vector(to_unsigned(87,8) ,
8429	 => std_logic_vector(to_unsigned(88,8) ,
8430	 => std_logic_vector(to_unsigned(85,8) ,
8431	 => std_logic_vector(to_unsigned(86,8) ,
8432	 => std_logic_vector(to_unsigned(90,8) ,
8433	 => std_logic_vector(to_unsigned(92,8) ,
8434	 => std_logic_vector(to_unsigned(91,8) ,
8435	 => std_logic_vector(to_unsigned(91,8) ,
8436	 => std_logic_vector(to_unsigned(92,8) ,
8437	 => std_logic_vector(to_unsigned(100,8) ,
8438	 => std_logic_vector(to_unsigned(107,8) ,
8439	 => std_logic_vector(to_unsigned(108,8) ,
8440	 => std_logic_vector(to_unsigned(108,8) ,
8441	 => std_logic_vector(to_unsigned(107,8) ,
8442	 => std_logic_vector(to_unsigned(111,8) ,
8443	 => std_logic_vector(to_unsigned(108,8) ,
8444	 => std_logic_vector(to_unsigned(103,8) ,
8445	 => std_logic_vector(to_unsigned(107,8) ,
8446	 => std_logic_vector(to_unsigned(115,8) ,
8447	 => std_logic_vector(to_unsigned(114,8) ,
8448	 => std_logic_vector(to_unsigned(119,8) ,
8449	 => std_logic_vector(to_unsigned(119,8) ,
8450	 => std_logic_vector(to_unsigned(118,8) ,
8451	 => std_logic_vector(to_unsigned(114,8) ,
8452	 => std_logic_vector(to_unsigned(114,8) ,
8453	 => std_logic_vector(to_unsigned(118,8) ,
8454	 => std_logic_vector(to_unsigned(115,8) ,
8455	 => std_logic_vector(to_unsigned(111,8) ,
8456	 => std_logic_vector(to_unsigned(118,8) ,
8457	 => std_logic_vector(to_unsigned(114,8) ,
8458	 => std_logic_vector(to_unsigned(111,8) ,
8459	 => std_logic_vector(to_unsigned(122,8) ,
8460	 => std_logic_vector(to_unsigned(125,8) ,
8461	 => std_logic_vector(to_unsigned(121,8) ,
8462	 => std_logic_vector(to_unsigned(119,8) ,
8463	 => std_logic_vector(to_unsigned(112,8) ,
8464	 => std_logic_vector(to_unsigned(119,8) ,
8465	 => std_logic_vector(to_unsigned(122,8) ,
8466	 => std_logic_vector(to_unsigned(122,8) ,
8467	 => std_logic_vector(to_unsigned(116,8) ,
8468	 => std_logic_vector(to_unsigned(112,8) ,
8469	 => std_logic_vector(to_unsigned(114,8) ,
8470	 => std_logic_vector(to_unsigned(112,8) ,
8471	 => std_logic_vector(to_unsigned(108,8) ,
8472	 => std_logic_vector(to_unsigned(111,8) ,
8473	 => std_logic_vector(to_unsigned(111,8) ,
8474	 => std_logic_vector(to_unsigned(115,8) ,
8475	 => std_logic_vector(to_unsigned(109,8) ,
8476	 => std_logic_vector(to_unsigned(104,8) ,
8477	 => std_logic_vector(to_unsigned(108,8) ,
8478	 => std_logic_vector(to_unsigned(100,8) ,
8479	 => std_logic_vector(to_unsigned(104,8) ,
8480	 => std_logic_vector(to_unsigned(105,8) ,
8481	 => std_logic_vector(to_unsigned(103,8) ,
8482	 => std_logic_vector(to_unsigned(93,8) ,
8483	 => std_logic_vector(to_unsigned(97,8) ,
8484	 => std_logic_vector(to_unsigned(97,8) ,
8485	 => std_logic_vector(to_unsigned(87,8) ,
8486	 => std_logic_vector(to_unsigned(91,8) ,
8487	 => std_logic_vector(to_unsigned(90,8) ,
8488	 => std_logic_vector(to_unsigned(88,8) ,
8489	 => std_logic_vector(to_unsigned(84,8) ,
8490	 => std_logic_vector(to_unsigned(74,8) ,
8491	 => std_logic_vector(to_unsigned(73,8) ,
8492	 => std_logic_vector(to_unsigned(70,8) ,
8493	 => std_logic_vector(to_unsigned(65,8) ,
8494	 => std_logic_vector(to_unsigned(78,8) ,
8495	 => std_logic_vector(to_unsigned(74,8) ,
8496	 => std_logic_vector(to_unsigned(76,8) ,
8497	 => std_logic_vector(to_unsigned(78,8) ,
8498	 => std_logic_vector(to_unsigned(74,8) ,
8499	 => std_logic_vector(to_unsigned(84,8) ,
8500	 => std_logic_vector(to_unsigned(84,8) ,
8501	 => std_logic_vector(to_unsigned(72,8) ,
8502	 => std_logic_vector(to_unsigned(76,8) ,
8503	 => std_logic_vector(to_unsigned(78,8) ,
8504	 => std_logic_vector(to_unsigned(78,8) ,
8505	 => std_logic_vector(to_unsigned(80,8) ,
8506	 => std_logic_vector(to_unsigned(74,8) ,
8507	 => std_logic_vector(to_unsigned(76,8) ,
8508	 => std_logic_vector(to_unsigned(74,8) ,
8509	 => std_logic_vector(to_unsigned(74,8) ,
8510	 => std_logic_vector(to_unsigned(72,8) ,
8511	 => std_logic_vector(to_unsigned(72,8) ,
8512	 => std_logic_vector(to_unsigned(63,8) ,
8513	 => std_logic_vector(to_unsigned(70,8) ,
8514	 => std_logic_vector(to_unsigned(79,8) ,
8515	 => std_logic_vector(to_unsigned(79,8) ,
8516	 => std_logic_vector(to_unsigned(77,8) ,
8517	 => std_logic_vector(to_unsigned(72,8) ,
8518	 => std_logic_vector(to_unsigned(63,8) ,
8519	 => std_logic_vector(to_unsigned(73,8) ,
8520	 => std_logic_vector(to_unsigned(61,8) ,
8521	 => std_logic_vector(to_unsigned(62,8) ,
8522	 => std_logic_vector(to_unsigned(74,8) ,
8523	 => std_logic_vector(to_unsigned(79,8) ,
8524	 => std_logic_vector(to_unsigned(78,8) ,
8525	 => std_logic_vector(to_unsigned(78,8) ,
8526	 => std_logic_vector(to_unsigned(79,8) ,
8527	 => std_logic_vector(to_unsigned(79,8) ,
8528	 => std_logic_vector(to_unsigned(87,8) ,
8529	 => std_logic_vector(to_unsigned(85,8) ,
8530	 => std_logic_vector(to_unsigned(87,8) ,
8531	 => std_logic_vector(to_unsigned(85,8) ,
8532	 => std_logic_vector(to_unsigned(73,8) ,
8533	 => std_logic_vector(to_unsigned(69,8) ,
8534	 => std_logic_vector(to_unsigned(68,8) ,
8535	 => std_logic_vector(to_unsigned(68,8) ,
8536	 => std_logic_vector(to_unsigned(73,8) ,
8537	 => std_logic_vector(to_unsigned(76,8) ,
8538	 => std_logic_vector(to_unsigned(73,8) ,
8539	 => std_logic_vector(to_unsigned(76,8) ,
8540	 => std_logic_vector(to_unsigned(74,8) ,
8541	 => std_logic_vector(to_unsigned(76,8) ,
8542	 => std_logic_vector(to_unsigned(70,8) ,
8543	 => std_logic_vector(to_unsigned(62,8) ,
8544	 => std_logic_vector(to_unsigned(62,8) ,
8545	 => std_logic_vector(to_unsigned(59,8) ,
8546	 => std_logic_vector(to_unsigned(59,8) ,
8547	 => std_logic_vector(to_unsigned(64,8) ,
8548	 => std_logic_vector(to_unsigned(62,8) ,
8549	 => std_logic_vector(to_unsigned(58,8) ,
8550	 => std_logic_vector(to_unsigned(59,8) ,
8551	 => std_logic_vector(to_unsigned(58,8) ,
8552	 => std_logic_vector(to_unsigned(68,8) ,
8553	 => std_logic_vector(to_unsigned(74,8) ,
8554	 => std_logic_vector(to_unsigned(77,8) ,
8555	 => std_logic_vector(to_unsigned(64,8) ,
8556	 => std_logic_vector(to_unsigned(63,8) ,
8557	 => std_logic_vector(to_unsigned(60,8) ,
8558	 => std_logic_vector(to_unsigned(56,8) ,
8559	 => std_logic_vector(to_unsigned(51,8) ,
8560	 => std_logic_vector(to_unsigned(52,8) ,
8561	 => std_logic_vector(to_unsigned(20,8) ,
8562	 => std_logic_vector(to_unsigned(1,8) ,
8563	 => std_logic_vector(to_unsigned(0,8) ,
8564	 => std_logic_vector(to_unsigned(2,8) ,
8565	 => std_logic_vector(to_unsigned(52,8) ,
8566	 => std_logic_vector(to_unsigned(74,8) ,
8567	 => std_logic_vector(to_unsigned(69,8) ,
8568	 => std_logic_vector(to_unsigned(77,8) ,
8569	 => std_logic_vector(to_unsigned(76,8) ,
8570	 => std_logic_vector(to_unsigned(96,8) ,
8571	 => std_logic_vector(to_unsigned(109,8) ,
8572	 => std_logic_vector(to_unsigned(96,8) ,
8573	 => std_logic_vector(to_unsigned(92,8) ,
8574	 => std_logic_vector(to_unsigned(91,8) ,
8575	 => std_logic_vector(to_unsigned(87,8) ,
8576	 => std_logic_vector(to_unsigned(87,8) ,
8577	 => std_logic_vector(to_unsigned(91,8) ,
8578	 => std_logic_vector(to_unsigned(93,8) ,
8579	 => std_logic_vector(to_unsigned(79,8) ,
8580	 => std_logic_vector(to_unsigned(81,8) ,
8581	 => std_logic_vector(to_unsigned(90,8) ,
8582	 => std_logic_vector(to_unsigned(87,8) ,
8583	 => std_logic_vector(to_unsigned(87,8) ,
8584	 => std_logic_vector(to_unsigned(86,8) ,
8585	 => std_logic_vector(to_unsigned(85,8) ,
8586	 => std_logic_vector(to_unsigned(80,8) ,
8587	 => std_logic_vector(to_unsigned(77,8) ,
8588	 => std_logic_vector(to_unsigned(81,8) ,
8589	 => std_logic_vector(to_unsigned(86,8) ,
8590	 => std_logic_vector(to_unsigned(77,8) ,
8591	 => std_logic_vector(to_unsigned(81,8) ,
8592	 => std_logic_vector(to_unsigned(84,8) ,
8593	 => std_logic_vector(to_unsigned(91,8) ,
8594	 => std_logic_vector(to_unsigned(85,8) ,
8595	 => std_logic_vector(to_unsigned(81,8) ,
8596	 => std_logic_vector(to_unsigned(86,8) ,
8597	 => std_logic_vector(to_unsigned(90,8) ,
8598	 => std_logic_vector(to_unsigned(91,8) ,
8599	 => std_logic_vector(to_unsigned(93,8) ,
8600	 => std_logic_vector(to_unsigned(99,8) ,
8601	 => std_logic_vector(to_unsigned(97,8) ,
8602	 => std_logic_vector(to_unsigned(101,8) ,
8603	 => std_logic_vector(to_unsigned(100,8) ,
8604	 => std_logic_vector(to_unsigned(99,8) ,
8605	 => std_logic_vector(to_unsigned(105,8) ,
8606	 => std_logic_vector(to_unsigned(104,8) ,
8607	 => std_logic_vector(to_unsigned(104,8) ,
8608	 => std_logic_vector(to_unsigned(100,8) ,
8609	 => std_logic_vector(to_unsigned(100,8) ,
8610	 => std_logic_vector(to_unsigned(105,8) ,
8611	 => std_logic_vector(to_unsigned(118,8) ,
8612	 => std_logic_vector(to_unsigned(115,8) ,
8613	 => std_logic_vector(to_unsigned(108,8) ,
8614	 => std_logic_vector(to_unsigned(103,8) ,
8615	 => std_logic_vector(to_unsigned(111,8) ,
8616	 => std_logic_vector(to_unsigned(116,8) ,
8617	 => std_logic_vector(to_unsigned(111,8) ,
8618	 => std_logic_vector(to_unsigned(121,8) ,
8619	 => std_logic_vector(to_unsigned(128,8) ,
8620	 => std_logic_vector(to_unsigned(128,8) ,
8621	 => std_logic_vector(to_unsigned(125,8) ,
8622	 => std_logic_vector(to_unsigned(124,8) ,
8623	 => std_logic_vector(to_unsigned(130,8) ,
8624	 => std_logic_vector(to_unsigned(133,8) ,
8625	 => std_logic_vector(to_unsigned(138,8) ,
8626	 => std_logic_vector(to_unsigned(142,8) ,
8627	 => std_logic_vector(to_unsigned(144,8) ,
8628	 => std_logic_vector(to_unsigned(146,8) ,
8629	 => std_logic_vector(to_unsigned(149,8) ,
8630	 => std_logic_vector(to_unsigned(151,8) ,
8631	 => std_logic_vector(to_unsigned(147,8) ,
8632	 => std_logic_vector(to_unsigned(149,8) ,
8633	 => std_logic_vector(to_unsigned(152,8) ,
8634	 => std_logic_vector(to_unsigned(151,8) ,
8635	 => std_logic_vector(to_unsigned(151,8) ,
8636	 => std_logic_vector(to_unsigned(151,8) ,
8637	 => std_logic_vector(to_unsigned(146,8) ,
8638	 => std_logic_vector(to_unsigned(147,8) ,
8639	 => std_logic_vector(to_unsigned(152,8) ,
8640	 => std_logic_vector(to_unsigned(152,8) ,
8641	 => std_logic_vector(to_unsigned(81,8) ,
8642	 => std_logic_vector(to_unsigned(82,8) ,
8643	 => std_logic_vector(to_unsigned(78,8) ,
8644	 => std_logic_vector(to_unsigned(69,8) ,
8645	 => std_logic_vector(to_unsigned(72,8) ,
8646	 => std_logic_vector(to_unsigned(72,8) ,
8647	 => std_logic_vector(to_unsigned(72,8) ,
8648	 => std_logic_vector(to_unsigned(73,8) ,
8649	 => std_logic_vector(to_unsigned(71,8) ,
8650	 => std_logic_vector(to_unsigned(72,8) ,
8651	 => std_logic_vector(to_unsigned(74,8) ,
8652	 => std_logic_vector(to_unsigned(79,8) ,
8653	 => std_logic_vector(to_unsigned(80,8) ,
8654	 => std_logic_vector(to_unsigned(78,8) ,
8655	 => std_logic_vector(to_unsigned(77,8) ,
8656	 => std_logic_vector(to_unsigned(80,8) ,
8657	 => std_logic_vector(to_unsigned(80,8) ,
8658	 => std_logic_vector(to_unsigned(79,8) ,
8659	 => std_logic_vector(to_unsigned(82,8) ,
8660	 => std_logic_vector(to_unsigned(79,8) ,
8661	 => std_logic_vector(to_unsigned(81,8) ,
8662	 => std_logic_vector(to_unsigned(91,8) ,
8663	 => std_logic_vector(to_unsigned(86,8) ,
8664	 => std_logic_vector(to_unsigned(84,8) ,
8665	 => std_logic_vector(to_unsigned(86,8) ,
8666	 => std_logic_vector(to_unsigned(86,8) ,
8667	 => std_logic_vector(to_unsigned(87,8) ,
8668	 => std_logic_vector(to_unsigned(88,8) ,
8669	 => std_logic_vector(to_unsigned(84,8) ,
8670	 => std_logic_vector(to_unsigned(78,8) ,
8671	 => std_logic_vector(to_unsigned(79,8) ,
8672	 => std_logic_vector(to_unsigned(82,8) ,
8673	 => std_logic_vector(to_unsigned(80,8) ,
8674	 => std_logic_vector(to_unsigned(81,8) ,
8675	 => std_logic_vector(to_unsigned(82,8) ,
8676	 => std_logic_vector(to_unsigned(79,8) ,
8677	 => std_logic_vector(to_unsigned(84,8) ,
8678	 => std_logic_vector(to_unsigned(84,8) ,
8679	 => std_logic_vector(to_unsigned(84,8) ,
8680	 => std_logic_vector(to_unsigned(86,8) ,
8681	 => std_logic_vector(to_unsigned(88,8) ,
8682	 => std_logic_vector(to_unsigned(95,8) ,
8683	 => std_logic_vector(to_unsigned(93,8) ,
8684	 => std_logic_vector(to_unsigned(92,8) ,
8685	 => std_logic_vector(to_unsigned(96,8) ,
8686	 => std_logic_vector(to_unsigned(95,8) ,
8687	 => std_logic_vector(to_unsigned(93,8) ,
8688	 => std_logic_vector(to_unsigned(97,8) ,
8689	 => std_logic_vector(to_unsigned(107,8) ,
8690	 => std_logic_vector(to_unsigned(108,8) ,
8691	 => std_logic_vector(to_unsigned(105,8) ,
8692	 => std_logic_vector(to_unsigned(109,8) ,
8693	 => std_logic_vector(to_unsigned(108,8) ,
8694	 => std_logic_vector(to_unsigned(100,8) ,
8695	 => std_logic_vector(to_unsigned(101,8) ,
8696	 => std_logic_vector(to_unsigned(107,8) ,
8697	 => std_logic_vector(to_unsigned(104,8) ,
8698	 => std_logic_vector(to_unsigned(109,8) ,
8699	 => std_logic_vector(to_unsigned(105,8) ,
8700	 => std_logic_vector(to_unsigned(104,8) ,
8701	 => std_logic_vector(to_unsigned(112,8) ,
8702	 => std_logic_vector(to_unsigned(114,8) ,
8703	 => std_logic_vector(to_unsigned(112,8) ,
8704	 => std_logic_vector(to_unsigned(111,8) ,
8705	 => std_logic_vector(to_unsigned(118,8) ,
8706	 => std_logic_vector(to_unsigned(124,8) ,
8707	 => std_logic_vector(to_unsigned(124,8) ,
8708	 => std_logic_vector(to_unsigned(122,8) ,
8709	 => std_logic_vector(to_unsigned(121,8) ,
8710	 => std_logic_vector(to_unsigned(116,8) ,
8711	 => std_logic_vector(to_unsigned(119,8) ,
8712	 => std_logic_vector(to_unsigned(115,8) ,
8713	 => std_logic_vector(to_unsigned(114,8) ,
8714	 => std_logic_vector(to_unsigned(121,8) ,
8715	 => std_logic_vector(to_unsigned(119,8) ,
8716	 => std_logic_vector(to_unsigned(114,8) ,
8717	 => std_logic_vector(to_unsigned(116,8) ,
8718	 => std_logic_vector(to_unsigned(119,8) ,
8719	 => std_logic_vector(to_unsigned(115,8) ,
8720	 => std_logic_vector(to_unsigned(118,8) ,
8721	 => std_logic_vector(to_unsigned(116,8) ,
8722	 => std_logic_vector(to_unsigned(118,8) ,
8723	 => std_logic_vector(to_unsigned(114,8) ,
8724	 => std_logic_vector(to_unsigned(109,8) ,
8725	 => std_logic_vector(to_unsigned(112,8) ,
8726	 => std_logic_vector(to_unsigned(108,8) ,
8727	 => std_logic_vector(to_unsigned(103,8) ,
8728	 => std_logic_vector(to_unsigned(105,8) ,
8729	 => std_logic_vector(to_unsigned(105,8) ,
8730	 => std_logic_vector(to_unsigned(112,8) ,
8731	 => std_logic_vector(to_unsigned(116,8) ,
8732	 => std_logic_vector(to_unsigned(114,8) ,
8733	 => std_logic_vector(to_unsigned(114,8) ,
8734	 => std_logic_vector(to_unsigned(108,8) ,
8735	 => std_logic_vector(to_unsigned(103,8) ,
8736	 => std_logic_vector(to_unsigned(101,8) ,
8737	 => std_logic_vector(to_unsigned(101,8) ,
8738	 => std_logic_vector(to_unsigned(103,8) ,
8739	 => std_logic_vector(to_unsigned(99,8) ,
8740	 => std_logic_vector(to_unsigned(92,8) ,
8741	 => std_logic_vector(to_unsigned(92,8) ,
8742	 => std_logic_vector(to_unsigned(90,8) ,
8743	 => std_logic_vector(to_unsigned(88,8) ,
8744	 => std_logic_vector(to_unsigned(91,8) ,
8745	 => std_logic_vector(to_unsigned(92,8) ,
8746	 => std_logic_vector(to_unsigned(91,8) ,
8747	 => std_logic_vector(to_unsigned(90,8) ,
8748	 => std_logic_vector(to_unsigned(87,8) ,
8749	 => std_logic_vector(to_unsigned(88,8) ,
8750	 => std_logic_vector(to_unsigned(90,8) ,
8751	 => std_logic_vector(to_unsigned(93,8) ,
8752	 => std_logic_vector(to_unsigned(96,8) ,
8753	 => std_logic_vector(to_unsigned(92,8) ,
8754	 => std_logic_vector(to_unsigned(96,8) ,
8755	 => std_logic_vector(to_unsigned(95,8) ,
8756	 => std_logic_vector(to_unsigned(92,8) ,
8757	 => std_logic_vector(to_unsigned(99,8) ,
8758	 => std_logic_vector(to_unsigned(105,8) ,
8759	 => std_logic_vector(to_unsigned(103,8) ,
8760	 => std_logic_vector(to_unsigned(103,8) ,
8761	 => std_logic_vector(to_unsigned(104,8) ,
8762	 => std_logic_vector(to_unsigned(104,8) ,
8763	 => std_logic_vector(to_unsigned(108,8) ,
8764	 => std_logic_vector(to_unsigned(103,8) ,
8765	 => std_logic_vector(to_unsigned(95,8) ,
8766	 => std_logic_vector(to_unsigned(104,8) ,
8767	 => std_logic_vector(to_unsigned(115,8) ,
8768	 => std_logic_vector(to_unsigned(118,8) ,
8769	 => std_logic_vector(to_unsigned(115,8) ,
8770	 => std_logic_vector(to_unsigned(121,8) ,
8771	 => std_logic_vector(to_unsigned(122,8) ,
8772	 => std_logic_vector(to_unsigned(116,8) ,
8773	 => std_logic_vector(to_unsigned(114,8) ,
8774	 => std_logic_vector(to_unsigned(114,8) ,
8775	 => std_logic_vector(to_unsigned(111,8) ,
8776	 => std_logic_vector(to_unsigned(112,8) ,
8777	 => std_logic_vector(to_unsigned(111,8) ,
8778	 => std_logic_vector(to_unsigned(116,8) ,
8779	 => std_logic_vector(to_unsigned(114,8) ,
8780	 => std_logic_vector(to_unsigned(112,8) ,
8781	 => std_logic_vector(to_unsigned(121,8) ,
8782	 => std_logic_vector(to_unsigned(122,8) ,
8783	 => std_logic_vector(to_unsigned(105,8) ,
8784	 => std_logic_vector(to_unsigned(109,8) ,
8785	 => std_logic_vector(to_unsigned(112,8) ,
8786	 => std_logic_vector(to_unsigned(103,8) ,
8787	 => std_logic_vector(to_unsigned(108,8) ,
8788	 => std_logic_vector(to_unsigned(114,8) ,
8789	 => std_logic_vector(to_unsigned(104,8) ,
8790	 => std_logic_vector(to_unsigned(91,8) ,
8791	 => std_logic_vector(to_unsigned(91,8) ,
8792	 => std_logic_vector(to_unsigned(107,8) ,
8793	 => std_logic_vector(to_unsigned(107,8) ,
8794	 => std_logic_vector(to_unsigned(99,8) ,
8795	 => std_logic_vector(to_unsigned(96,8) ,
8796	 => std_logic_vector(to_unsigned(88,8) ,
8797	 => std_logic_vector(to_unsigned(91,8) ,
8798	 => std_logic_vector(to_unsigned(96,8) ,
8799	 => std_logic_vector(to_unsigned(101,8) ,
8800	 => std_logic_vector(to_unsigned(109,8) ,
8801	 => std_logic_vector(to_unsigned(104,8) ,
8802	 => std_logic_vector(to_unsigned(100,8) ,
8803	 => std_logic_vector(to_unsigned(93,8) ,
8804	 => std_logic_vector(to_unsigned(91,8) ,
8805	 => std_logic_vector(to_unsigned(86,8) ,
8806	 => std_logic_vector(to_unsigned(80,8) ,
8807	 => std_logic_vector(to_unsigned(87,8) ,
8808	 => std_logic_vector(to_unsigned(96,8) ,
8809	 => std_logic_vector(to_unsigned(81,8) ,
8810	 => std_logic_vector(to_unsigned(69,8) ,
8811	 => std_logic_vector(to_unsigned(74,8) ,
8812	 => std_logic_vector(to_unsigned(76,8) ,
8813	 => std_logic_vector(to_unsigned(72,8) ,
8814	 => std_logic_vector(to_unsigned(78,8) ,
8815	 => std_logic_vector(to_unsigned(71,8) ,
8816	 => std_logic_vector(to_unsigned(72,8) ,
8817	 => std_logic_vector(to_unsigned(68,8) ,
8818	 => std_logic_vector(to_unsigned(76,8) ,
8819	 => std_logic_vector(to_unsigned(79,8) ,
8820	 => std_logic_vector(to_unsigned(74,8) ,
8821	 => std_logic_vector(to_unsigned(77,8) ,
8822	 => std_logic_vector(to_unsigned(72,8) ,
8823	 => std_logic_vector(to_unsigned(78,8) ,
8824	 => std_logic_vector(to_unsigned(67,8) ,
8825	 => std_logic_vector(to_unsigned(66,8) ,
8826	 => std_logic_vector(to_unsigned(69,8) ,
8827	 => std_logic_vector(to_unsigned(70,8) ,
8828	 => std_logic_vector(to_unsigned(72,8) ,
8829	 => std_logic_vector(to_unsigned(69,8) ,
8830	 => std_logic_vector(to_unsigned(67,8) ,
8831	 => std_logic_vector(to_unsigned(60,8) ,
8832	 => std_logic_vector(to_unsigned(66,8) ,
8833	 => std_logic_vector(to_unsigned(77,8) ,
8834	 => std_logic_vector(to_unsigned(76,8) ,
8835	 => std_logic_vector(to_unsigned(81,8) ,
8836	 => std_logic_vector(to_unsigned(84,8) ,
8837	 => std_logic_vector(to_unsigned(80,8) ,
8838	 => std_logic_vector(to_unsigned(63,8) ,
8839	 => std_logic_vector(to_unsigned(72,8) ,
8840	 => std_logic_vector(to_unsigned(71,8) ,
8841	 => std_logic_vector(to_unsigned(65,8) ,
8842	 => std_logic_vector(to_unsigned(64,8) ,
8843	 => std_logic_vector(to_unsigned(82,8) ,
8844	 => std_logic_vector(to_unsigned(85,8) ,
8845	 => std_logic_vector(to_unsigned(81,8) ,
8846	 => std_logic_vector(to_unsigned(80,8) ,
8847	 => std_logic_vector(to_unsigned(74,8) ,
8848	 => std_logic_vector(to_unsigned(80,8) ,
8849	 => std_logic_vector(to_unsigned(80,8) ,
8850	 => std_logic_vector(to_unsigned(87,8) ,
8851	 => std_logic_vector(to_unsigned(87,8) ,
8852	 => std_logic_vector(to_unsigned(79,8) ,
8853	 => std_logic_vector(to_unsigned(73,8) ,
8854	 => std_logic_vector(to_unsigned(67,8) ,
8855	 => std_logic_vector(to_unsigned(70,8) ,
8856	 => std_logic_vector(to_unsigned(78,8) ,
8857	 => std_logic_vector(to_unsigned(77,8) ,
8858	 => std_logic_vector(to_unsigned(79,8) ,
8859	 => std_logic_vector(to_unsigned(73,8) ,
8860	 => std_logic_vector(to_unsigned(64,8) ,
8861	 => std_logic_vector(to_unsigned(85,8) ,
8862	 => std_logic_vector(to_unsigned(73,8) ,
8863	 => std_logic_vector(to_unsigned(66,8) ,
8864	 => std_logic_vector(to_unsigned(67,8) ,
8865	 => std_logic_vector(to_unsigned(63,8) ,
8866	 => std_logic_vector(to_unsigned(66,8) ,
8867	 => std_logic_vector(to_unsigned(67,8) ,
8868	 => std_logic_vector(to_unsigned(66,8) ,
8869	 => std_logic_vector(to_unsigned(62,8) ,
8870	 => std_logic_vector(to_unsigned(63,8) ,
8871	 => std_logic_vector(to_unsigned(68,8) ,
8872	 => std_logic_vector(to_unsigned(60,8) ,
8873	 => std_logic_vector(to_unsigned(62,8) ,
8874	 => std_logic_vector(to_unsigned(53,8) ,
8875	 => std_logic_vector(to_unsigned(45,8) ,
8876	 => std_logic_vector(to_unsigned(64,8) ,
8877	 => std_logic_vector(to_unsigned(65,8) ,
8878	 => std_logic_vector(to_unsigned(54,8) ,
8879	 => std_logic_vector(to_unsigned(56,8) ,
8880	 => std_logic_vector(to_unsigned(66,8) ,
8881	 => std_logic_vector(to_unsigned(38,8) ,
8882	 => std_logic_vector(to_unsigned(2,8) ,
8883	 => std_logic_vector(to_unsigned(0,8) ,
8884	 => std_logic_vector(to_unsigned(1,8) ,
8885	 => std_logic_vector(to_unsigned(41,8) ,
8886	 => std_logic_vector(to_unsigned(82,8) ,
8887	 => std_logic_vector(to_unsigned(73,8) ,
8888	 => std_logic_vector(to_unsigned(85,8) ,
8889	 => std_logic_vector(to_unsigned(87,8) ,
8890	 => std_logic_vector(to_unsigned(93,8) ,
8891	 => std_logic_vector(to_unsigned(91,8) ,
8892	 => std_logic_vector(to_unsigned(95,8) ,
8893	 => std_logic_vector(to_unsigned(105,8) ,
8894	 => std_logic_vector(to_unsigned(97,8) ,
8895	 => std_logic_vector(to_unsigned(92,8) ,
8896	 => std_logic_vector(to_unsigned(87,8) ,
8897	 => std_logic_vector(to_unsigned(85,8) ,
8898	 => std_logic_vector(to_unsigned(86,8) ,
8899	 => std_logic_vector(to_unsigned(84,8) ,
8900	 => std_logic_vector(to_unsigned(90,8) ,
8901	 => std_logic_vector(to_unsigned(90,8) ,
8902	 => std_logic_vector(to_unsigned(92,8) ,
8903	 => std_logic_vector(to_unsigned(101,8) ,
8904	 => std_logic_vector(to_unsigned(86,8) ,
8905	 => std_logic_vector(to_unsigned(86,8) ,
8906	 => std_logic_vector(to_unsigned(90,8) ,
8907	 => std_logic_vector(to_unsigned(91,8) ,
8908	 => std_logic_vector(to_unsigned(93,8) ,
8909	 => std_logic_vector(to_unsigned(85,8) ,
8910	 => std_logic_vector(to_unsigned(80,8) ,
8911	 => std_logic_vector(to_unsigned(90,8) ,
8912	 => std_logic_vector(to_unsigned(86,8) ,
8913	 => std_logic_vector(to_unsigned(92,8) ,
8914	 => std_logic_vector(to_unsigned(91,8) ,
8915	 => std_logic_vector(to_unsigned(85,8) ,
8916	 => std_logic_vector(to_unsigned(92,8) ,
8917	 => std_logic_vector(to_unsigned(95,8) ,
8918	 => std_logic_vector(to_unsigned(100,8) ,
8919	 => std_logic_vector(to_unsigned(99,8) ,
8920	 => std_logic_vector(to_unsigned(101,8) ,
8921	 => std_logic_vector(to_unsigned(100,8) ,
8922	 => std_logic_vector(to_unsigned(104,8) ,
8923	 => std_logic_vector(to_unsigned(100,8) ,
8924	 => std_logic_vector(to_unsigned(101,8) ,
8925	 => std_logic_vector(to_unsigned(105,8) ,
8926	 => std_logic_vector(to_unsigned(105,8) ,
8927	 => std_logic_vector(to_unsigned(109,8) ,
8928	 => std_logic_vector(to_unsigned(104,8) ,
8929	 => std_logic_vector(to_unsigned(108,8) ,
8930	 => std_logic_vector(to_unsigned(115,8) ,
8931	 => std_logic_vector(to_unsigned(114,8) ,
8932	 => std_logic_vector(to_unsigned(116,8) ,
8933	 => std_logic_vector(to_unsigned(115,8) ,
8934	 => std_logic_vector(to_unsigned(105,8) ,
8935	 => std_logic_vector(to_unsigned(108,8) ,
8936	 => std_logic_vector(to_unsigned(118,8) ,
8937	 => std_logic_vector(to_unsigned(114,8) ,
8938	 => std_logic_vector(to_unsigned(116,8) ,
8939	 => std_logic_vector(to_unsigned(128,8) ,
8940	 => std_logic_vector(to_unsigned(130,8) ,
8941	 => std_logic_vector(to_unsigned(128,8) ,
8942	 => std_logic_vector(to_unsigned(134,8) ,
8943	 => std_logic_vector(to_unsigned(142,8) ,
8944	 => std_logic_vector(to_unsigned(138,8) ,
8945	 => std_logic_vector(to_unsigned(138,8) ,
8946	 => std_logic_vector(to_unsigned(144,8) ,
8947	 => std_logic_vector(to_unsigned(146,8) ,
8948	 => std_logic_vector(to_unsigned(146,8) ,
8949	 => std_logic_vector(to_unsigned(144,8) ,
8950	 => std_logic_vector(to_unsigned(146,8) ,
8951	 => std_logic_vector(to_unsigned(149,8) ,
8952	 => std_logic_vector(to_unsigned(147,8) ,
8953	 => std_logic_vector(to_unsigned(151,8) ,
8954	 => std_logic_vector(to_unsigned(151,8) ,
8955	 => std_logic_vector(to_unsigned(154,8) ,
8956	 => std_logic_vector(to_unsigned(149,8) ,
8957	 => std_logic_vector(to_unsigned(141,8) ,
8958	 => std_logic_vector(to_unsigned(146,8) ,
8959	 => std_logic_vector(to_unsigned(149,8) ,
8960	 => std_logic_vector(to_unsigned(147,8) ,
8961	 => std_logic_vector(to_unsigned(76,8) ,
8962	 => std_logic_vector(to_unsigned(73,8) ,
8963	 => std_logic_vector(to_unsigned(77,8) ,
8964	 => std_logic_vector(to_unsigned(72,8) ,
8965	 => std_logic_vector(to_unsigned(77,8) ,
8966	 => std_logic_vector(to_unsigned(73,8) ,
8967	 => std_logic_vector(to_unsigned(77,8) ,
8968	 => std_logic_vector(to_unsigned(80,8) ,
8969	 => std_logic_vector(to_unsigned(78,8) ,
8970	 => std_logic_vector(to_unsigned(79,8) ,
8971	 => std_logic_vector(to_unsigned(80,8) ,
8972	 => std_logic_vector(to_unsigned(81,8) ,
8973	 => std_logic_vector(to_unsigned(82,8) ,
8974	 => std_logic_vector(to_unsigned(85,8) ,
8975	 => std_logic_vector(to_unsigned(86,8) ,
8976	 => std_logic_vector(to_unsigned(86,8) ,
8977	 => std_logic_vector(to_unsigned(84,8) ,
8978	 => std_logic_vector(to_unsigned(80,8) ,
8979	 => std_logic_vector(to_unsigned(82,8) ,
8980	 => std_logic_vector(to_unsigned(81,8) ,
8981	 => std_logic_vector(to_unsigned(85,8) ,
8982	 => std_logic_vector(to_unsigned(90,8) ,
8983	 => std_logic_vector(to_unsigned(85,8) ,
8984	 => std_logic_vector(to_unsigned(84,8) ,
8985	 => std_logic_vector(to_unsigned(82,8) ,
8986	 => std_logic_vector(to_unsigned(86,8) ,
8987	 => std_logic_vector(to_unsigned(87,8) ,
8988	 => std_logic_vector(to_unsigned(79,8) ,
8989	 => std_logic_vector(to_unsigned(85,8) ,
8990	 => std_logic_vector(to_unsigned(80,8) ,
8991	 => std_logic_vector(to_unsigned(80,8) ,
8992	 => std_logic_vector(to_unsigned(84,8) ,
8993	 => std_logic_vector(to_unsigned(81,8) ,
8994	 => std_logic_vector(to_unsigned(84,8) ,
8995	 => std_logic_vector(to_unsigned(86,8) ,
8996	 => std_logic_vector(to_unsigned(81,8) ,
8997	 => std_logic_vector(to_unsigned(82,8) ,
8998	 => std_logic_vector(to_unsigned(85,8) ,
8999	 => std_logic_vector(to_unsigned(86,8) ,
9000	 => std_logic_vector(to_unsigned(88,8) ,
9001	 => std_logic_vector(to_unsigned(87,8) ,
9002	 => std_logic_vector(to_unsigned(92,8) ,
9003	 => std_logic_vector(to_unsigned(93,8) ,
9004	 => std_logic_vector(to_unsigned(91,8) ,
9005	 => std_logic_vector(to_unsigned(95,8) ,
9006	 => std_logic_vector(to_unsigned(97,8) ,
9007	 => std_logic_vector(to_unsigned(100,8) ,
9008	 => std_logic_vector(to_unsigned(100,8) ,
9009	 => std_logic_vector(to_unsigned(104,8) ,
9010	 => std_logic_vector(to_unsigned(101,8) ,
9011	 => std_logic_vector(to_unsigned(99,8) ,
9012	 => std_logic_vector(to_unsigned(105,8) ,
9013	 => std_logic_vector(to_unsigned(111,8) ,
9014	 => std_logic_vector(to_unsigned(104,8) ,
9015	 => std_logic_vector(to_unsigned(101,8) ,
9016	 => std_logic_vector(to_unsigned(96,8) ,
9017	 => std_logic_vector(to_unsigned(99,8) ,
9018	 => std_logic_vector(to_unsigned(104,8) ,
9019	 => std_logic_vector(to_unsigned(107,8) ,
9020	 => std_logic_vector(to_unsigned(108,8) ,
9021	 => std_logic_vector(to_unsigned(116,8) ,
9022	 => std_logic_vector(to_unsigned(118,8) ,
9023	 => std_logic_vector(to_unsigned(119,8) ,
9024	 => std_logic_vector(to_unsigned(115,8) ,
9025	 => std_logic_vector(to_unsigned(122,8) ,
9026	 => std_logic_vector(to_unsigned(122,8) ,
9027	 => std_logic_vector(to_unsigned(121,8) ,
9028	 => std_logic_vector(to_unsigned(125,8) ,
9029	 => std_logic_vector(to_unsigned(128,8) ,
9030	 => std_logic_vector(to_unsigned(118,8) ,
9031	 => std_logic_vector(to_unsigned(115,8) ,
9032	 => std_logic_vector(to_unsigned(118,8) ,
9033	 => std_logic_vector(to_unsigned(119,8) ,
9034	 => std_logic_vector(to_unsigned(119,8) ,
9035	 => std_logic_vector(to_unsigned(116,8) ,
9036	 => std_logic_vector(to_unsigned(114,8) ,
9037	 => std_logic_vector(to_unsigned(121,8) ,
9038	 => std_logic_vector(to_unsigned(127,8) ,
9039	 => std_logic_vector(to_unsigned(124,8) ,
9040	 => std_logic_vector(to_unsigned(124,8) ,
9041	 => std_logic_vector(to_unsigned(119,8) ,
9042	 => std_logic_vector(to_unsigned(122,8) ,
9043	 => std_logic_vector(to_unsigned(121,8) ,
9044	 => std_logic_vector(to_unsigned(118,8) ,
9045	 => std_logic_vector(to_unsigned(119,8) ,
9046	 => std_logic_vector(to_unsigned(114,8) ,
9047	 => std_logic_vector(to_unsigned(112,8) ,
9048	 => std_logic_vector(to_unsigned(109,8) ,
9049	 => std_logic_vector(to_unsigned(114,8) ,
9050	 => std_logic_vector(to_unsigned(122,8) ,
9051	 => std_logic_vector(to_unsigned(118,8) ,
9052	 => std_logic_vector(to_unsigned(112,8) ,
9053	 => std_logic_vector(to_unsigned(121,8) ,
9054	 => std_logic_vector(to_unsigned(119,8) ,
9055	 => std_logic_vector(to_unsigned(116,8) ,
9056	 => std_logic_vector(to_unsigned(109,8) ,
9057	 => std_logic_vector(to_unsigned(104,8) ,
9058	 => std_logic_vector(to_unsigned(109,8) ,
9059	 => std_logic_vector(to_unsigned(101,8) ,
9060	 => std_logic_vector(to_unsigned(99,8) ,
9061	 => std_logic_vector(to_unsigned(101,8) ,
9062	 => std_logic_vector(to_unsigned(101,8) ,
9063	 => std_logic_vector(to_unsigned(96,8) ,
9064	 => std_logic_vector(to_unsigned(96,8) ,
9065	 => std_logic_vector(to_unsigned(101,8) ,
9066	 => std_logic_vector(to_unsigned(100,8) ,
9067	 => std_logic_vector(to_unsigned(95,8) ,
9068	 => std_logic_vector(to_unsigned(90,8) ,
9069	 => std_logic_vector(to_unsigned(91,8) ,
9070	 => std_logic_vector(to_unsigned(95,8) ,
9071	 => std_logic_vector(to_unsigned(95,8) ,
9072	 => std_logic_vector(to_unsigned(97,8) ,
9073	 => std_logic_vector(to_unsigned(95,8) ,
9074	 => std_logic_vector(to_unsigned(97,8) ,
9075	 => std_logic_vector(to_unsigned(103,8) ,
9076	 => std_logic_vector(to_unsigned(101,8) ,
9077	 => std_logic_vector(to_unsigned(99,8) ,
9078	 => std_logic_vector(to_unsigned(103,8) ,
9079	 => std_logic_vector(to_unsigned(108,8) ,
9080	 => std_logic_vector(to_unsigned(104,8) ,
9081	 => std_logic_vector(to_unsigned(99,8) ,
9082	 => std_logic_vector(to_unsigned(96,8) ,
9083	 => std_logic_vector(to_unsigned(95,8) ,
9084	 => std_logic_vector(to_unsigned(96,8) ,
9085	 => std_logic_vector(to_unsigned(93,8) ,
9086	 => std_logic_vector(to_unsigned(91,8) ,
9087	 => std_logic_vector(to_unsigned(103,8) ,
9088	 => std_logic_vector(to_unsigned(109,8) ,
9089	 => std_logic_vector(to_unsigned(107,8) ,
9090	 => std_logic_vector(to_unsigned(109,8) ,
9091	 => std_logic_vector(to_unsigned(122,8) ,
9092	 => std_logic_vector(to_unsigned(121,8) ,
9093	 => std_logic_vector(to_unsigned(112,8) ,
9094	 => std_logic_vector(to_unsigned(109,8) ,
9095	 => std_logic_vector(to_unsigned(103,8) ,
9096	 => std_logic_vector(to_unsigned(100,8) ,
9097	 => std_logic_vector(to_unsigned(103,8) ,
9098	 => std_logic_vector(to_unsigned(105,8) ,
9099	 => std_logic_vector(to_unsigned(105,8) ,
9100	 => std_logic_vector(to_unsigned(105,8) ,
9101	 => std_logic_vector(to_unsigned(112,8) ,
9102	 => std_logic_vector(to_unsigned(118,8) ,
9103	 => std_logic_vector(to_unsigned(114,8) ,
9104	 => std_logic_vector(to_unsigned(108,8) ,
9105	 => std_logic_vector(to_unsigned(99,8) ,
9106	 => std_logic_vector(to_unsigned(93,8) ,
9107	 => std_logic_vector(to_unsigned(95,8) ,
9108	 => std_logic_vector(to_unsigned(92,8) ,
9109	 => std_logic_vector(to_unsigned(88,8) ,
9110	 => std_logic_vector(to_unsigned(86,8) ,
9111	 => std_logic_vector(to_unsigned(84,8) ,
9112	 => std_logic_vector(to_unsigned(95,8) ,
9113	 => std_logic_vector(to_unsigned(96,8) ,
9114	 => std_logic_vector(to_unsigned(93,8) ,
9115	 => std_logic_vector(to_unsigned(92,8) ,
9116	 => std_logic_vector(to_unsigned(85,8) ,
9117	 => std_logic_vector(to_unsigned(86,8) ,
9118	 => std_logic_vector(to_unsigned(91,8) ,
9119	 => std_logic_vector(to_unsigned(88,8) ,
9120	 => std_logic_vector(to_unsigned(92,8) ,
9121	 => std_logic_vector(to_unsigned(91,8) ,
9122	 => std_logic_vector(to_unsigned(95,8) ,
9123	 => std_logic_vector(to_unsigned(88,8) ,
9124	 => std_logic_vector(to_unsigned(90,8) ,
9125	 => std_logic_vector(to_unsigned(92,8) ,
9126	 => std_logic_vector(to_unsigned(85,8) ,
9127	 => std_logic_vector(to_unsigned(85,8) ,
9128	 => std_logic_vector(to_unsigned(84,8) ,
9129	 => std_logic_vector(to_unsigned(84,8) ,
9130	 => std_logic_vector(to_unsigned(90,8) ,
9131	 => std_logic_vector(to_unsigned(90,8) ,
9132	 => std_logic_vector(to_unsigned(85,8) ,
9133	 => std_logic_vector(to_unsigned(85,8) ,
9134	 => std_logic_vector(to_unsigned(82,8) ,
9135	 => std_logic_vector(to_unsigned(63,8) ,
9136	 => std_logic_vector(to_unsigned(69,8) ,
9137	 => std_logic_vector(to_unsigned(70,8) ,
9138	 => std_logic_vector(to_unsigned(68,8) ,
9139	 => std_logic_vector(to_unsigned(68,8) ,
9140	 => std_logic_vector(to_unsigned(68,8) ,
9141	 => std_logic_vector(to_unsigned(78,8) ,
9142	 => std_logic_vector(to_unsigned(73,8) ,
9143	 => std_logic_vector(to_unsigned(69,8) ,
9144	 => std_logic_vector(to_unsigned(59,8) ,
9145	 => std_logic_vector(to_unsigned(62,8) ,
9146	 => std_logic_vector(to_unsigned(61,8) ,
9147	 => std_logic_vector(to_unsigned(60,8) ,
9148	 => std_logic_vector(to_unsigned(61,8) ,
9149	 => std_logic_vector(to_unsigned(63,8) ,
9150	 => std_logic_vector(to_unsigned(70,8) ,
9151	 => std_logic_vector(to_unsigned(71,8) ,
9152	 => std_logic_vector(to_unsigned(77,8) ,
9153	 => std_logic_vector(to_unsigned(81,8) ,
9154	 => std_logic_vector(to_unsigned(73,8) ,
9155	 => std_logic_vector(to_unsigned(74,8) ,
9156	 => std_logic_vector(to_unsigned(76,8) ,
9157	 => std_logic_vector(to_unsigned(73,8) ,
9158	 => std_logic_vector(to_unsigned(73,8) ,
9159	 => std_logic_vector(to_unsigned(61,8) ,
9160	 => std_logic_vector(to_unsigned(73,8) ,
9161	 => std_logic_vector(to_unsigned(72,8) ,
9162	 => std_logic_vector(to_unsigned(65,8) ,
9163	 => std_logic_vector(to_unsigned(84,8) ,
9164	 => std_logic_vector(to_unsigned(88,8) ,
9165	 => std_logic_vector(to_unsigned(91,8) ,
9166	 => std_logic_vector(to_unsigned(82,8) ,
9167	 => std_logic_vector(to_unsigned(73,8) ,
9168	 => std_logic_vector(to_unsigned(78,8) ,
9169	 => std_logic_vector(to_unsigned(76,8) ,
9170	 => std_logic_vector(to_unsigned(84,8) ,
9171	 => std_logic_vector(to_unsigned(88,8) ,
9172	 => std_logic_vector(to_unsigned(80,8) ,
9173	 => std_logic_vector(to_unsigned(77,8) ,
9174	 => std_logic_vector(to_unsigned(74,8) ,
9175	 => std_logic_vector(to_unsigned(78,8) ,
9176	 => std_logic_vector(to_unsigned(79,8) ,
9177	 => std_logic_vector(to_unsigned(78,8) ,
9178	 => std_logic_vector(to_unsigned(84,8) ,
9179	 => std_logic_vector(to_unsigned(70,8) ,
9180	 => std_logic_vector(to_unsigned(62,8) ,
9181	 => std_logic_vector(to_unsigned(82,8) ,
9182	 => std_logic_vector(to_unsigned(76,8) ,
9183	 => std_logic_vector(to_unsigned(64,8) ,
9184	 => std_logic_vector(to_unsigned(84,8) ,
9185	 => std_logic_vector(to_unsigned(79,8) ,
9186	 => std_logic_vector(to_unsigned(86,8) ,
9187	 => std_logic_vector(to_unsigned(81,8) ,
9188	 => std_logic_vector(to_unsigned(64,8) ,
9189	 => std_logic_vector(to_unsigned(66,8) ,
9190	 => std_logic_vector(to_unsigned(72,8) ,
9191	 => std_logic_vector(to_unsigned(67,8) ,
9192	 => std_logic_vector(to_unsigned(57,8) ,
9193	 => std_logic_vector(to_unsigned(65,8) ,
9194	 => std_logic_vector(to_unsigned(51,8) ,
9195	 => std_logic_vector(to_unsigned(56,8) ,
9196	 => std_logic_vector(to_unsigned(59,8) ,
9197	 => std_logic_vector(to_unsigned(59,8) ,
9198	 => std_logic_vector(to_unsigned(57,8) ,
9199	 => std_logic_vector(to_unsigned(55,8) ,
9200	 => std_logic_vector(to_unsigned(63,8) ,
9201	 => std_logic_vector(to_unsigned(47,8) ,
9202	 => std_logic_vector(to_unsigned(3,8) ,
9203	 => std_logic_vector(to_unsigned(0,8) ,
9204	 => std_logic_vector(to_unsigned(0,8) ,
9205	 => std_logic_vector(to_unsigned(28,8) ,
9206	 => std_logic_vector(to_unsigned(90,8) ,
9207	 => std_logic_vector(to_unsigned(81,8) ,
9208	 => std_logic_vector(to_unsigned(81,8) ,
9209	 => std_logic_vector(to_unsigned(81,8) ,
9210	 => std_logic_vector(to_unsigned(87,8) ,
9211	 => std_logic_vector(to_unsigned(92,8) ,
9212	 => std_logic_vector(to_unsigned(92,8) ,
9213	 => std_logic_vector(to_unsigned(90,8) ,
9214	 => std_logic_vector(to_unsigned(99,8) ,
9215	 => std_logic_vector(to_unsigned(92,8) ,
9216	 => std_logic_vector(to_unsigned(82,8) ,
9217	 => std_logic_vector(to_unsigned(87,8) ,
9218	 => std_logic_vector(to_unsigned(80,8) ,
9219	 => std_logic_vector(to_unsigned(82,8) ,
9220	 => std_logic_vector(to_unsigned(90,8) ,
9221	 => std_logic_vector(to_unsigned(90,8) ,
9222	 => std_logic_vector(to_unsigned(103,8) ,
9223	 => std_logic_vector(to_unsigned(103,8) ,
9224	 => std_logic_vector(to_unsigned(85,8) ,
9225	 => std_logic_vector(to_unsigned(85,8) ,
9226	 => std_logic_vector(to_unsigned(87,8) ,
9227	 => std_logic_vector(to_unsigned(88,8) ,
9228	 => std_logic_vector(to_unsigned(88,8) ,
9229	 => std_logic_vector(to_unsigned(85,8) ,
9230	 => std_logic_vector(to_unsigned(88,8) ,
9231	 => std_logic_vector(to_unsigned(90,8) ,
9232	 => std_logic_vector(to_unsigned(87,8) ,
9233	 => std_logic_vector(to_unsigned(92,8) ,
9234	 => std_logic_vector(to_unsigned(88,8) ,
9235	 => std_logic_vector(to_unsigned(88,8) ,
9236	 => std_logic_vector(to_unsigned(90,8) ,
9237	 => std_logic_vector(to_unsigned(88,8) ,
9238	 => std_logic_vector(to_unsigned(97,8) ,
9239	 => std_logic_vector(to_unsigned(96,8) ,
9240	 => std_logic_vector(to_unsigned(100,8) ,
9241	 => std_logic_vector(to_unsigned(103,8) ,
9242	 => std_logic_vector(to_unsigned(97,8) ,
9243	 => std_logic_vector(to_unsigned(97,8) ,
9244	 => std_logic_vector(to_unsigned(97,8) ,
9245	 => std_logic_vector(to_unsigned(105,8) ,
9246	 => std_logic_vector(to_unsigned(108,8) ,
9247	 => std_logic_vector(to_unsigned(108,8) ,
9248	 => std_logic_vector(to_unsigned(105,8) ,
9249	 => std_logic_vector(to_unsigned(105,8) ,
9250	 => std_logic_vector(to_unsigned(109,8) ,
9251	 => std_logic_vector(to_unsigned(103,8) ,
9252	 => std_logic_vector(to_unsigned(107,8) ,
9253	 => std_logic_vector(to_unsigned(111,8) ,
9254	 => std_logic_vector(to_unsigned(109,8) ,
9255	 => std_logic_vector(to_unsigned(108,8) ,
9256	 => std_logic_vector(to_unsigned(111,8) ,
9257	 => std_logic_vector(to_unsigned(112,8) ,
9258	 => std_logic_vector(to_unsigned(111,8) ,
9259	 => std_logic_vector(to_unsigned(116,8) ,
9260	 => std_logic_vector(to_unsigned(122,8) ,
9261	 => std_logic_vector(to_unsigned(127,8) ,
9262	 => std_logic_vector(to_unsigned(131,8) ,
9263	 => std_logic_vector(to_unsigned(134,8) ,
9264	 => std_logic_vector(to_unsigned(133,8) ,
9265	 => std_logic_vector(to_unsigned(136,8) ,
9266	 => std_logic_vector(to_unsigned(142,8) ,
9267	 => std_logic_vector(to_unsigned(142,8) ,
9268	 => std_logic_vector(to_unsigned(142,8) ,
9269	 => std_logic_vector(to_unsigned(144,8) ,
9270	 => std_logic_vector(to_unsigned(147,8) ,
9271	 => std_logic_vector(to_unsigned(151,8) ,
9272	 => std_logic_vector(to_unsigned(151,8) ,
9273	 => std_logic_vector(to_unsigned(147,8) ,
9274	 => std_logic_vector(to_unsigned(149,8) ,
9275	 => std_logic_vector(to_unsigned(151,8) ,
9276	 => std_logic_vector(to_unsigned(146,8) ,
9277	 => std_logic_vector(to_unsigned(138,8) ,
9278	 => std_logic_vector(to_unsigned(141,8) ,
9279	 => std_logic_vector(to_unsigned(146,8) ,
9280	 => std_logic_vector(to_unsigned(146,8) ,
9281	 => std_logic_vector(to_unsigned(87,8) ,
9282	 => std_logic_vector(to_unsigned(87,8) ,
9283	 => std_logic_vector(to_unsigned(81,8) ,
9284	 => std_logic_vector(to_unsigned(71,8) ,
9285	 => std_logic_vector(to_unsigned(77,8) ,
9286	 => std_logic_vector(to_unsigned(81,8) ,
9287	 => std_logic_vector(to_unsigned(84,8) ,
9288	 => std_logic_vector(to_unsigned(82,8) ,
9289	 => std_logic_vector(to_unsigned(80,8) ,
9290	 => std_logic_vector(to_unsigned(82,8) ,
9291	 => std_logic_vector(to_unsigned(86,8) ,
9292	 => std_logic_vector(to_unsigned(85,8) ,
9293	 => std_logic_vector(to_unsigned(84,8) ,
9294	 => std_logic_vector(to_unsigned(87,8) ,
9295	 => std_logic_vector(to_unsigned(88,8) ,
9296	 => std_logic_vector(to_unsigned(87,8) ,
9297	 => std_logic_vector(to_unsigned(87,8) ,
9298	 => std_logic_vector(to_unsigned(82,8) ,
9299	 => std_logic_vector(to_unsigned(79,8) ,
9300	 => std_logic_vector(to_unsigned(90,8) ,
9301	 => std_logic_vector(to_unsigned(93,8) ,
9302	 => std_logic_vector(to_unsigned(84,8) ,
9303	 => std_logic_vector(to_unsigned(82,8) ,
9304	 => std_logic_vector(to_unsigned(81,8) ,
9305	 => std_logic_vector(to_unsigned(85,8) ,
9306	 => std_logic_vector(to_unsigned(91,8) ,
9307	 => std_logic_vector(to_unsigned(85,8) ,
9308	 => std_logic_vector(to_unsigned(80,8) ,
9309	 => std_logic_vector(to_unsigned(85,8) ,
9310	 => std_logic_vector(to_unsigned(84,8) ,
9311	 => std_logic_vector(to_unsigned(90,8) ,
9312	 => std_logic_vector(to_unsigned(86,8) ,
9313	 => std_logic_vector(to_unsigned(84,8) ,
9314	 => std_logic_vector(to_unsigned(88,8) ,
9315	 => std_logic_vector(to_unsigned(90,8) ,
9316	 => std_logic_vector(to_unsigned(86,8) ,
9317	 => std_logic_vector(to_unsigned(87,8) ,
9318	 => std_logic_vector(to_unsigned(88,8) ,
9319	 => std_logic_vector(to_unsigned(87,8) ,
9320	 => std_logic_vector(to_unsigned(86,8) ,
9321	 => std_logic_vector(to_unsigned(85,8) ,
9322	 => std_logic_vector(to_unsigned(90,8) ,
9323	 => std_logic_vector(to_unsigned(97,8) ,
9324	 => std_logic_vector(to_unsigned(93,8) ,
9325	 => std_logic_vector(to_unsigned(95,8) ,
9326	 => std_logic_vector(to_unsigned(99,8) ,
9327	 => std_logic_vector(to_unsigned(100,8) ,
9328	 => std_logic_vector(to_unsigned(100,8) ,
9329	 => std_logic_vector(to_unsigned(101,8) ,
9330	 => std_logic_vector(to_unsigned(100,8) ,
9331	 => std_logic_vector(to_unsigned(100,8) ,
9332	 => std_logic_vector(to_unsigned(105,8) ,
9333	 => std_logic_vector(to_unsigned(104,8) ,
9334	 => std_logic_vector(to_unsigned(101,8) ,
9335	 => std_logic_vector(to_unsigned(101,8) ,
9336	 => std_logic_vector(to_unsigned(99,8) ,
9337	 => std_logic_vector(to_unsigned(107,8) ,
9338	 => std_logic_vector(to_unsigned(115,8) ,
9339	 => std_logic_vector(to_unsigned(116,8) ,
9340	 => std_logic_vector(to_unsigned(119,8) ,
9341	 => std_logic_vector(to_unsigned(127,8) ,
9342	 => std_logic_vector(to_unsigned(124,8) ,
9343	 => std_logic_vector(to_unsigned(130,8) ,
9344	 => std_logic_vector(to_unsigned(134,8) ,
9345	 => std_logic_vector(to_unsigned(128,8) ,
9346	 => std_logic_vector(to_unsigned(127,8) ,
9347	 => std_logic_vector(to_unsigned(131,8) ,
9348	 => std_logic_vector(to_unsigned(130,8) ,
9349	 => std_logic_vector(to_unsigned(136,8) ,
9350	 => std_logic_vector(to_unsigned(133,8) ,
9351	 => std_logic_vector(to_unsigned(130,8) ,
9352	 => std_logic_vector(to_unsigned(131,8) ,
9353	 => std_logic_vector(to_unsigned(127,8) ,
9354	 => std_logic_vector(to_unsigned(133,8) ,
9355	 => std_logic_vector(to_unsigned(134,8) ,
9356	 => std_logic_vector(to_unsigned(121,8) ,
9357	 => std_logic_vector(to_unsigned(128,8) ,
9358	 => std_logic_vector(to_unsigned(134,8) ,
9359	 => std_logic_vector(to_unsigned(131,8) ,
9360	 => std_logic_vector(to_unsigned(128,8) ,
9361	 => std_logic_vector(to_unsigned(128,8) ,
9362	 => std_logic_vector(to_unsigned(130,8) ,
9363	 => std_logic_vector(to_unsigned(127,8) ,
9364	 => std_logic_vector(to_unsigned(128,8) ,
9365	 => std_logic_vector(to_unsigned(131,8) ,
9366	 => std_logic_vector(to_unsigned(125,8) ,
9367	 => std_logic_vector(to_unsigned(119,8) ,
9368	 => std_logic_vector(to_unsigned(118,8) ,
9369	 => std_logic_vector(to_unsigned(121,8) ,
9370	 => std_logic_vector(to_unsigned(128,8) ,
9371	 => std_logic_vector(to_unsigned(125,8) ,
9372	 => std_logic_vector(to_unsigned(119,8) ,
9373	 => std_logic_vector(to_unsigned(121,8) ,
9374	 => std_logic_vector(to_unsigned(125,8) ,
9375	 => std_logic_vector(to_unsigned(122,8) ,
9376	 => std_logic_vector(to_unsigned(121,8) ,
9377	 => std_logic_vector(to_unsigned(109,8) ,
9378	 => std_logic_vector(to_unsigned(103,8) ,
9379	 => std_logic_vector(to_unsigned(105,8) ,
9380	 => std_logic_vector(to_unsigned(105,8) ,
9381	 => std_logic_vector(to_unsigned(105,8) ,
9382	 => std_logic_vector(to_unsigned(105,8) ,
9383	 => std_logic_vector(to_unsigned(99,8) ,
9384	 => std_logic_vector(to_unsigned(97,8) ,
9385	 => std_logic_vector(to_unsigned(103,8) ,
9386	 => std_logic_vector(to_unsigned(100,8) ,
9387	 => std_logic_vector(to_unsigned(101,8) ,
9388	 => std_logic_vector(to_unsigned(99,8) ,
9389	 => std_logic_vector(to_unsigned(97,8) ,
9390	 => std_logic_vector(to_unsigned(97,8) ,
9391	 => std_logic_vector(to_unsigned(82,8) ,
9392	 => std_logic_vector(to_unsigned(85,8) ,
9393	 => std_logic_vector(to_unsigned(90,8) ,
9394	 => std_logic_vector(to_unsigned(92,8) ,
9395	 => std_logic_vector(to_unsigned(97,8) ,
9396	 => std_logic_vector(to_unsigned(103,8) ,
9397	 => std_logic_vector(to_unsigned(97,8) ,
9398	 => std_logic_vector(to_unsigned(104,8) ,
9399	 => std_logic_vector(to_unsigned(107,8) ,
9400	 => std_logic_vector(to_unsigned(97,8) ,
9401	 => std_logic_vector(to_unsigned(92,8) ,
9402	 => std_logic_vector(to_unsigned(88,8) ,
9403	 => std_logic_vector(to_unsigned(87,8) ,
9404	 => std_logic_vector(to_unsigned(93,8) ,
9405	 => std_logic_vector(to_unsigned(99,8) ,
9406	 => std_logic_vector(to_unsigned(99,8) ,
9407	 => std_logic_vector(to_unsigned(97,8) ,
9408	 => std_logic_vector(to_unsigned(101,8) ,
9409	 => std_logic_vector(to_unsigned(105,8) ,
9410	 => std_logic_vector(to_unsigned(111,8) ,
9411	 => std_logic_vector(to_unsigned(115,8) ,
9412	 => std_logic_vector(to_unsigned(121,8) ,
9413	 => std_logic_vector(to_unsigned(119,8) ,
9414	 => std_logic_vector(to_unsigned(109,8) ,
9415	 => std_logic_vector(to_unsigned(101,8) ,
9416	 => std_logic_vector(to_unsigned(105,8) ,
9417	 => std_logic_vector(to_unsigned(111,8) ,
9418	 => std_logic_vector(to_unsigned(101,8) ,
9419	 => std_logic_vector(to_unsigned(104,8) ,
9420	 => std_logic_vector(to_unsigned(105,8) ,
9421	 => std_logic_vector(to_unsigned(108,8) ,
9422	 => std_logic_vector(to_unsigned(114,8) ,
9423	 => std_logic_vector(to_unsigned(114,8) ,
9424	 => std_logic_vector(to_unsigned(108,8) ,
9425	 => std_logic_vector(to_unsigned(103,8) ,
9426	 => std_logic_vector(to_unsigned(104,8) ,
9427	 => std_logic_vector(to_unsigned(97,8) ,
9428	 => std_logic_vector(to_unsigned(84,8) ,
9429	 => std_logic_vector(to_unsigned(87,8) ,
9430	 => std_logic_vector(to_unsigned(92,8) ,
9431	 => std_logic_vector(to_unsigned(84,8) ,
9432	 => std_logic_vector(to_unsigned(88,8) ,
9433	 => std_logic_vector(to_unsigned(95,8) ,
9434	 => std_logic_vector(to_unsigned(92,8) ,
9435	 => std_logic_vector(to_unsigned(99,8) ,
9436	 => std_logic_vector(to_unsigned(95,8) ,
9437	 => std_logic_vector(to_unsigned(91,8) ,
9438	 => std_logic_vector(to_unsigned(93,8) ,
9439	 => std_logic_vector(to_unsigned(90,8) ,
9440	 => std_logic_vector(to_unsigned(80,8) ,
9441	 => std_logic_vector(to_unsigned(79,8) ,
9442	 => std_logic_vector(to_unsigned(80,8) ,
9443	 => std_logic_vector(to_unsigned(90,8) ,
9444	 => std_logic_vector(to_unsigned(100,8) ,
9445	 => std_logic_vector(to_unsigned(93,8) ,
9446	 => std_logic_vector(to_unsigned(90,8) ,
9447	 => std_logic_vector(to_unsigned(88,8) ,
9448	 => std_logic_vector(to_unsigned(79,8) ,
9449	 => std_logic_vector(to_unsigned(82,8) ,
9450	 => std_logic_vector(to_unsigned(96,8) ,
9451	 => std_logic_vector(to_unsigned(99,8) ,
9452	 => std_logic_vector(to_unsigned(91,8) ,
9453	 => std_logic_vector(to_unsigned(80,8) ,
9454	 => std_logic_vector(to_unsigned(74,8) ,
9455	 => std_logic_vector(to_unsigned(68,8) ,
9456	 => std_logic_vector(to_unsigned(74,8) ,
9457	 => std_logic_vector(to_unsigned(76,8) ,
9458	 => std_logic_vector(to_unsigned(65,8) ,
9459	 => std_logic_vector(to_unsigned(73,8) ,
9460	 => std_logic_vector(to_unsigned(78,8) ,
9461	 => std_logic_vector(to_unsigned(65,8) ,
9462	 => std_logic_vector(to_unsigned(65,8) ,
9463	 => std_logic_vector(to_unsigned(73,8) ,
9464	 => std_logic_vector(to_unsigned(72,8) ,
9465	 => std_logic_vector(to_unsigned(73,8) ,
9466	 => std_logic_vector(to_unsigned(70,8) ,
9467	 => std_logic_vector(to_unsigned(67,8) ,
9468	 => std_logic_vector(to_unsigned(74,8) ,
9469	 => std_logic_vector(to_unsigned(73,8) ,
9470	 => std_logic_vector(to_unsigned(81,8) ,
9471	 => std_logic_vector(to_unsigned(101,8) ,
9472	 => std_logic_vector(to_unsigned(84,8) ,
9473	 => std_logic_vector(to_unsigned(73,8) ,
9474	 => std_logic_vector(to_unsigned(80,8) ,
9475	 => std_logic_vector(to_unsigned(68,8) ,
9476	 => std_logic_vector(to_unsigned(61,8) ,
9477	 => std_logic_vector(to_unsigned(68,8) ,
9478	 => std_logic_vector(to_unsigned(78,8) ,
9479	 => std_logic_vector(to_unsigned(62,8) ,
9480	 => std_logic_vector(to_unsigned(76,8) ,
9481	 => std_logic_vector(to_unsigned(79,8) ,
9482	 => std_logic_vector(to_unsigned(72,8) ,
9483	 => std_logic_vector(to_unsigned(74,8) ,
9484	 => std_logic_vector(to_unsigned(76,8) ,
9485	 => std_logic_vector(to_unsigned(90,8) ,
9486	 => std_logic_vector(to_unsigned(87,8) ,
9487	 => std_logic_vector(to_unsigned(73,8) ,
9488	 => std_logic_vector(to_unsigned(77,8) ,
9489	 => std_logic_vector(to_unsigned(76,8) ,
9490	 => std_logic_vector(to_unsigned(81,8) ,
9491	 => std_logic_vector(to_unsigned(80,8) ,
9492	 => std_logic_vector(to_unsigned(76,8) ,
9493	 => std_logic_vector(to_unsigned(77,8) ,
9494	 => std_logic_vector(to_unsigned(72,8) ,
9495	 => std_logic_vector(to_unsigned(71,8) ,
9496	 => std_logic_vector(to_unsigned(70,8) ,
9497	 => std_logic_vector(to_unsigned(70,8) ,
9498	 => std_logic_vector(to_unsigned(77,8) ,
9499	 => std_logic_vector(to_unsigned(68,8) ,
9500	 => std_logic_vector(to_unsigned(57,8) ,
9501	 => std_logic_vector(to_unsigned(64,8) ,
9502	 => std_logic_vector(to_unsigned(77,8) ,
9503	 => std_logic_vector(to_unsigned(76,8) ,
9504	 => std_logic_vector(to_unsigned(79,8) ,
9505	 => std_logic_vector(to_unsigned(76,8) ,
9506	 => std_logic_vector(to_unsigned(85,8) ,
9507	 => std_logic_vector(to_unsigned(79,8) ,
9508	 => std_logic_vector(to_unsigned(69,8) ,
9509	 => std_logic_vector(to_unsigned(78,8) ,
9510	 => std_logic_vector(to_unsigned(71,8) ,
9511	 => std_logic_vector(to_unsigned(60,8) ,
9512	 => std_logic_vector(to_unsigned(65,8) ,
9513	 => std_logic_vector(to_unsigned(77,8) ,
9514	 => std_logic_vector(to_unsigned(69,8) ,
9515	 => std_logic_vector(to_unsigned(73,8) ,
9516	 => std_logic_vector(to_unsigned(56,8) ,
9517	 => std_logic_vector(to_unsigned(49,8) ,
9518	 => std_logic_vector(to_unsigned(53,8) ,
9519	 => std_logic_vector(to_unsigned(55,8) ,
9520	 => std_logic_vector(to_unsigned(68,8) ,
9521	 => std_logic_vector(to_unsigned(58,8) ,
9522	 => std_logic_vector(to_unsigned(5,8) ,
9523	 => std_logic_vector(to_unsigned(0,8) ,
9524	 => std_logic_vector(to_unsigned(0,8) ,
9525	 => std_logic_vector(to_unsigned(18,8) ,
9526	 => std_logic_vector(to_unsigned(85,8) ,
9527	 => std_logic_vector(to_unsigned(81,8) ,
9528	 => std_logic_vector(to_unsigned(90,8) ,
9529	 => std_logic_vector(to_unsigned(93,8) ,
9530	 => std_logic_vector(to_unsigned(96,8) ,
9531	 => std_logic_vector(to_unsigned(108,8) ,
9532	 => std_logic_vector(to_unsigned(99,8) ,
9533	 => std_logic_vector(to_unsigned(78,8) ,
9534	 => std_logic_vector(to_unsigned(93,8) ,
9535	 => std_logic_vector(to_unsigned(92,8) ,
9536	 => std_logic_vector(to_unsigned(78,8) ,
9537	 => std_logic_vector(to_unsigned(77,8) ,
9538	 => std_logic_vector(to_unsigned(79,8) ,
9539	 => std_logic_vector(to_unsigned(86,8) ,
9540	 => std_logic_vector(to_unsigned(87,8) ,
9541	 => std_logic_vector(to_unsigned(97,8) ,
9542	 => std_logic_vector(to_unsigned(112,8) ,
9543	 => std_logic_vector(to_unsigned(101,8) ,
9544	 => std_logic_vector(to_unsigned(84,8) ,
9545	 => std_logic_vector(to_unsigned(88,8) ,
9546	 => std_logic_vector(to_unsigned(88,8) ,
9547	 => std_logic_vector(to_unsigned(90,8) ,
9548	 => std_logic_vector(to_unsigned(93,8) ,
9549	 => std_logic_vector(to_unsigned(87,8) ,
9550	 => std_logic_vector(to_unsigned(86,8) ,
9551	 => std_logic_vector(to_unsigned(90,8) ,
9552	 => std_logic_vector(to_unsigned(91,8) ,
9553	 => std_logic_vector(to_unsigned(92,8) ,
9554	 => std_logic_vector(to_unsigned(87,8) ,
9555	 => std_logic_vector(to_unsigned(88,8) ,
9556	 => std_logic_vector(to_unsigned(91,8) ,
9557	 => std_logic_vector(to_unsigned(88,8) ,
9558	 => std_logic_vector(to_unsigned(91,8) ,
9559	 => std_logic_vector(to_unsigned(90,8) ,
9560	 => std_logic_vector(to_unsigned(91,8) ,
9561	 => std_logic_vector(to_unsigned(91,8) ,
9562	 => std_logic_vector(to_unsigned(87,8) ,
9563	 => std_logic_vector(to_unsigned(90,8) ,
9564	 => std_logic_vector(to_unsigned(91,8) ,
9565	 => std_logic_vector(to_unsigned(95,8) ,
9566	 => std_logic_vector(to_unsigned(99,8) ,
9567	 => std_logic_vector(to_unsigned(99,8) ,
9568	 => std_logic_vector(to_unsigned(97,8) ,
9569	 => std_logic_vector(to_unsigned(95,8) ,
9570	 => std_logic_vector(to_unsigned(93,8) ,
9571	 => std_logic_vector(to_unsigned(99,8) ,
9572	 => std_logic_vector(to_unsigned(97,8) ,
9573	 => std_logic_vector(to_unsigned(100,8) ,
9574	 => std_logic_vector(to_unsigned(108,8) ,
9575	 => std_logic_vector(to_unsigned(112,8) ,
9576	 => std_logic_vector(to_unsigned(104,8) ,
9577	 => std_logic_vector(to_unsigned(107,8) ,
9578	 => std_logic_vector(to_unsigned(111,8) ,
9579	 => std_logic_vector(to_unsigned(111,8) ,
9580	 => std_logic_vector(to_unsigned(115,8) ,
9581	 => std_logic_vector(to_unsigned(122,8) ,
9582	 => std_logic_vector(to_unsigned(127,8) ,
9583	 => std_logic_vector(to_unsigned(125,8) ,
9584	 => std_logic_vector(to_unsigned(128,8) ,
9585	 => std_logic_vector(to_unsigned(130,8) ,
9586	 => std_logic_vector(to_unsigned(134,8) ,
9587	 => std_logic_vector(to_unsigned(142,8) ,
9588	 => std_logic_vector(to_unsigned(142,8) ,
9589	 => std_logic_vector(to_unsigned(146,8) ,
9590	 => std_logic_vector(to_unsigned(151,8) ,
9591	 => std_logic_vector(to_unsigned(154,8) ,
9592	 => std_logic_vector(to_unsigned(151,8) ,
9593	 => std_logic_vector(to_unsigned(151,8) ,
9594	 => std_logic_vector(to_unsigned(154,8) ,
9595	 => std_logic_vector(to_unsigned(151,8) ,
9596	 => std_logic_vector(to_unsigned(149,8) ,
9597	 => std_logic_vector(to_unsigned(146,8) ,
9598	 => std_logic_vector(to_unsigned(147,8) ,
9599	 => std_logic_vector(to_unsigned(149,8) ,
9600	 => std_logic_vector(to_unsigned(149,8) ,
9601	 => std_logic_vector(to_unsigned(105,8) ,
9602	 => std_logic_vector(to_unsigned(108,8) ,
9603	 => std_logic_vector(to_unsigned(99,8) ,
9604	 => std_logic_vector(to_unsigned(88,8) ,
9605	 => std_logic_vector(to_unsigned(93,8) ,
9606	 => std_logic_vector(to_unsigned(92,8) ,
9607	 => std_logic_vector(to_unsigned(82,8) ,
9608	 => std_logic_vector(to_unsigned(86,8) ,
9609	 => std_logic_vector(to_unsigned(91,8) ,
9610	 => std_logic_vector(to_unsigned(88,8) ,
9611	 => std_logic_vector(to_unsigned(87,8) ,
9612	 => std_logic_vector(to_unsigned(86,8) ,
9613	 => std_logic_vector(to_unsigned(85,8) ,
9614	 => std_logic_vector(to_unsigned(90,8) ,
9615	 => std_logic_vector(to_unsigned(90,8) ,
9616	 => std_logic_vector(to_unsigned(85,8) ,
9617	 => std_logic_vector(to_unsigned(86,8) ,
9618	 => std_logic_vector(to_unsigned(86,8) ,
9619	 => std_logic_vector(to_unsigned(81,8) ,
9620	 => std_logic_vector(to_unsigned(90,8) ,
9621	 => std_logic_vector(to_unsigned(95,8) ,
9622	 => std_logic_vector(to_unsigned(88,8) ,
9623	 => std_logic_vector(to_unsigned(91,8) ,
9624	 => std_logic_vector(to_unsigned(87,8) ,
9625	 => std_logic_vector(to_unsigned(97,8) ,
9626	 => std_logic_vector(to_unsigned(100,8) ,
9627	 => std_logic_vector(to_unsigned(97,8) ,
9628	 => std_logic_vector(to_unsigned(101,8) ,
9629	 => std_logic_vector(to_unsigned(93,8) ,
9630	 => std_logic_vector(to_unsigned(96,8) ,
9631	 => std_logic_vector(to_unsigned(103,8) ,
9632	 => std_logic_vector(to_unsigned(88,8) ,
9633	 => std_logic_vector(to_unsigned(88,8) ,
9634	 => std_logic_vector(to_unsigned(93,8) ,
9635	 => std_logic_vector(to_unsigned(92,8) ,
9636	 => std_logic_vector(to_unsigned(88,8) ,
9637	 => std_logic_vector(to_unsigned(87,8) ,
9638	 => std_logic_vector(to_unsigned(91,8) ,
9639	 => std_logic_vector(to_unsigned(90,8) ,
9640	 => std_logic_vector(to_unsigned(90,8) ,
9641	 => std_logic_vector(to_unsigned(93,8) ,
9642	 => std_logic_vector(to_unsigned(105,8) ,
9643	 => std_logic_vector(to_unsigned(105,8) ,
9644	 => std_logic_vector(to_unsigned(100,8) ,
9645	 => std_logic_vector(to_unsigned(108,8) ,
9646	 => std_logic_vector(to_unsigned(108,8) ,
9647	 => std_logic_vector(to_unsigned(103,8) ,
9648	 => std_logic_vector(to_unsigned(107,8) ,
9649	 => std_logic_vector(to_unsigned(118,8) ,
9650	 => std_logic_vector(to_unsigned(118,8) ,
9651	 => std_logic_vector(to_unsigned(115,8) ,
9652	 => std_logic_vector(to_unsigned(118,8) ,
9653	 => std_logic_vector(to_unsigned(121,8) ,
9654	 => std_logic_vector(to_unsigned(118,8) ,
9655	 => std_logic_vector(to_unsigned(114,8) ,
9656	 => std_logic_vector(to_unsigned(112,8) ,
9657	 => std_logic_vector(to_unsigned(118,8) ,
9658	 => std_logic_vector(to_unsigned(127,8) ,
9659	 => std_logic_vector(to_unsigned(130,8) ,
9660	 => std_logic_vector(to_unsigned(133,8) ,
9661	 => std_logic_vector(to_unsigned(136,8) ,
9662	 => std_logic_vector(to_unsigned(133,8) ,
9663	 => std_logic_vector(to_unsigned(141,8) ,
9664	 => std_logic_vector(to_unsigned(141,8) ,
9665	 => std_logic_vector(to_unsigned(134,8) ,
9666	 => std_logic_vector(to_unsigned(133,8) ,
9667	 => std_logic_vector(to_unsigned(142,8) ,
9668	 => std_logic_vector(to_unsigned(136,8) ,
9669	 => std_logic_vector(to_unsigned(133,8) ,
9670	 => std_logic_vector(to_unsigned(136,8) ,
9671	 => std_logic_vector(to_unsigned(142,8) ,
9672	 => std_logic_vector(to_unsigned(142,8) ,
9673	 => std_logic_vector(to_unsigned(138,8) ,
9674	 => std_logic_vector(to_unsigned(141,8) ,
9675	 => std_logic_vector(to_unsigned(139,8) ,
9676	 => std_logic_vector(to_unsigned(134,8) ,
9677	 => std_logic_vector(to_unsigned(138,8) ,
9678	 => std_logic_vector(to_unsigned(141,8) ,
9679	 => std_logic_vector(to_unsigned(136,8) ,
9680	 => std_logic_vector(to_unsigned(134,8) ,
9681	 => std_logic_vector(to_unsigned(134,8) ,
9682	 => std_logic_vector(to_unsigned(133,8) ,
9683	 => std_logic_vector(to_unsigned(127,8) ,
9684	 => std_logic_vector(to_unsigned(127,8) ,
9685	 => std_logic_vector(to_unsigned(134,8) ,
9686	 => std_logic_vector(to_unsigned(133,8) ,
9687	 => std_logic_vector(to_unsigned(130,8) ,
9688	 => std_logic_vector(to_unsigned(128,8) ,
9689	 => std_logic_vector(to_unsigned(127,8) ,
9690	 => std_logic_vector(to_unsigned(128,8) ,
9691	 => std_logic_vector(to_unsigned(131,8) ,
9692	 => std_logic_vector(to_unsigned(136,8) ,
9693	 => std_logic_vector(to_unsigned(130,8) ,
9694	 => std_logic_vector(to_unsigned(130,8) ,
9695	 => std_logic_vector(to_unsigned(127,8) ,
9696	 => std_logic_vector(to_unsigned(128,8) ,
9697	 => std_logic_vector(to_unsigned(122,8) ,
9698	 => std_logic_vector(to_unsigned(115,8) ,
9699	 => std_logic_vector(to_unsigned(115,8) ,
9700	 => std_logic_vector(to_unsigned(108,8) ,
9701	 => std_logic_vector(to_unsigned(107,8) ,
9702	 => std_logic_vector(to_unsigned(105,8) ,
9703	 => std_logic_vector(to_unsigned(99,8) ,
9704	 => std_logic_vector(to_unsigned(103,8) ,
9705	 => std_logic_vector(to_unsigned(101,8) ,
9706	 => std_logic_vector(to_unsigned(90,8) ,
9707	 => std_logic_vector(to_unsigned(92,8) ,
9708	 => std_logic_vector(to_unsigned(86,8) ,
9709	 => std_logic_vector(to_unsigned(81,8) ,
9710	 => std_logic_vector(to_unsigned(87,8) ,
9711	 => std_logic_vector(to_unsigned(73,8) ,
9712	 => std_logic_vector(to_unsigned(68,8) ,
9713	 => std_logic_vector(to_unsigned(74,8) ,
9714	 => std_logic_vector(to_unsigned(78,8) ,
9715	 => std_logic_vector(to_unsigned(79,8) ,
9716	 => std_logic_vector(to_unsigned(78,8) ,
9717	 => std_logic_vector(to_unsigned(77,8) ,
9718	 => std_logic_vector(to_unsigned(87,8) ,
9719	 => std_logic_vector(to_unsigned(95,8) ,
9720	 => std_logic_vector(to_unsigned(90,8) ,
9721	 => std_logic_vector(to_unsigned(90,8) ,
9722	 => std_logic_vector(to_unsigned(96,8) ,
9723	 => std_logic_vector(to_unsigned(92,8) ,
9724	 => std_logic_vector(to_unsigned(93,8) ,
9725	 => std_logic_vector(to_unsigned(108,8) ,
9726	 => std_logic_vector(to_unsigned(108,8) ,
9727	 => std_logic_vector(to_unsigned(93,8) ,
9728	 => std_logic_vector(to_unsigned(101,8) ,
9729	 => std_logic_vector(to_unsigned(105,8) ,
9730	 => std_logic_vector(to_unsigned(104,8) ,
9731	 => std_logic_vector(to_unsigned(108,8) ,
9732	 => std_logic_vector(to_unsigned(105,8) ,
9733	 => std_logic_vector(to_unsigned(107,8) ,
9734	 => std_logic_vector(to_unsigned(104,8) ,
9735	 => std_logic_vector(to_unsigned(100,8) ,
9736	 => std_logic_vector(to_unsigned(104,8) ,
9737	 => std_logic_vector(to_unsigned(107,8) ,
9738	 => std_logic_vector(to_unsigned(96,8) ,
9739	 => std_logic_vector(to_unsigned(92,8) ,
9740	 => std_logic_vector(to_unsigned(97,8) ,
9741	 => std_logic_vector(to_unsigned(108,8) ,
9742	 => std_logic_vector(to_unsigned(101,8) ,
9743	 => std_logic_vector(to_unsigned(96,8) ,
9744	 => std_logic_vector(to_unsigned(108,8) ,
9745	 => std_logic_vector(to_unsigned(111,8) ,
9746	 => std_logic_vector(to_unsigned(114,8) ,
9747	 => std_logic_vector(to_unsigned(116,8) ,
9748	 => std_logic_vector(to_unsigned(101,8) ,
9749	 => std_logic_vector(to_unsigned(92,8) ,
9750	 => std_logic_vector(to_unsigned(85,8) ,
9751	 => std_logic_vector(to_unsigned(77,8) ,
9752	 => std_logic_vector(to_unsigned(81,8) ,
9753	 => std_logic_vector(to_unsigned(92,8) ,
9754	 => std_logic_vector(to_unsigned(96,8) ,
9755	 => std_logic_vector(to_unsigned(103,8) ,
9756	 => std_logic_vector(to_unsigned(104,8) ,
9757	 => std_logic_vector(to_unsigned(95,8) ,
9758	 => std_logic_vector(to_unsigned(88,8) ,
9759	 => std_logic_vector(to_unsigned(86,8) ,
9760	 => std_logic_vector(to_unsigned(92,8) ,
9761	 => std_logic_vector(to_unsigned(82,8) ,
9762	 => std_logic_vector(to_unsigned(70,8) ,
9763	 => std_logic_vector(to_unsigned(84,8) ,
9764	 => std_logic_vector(to_unsigned(103,8) ,
9765	 => std_logic_vector(to_unsigned(96,8) ,
9766	 => std_logic_vector(to_unsigned(85,8) ,
9767	 => std_logic_vector(to_unsigned(80,8) ,
9768	 => std_logic_vector(to_unsigned(80,8) ,
9769	 => std_logic_vector(to_unsigned(82,8) ,
9770	 => std_logic_vector(to_unsigned(85,8) ,
9771	 => std_logic_vector(to_unsigned(92,8) ,
9772	 => std_logic_vector(to_unsigned(92,8) ,
9773	 => std_logic_vector(to_unsigned(77,8) ,
9774	 => std_logic_vector(to_unsigned(68,8) ,
9775	 => std_logic_vector(to_unsigned(76,8) ,
9776	 => std_logic_vector(to_unsigned(78,8) ,
9777	 => std_logic_vector(to_unsigned(82,8) ,
9778	 => std_logic_vector(to_unsigned(84,8) ,
9779	 => std_logic_vector(to_unsigned(85,8) ,
9780	 => std_logic_vector(to_unsigned(91,8) ,
9781	 => std_logic_vector(to_unsigned(79,8) ,
9782	 => std_logic_vector(to_unsigned(77,8) ,
9783	 => std_logic_vector(to_unsigned(81,8) ,
9784	 => std_logic_vector(to_unsigned(79,8) ,
9785	 => std_logic_vector(to_unsigned(79,8) ,
9786	 => std_logic_vector(to_unsigned(86,8) ,
9787	 => std_logic_vector(to_unsigned(87,8) ,
9788	 => std_logic_vector(to_unsigned(91,8) ,
9789	 => std_logic_vector(to_unsigned(92,8) ,
9790	 => std_logic_vector(to_unsigned(101,8) ,
9791	 => std_logic_vector(to_unsigned(100,8) ,
9792	 => std_logic_vector(to_unsigned(72,8) ,
9793	 => std_logic_vector(to_unsigned(76,8) ,
9794	 => std_logic_vector(to_unsigned(85,8) ,
9795	 => std_logic_vector(to_unsigned(76,8) ,
9796	 => std_logic_vector(to_unsigned(73,8) ,
9797	 => std_logic_vector(to_unsigned(81,8) ,
9798	 => std_logic_vector(to_unsigned(87,8) ,
9799	 => std_logic_vector(to_unsigned(74,8) ,
9800	 => std_logic_vector(to_unsigned(77,8) ,
9801	 => std_logic_vector(to_unsigned(87,8) ,
9802	 => std_logic_vector(to_unsigned(81,8) ,
9803	 => std_logic_vector(to_unsigned(80,8) ,
9804	 => std_logic_vector(to_unsigned(72,8) ,
9805	 => std_logic_vector(to_unsigned(77,8) ,
9806	 => std_logic_vector(to_unsigned(82,8) ,
9807	 => std_logic_vector(to_unsigned(79,8) ,
9808	 => std_logic_vector(to_unsigned(78,8) ,
9809	 => std_logic_vector(to_unsigned(86,8) ,
9810	 => std_logic_vector(to_unsigned(86,8) ,
9811	 => std_logic_vector(to_unsigned(78,8) ,
9812	 => std_logic_vector(to_unsigned(70,8) ,
9813	 => std_logic_vector(to_unsigned(71,8) ,
9814	 => std_logic_vector(to_unsigned(66,8) ,
9815	 => std_logic_vector(to_unsigned(61,8) ,
9816	 => std_logic_vector(to_unsigned(62,8) ,
9817	 => std_logic_vector(to_unsigned(66,8) ,
9818	 => std_logic_vector(to_unsigned(70,8) ,
9819	 => std_logic_vector(to_unsigned(73,8) ,
9820	 => std_logic_vector(to_unsigned(65,8) ,
9821	 => std_logic_vector(to_unsigned(64,8) ,
9822	 => std_logic_vector(to_unsigned(86,8) ,
9823	 => std_logic_vector(to_unsigned(100,8) ,
9824	 => std_logic_vector(to_unsigned(86,8) ,
9825	 => std_logic_vector(to_unsigned(64,8) ,
9826	 => std_logic_vector(to_unsigned(79,8) ,
9827	 => std_logic_vector(to_unsigned(76,8) ,
9828	 => std_logic_vector(to_unsigned(74,8) ,
9829	 => std_logic_vector(to_unsigned(78,8) ,
9830	 => std_logic_vector(to_unsigned(79,8) ,
9831	 => std_logic_vector(to_unsigned(76,8) ,
9832	 => std_logic_vector(to_unsigned(74,8) ,
9833	 => std_logic_vector(to_unsigned(74,8) ,
9834	 => std_logic_vector(to_unsigned(67,8) ,
9835	 => std_logic_vector(to_unsigned(72,8) ,
9836	 => std_logic_vector(to_unsigned(54,8) ,
9837	 => std_logic_vector(to_unsigned(49,8) ,
9838	 => std_logic_vector(to_unsigned(52,8) ,
9839	 => std_logic_vector(to_unsigned(63,8) ,
9840	 => std_logic_vector(to_unsigned(82,8) ,
9841	 => std_logic_vector(to_unsigned(80,8) ,
9842	 => std_logic_vector(to_unsigned(15,8) ,
9843	 => std_logic_vector(to_unsigned(0,8) ,
9844	 => std_logic_vector(to_unsigned(0,8) ,
9845	 => std_logic_vector(to_unsigned(6,8) ,
9846	 => std_logic_vector(to_unsigned(66,8) ,
9847	 => std_logic_vector(to_unsigned(82,8) ,
9848	 => std_logic_vector(to_unsigned(97,8) ,
9849	 => std_logic_vector(to_unsigned(107,8) ,
9850	 => std_logic_vector(to_unsigned(103,8) ,
9851	 => std_logic_vector(to_unsigned(103,8) ,
9852	 => std_logic_vector(to_unsigned(101,8) ,
9853	 => std_logic_vector(to_unsigned(85,8) ,
9854	 => std_logic_vector(to_unsigned(78,8) ,
9855	 => std_logic_vector(to_unsigned(93,8) ,
9856	 => std_logic_vector(to_unsigned(84,8) ,
9857	 => std_logic_vector(to_unsigned(68,8) ,
9858	 => std_logic_vector(to_unsigned(74,8) ,
9859	 => std_logic_vector(to_unsigned(82,8) ,
9860	 => std_logic_vector(to_unsigned(70,8) ,
9861	 => std_logic_vector(to_unsigned(87,8) ,
9862	 => std_logic_vector(to_unsigned(107,8) ,
9863	 => std_logic_vector(to_unsigned(95,8) ,
9864	 => std_logic_vector(to_unsigned(71,8) ,
9865	 => std_logic_vector(to_unsigned(84,8) ,
9866	 => std_logic_vector(to_unsigned(90,8) ,
9867	 => std_logic_vector(to_unsigned(95,8) ,
9868	 => std_logic_vector(to_unsigned(96,8) ,
9869	 => std_logic_vector(to_unsigned(82,8) ,
9870	 => std_logic_vector(to_unsigned(78,8) ,
9871	 => std_logic_vector(to_unsigned(93,8) ,
9872	 => std_logic_vector(to_unsigned(92,8) ,
9873	 => std_logic_vector(to_unsigned(79,8) ,
9874	 => std_logic_vector(to_unsigned(74,8) ,
9875	 => std_logic_vector(to_unsigned(77,8) ,
9876	 => std_logic_vector(to_unsigned(82,8) ,
9877	 => std_logic_vector(to_unsigned(82,8) ,
9878	 => std_logic_vector(to_unsigned(86,8) ,
9879	 => std_logic_vector(to_unsigned(90,8) ,
9880	 => std_logic_vector(to_unsigned(90,8) ,
9881	 => std_logic_vector(to_unsigned(87,8) ,
9882	 => std_logic_vector(to_unsigned(85,8) ,
9883	 => std_logic_vector(to_unsigned(87,8) ,
9884	 => std_logic_vector(to_unsigned(88,8) ,
9885	 => std_logic_vector(to_unsigned(87,8) ,
9886	 => std_logic_vector(to_unsigned(92,8) ,
9887	 => std_logic_vector(to_unsigned(95,8) ,
9888	 => std_logic_vector(to_unsigned(92,8) ,
9889	 => std_logic_vector(to_unsigned(91,8) ,
9890	 => std_logic_vector(to_unsigned(97,8) ,
9891	 => std_logic_vector(to_unsigned(101,8) ,
9892	 => std_logic_vector(to_unsigned(105,8) ,
9893	 => std_logic_vector(to_unsigned(105,8) ,
9894	 => std_logic_vector(to_unsigned(107,8) ,
9895	 => std_logic_vector(to_unsigned(109,8) ,
9896	 => std_logic_vector(to_unsigned(105,8) ,
9897	 => std_logic_vector(to_unsigned(111,8) ,
9898	 => std_logic_vector(to_unsigned(115,8) ,
9899	 => std_logic_vector(to_unsigned(121,8) ,
9900	 => std_logic_vector(to_unsigned(125,8) ,
9901	 => std_logic_vector(to_unsigned(125,8) ,
9902	 => std_logic_vector(to_unsigned(127,8) ,
9903	 => std_logic_vector(to_unsigned(127,8) ,
9904	 => std_logic_vector(to_unsigned(134,8) ,
9905	 => std_logic_vector(to_unsigned(138,8) ,
9906	 => std_logic_vector(to_unsigned(136,8) ,
9907	 => std_logic_vector(to_unsigned(144,8) ,
9908	 => std_logic_vector(to_unsigned(146,8) ,
9909	 => std_logic_vector(to_unsigned(149,8) ,
9910	 => std_logic_vector(to_unsigned(152,8) ,
9911	 => std_logic_vector(to_unsigned(154,8) ,
9912	 => std_logic_vector(to_unsigned(151,8) ,
9913	 => std_logic_vector(to_unsigned(152,8) ,
9914	 => std_logic_vector(to_unsigned(154,8) ,
9915	 => std_logic_vector(to_unsigned(154,8) ,
9916	 => std_logic_vector(to_unsigned(156,8) ,
9917	 => std_logic_vector(to_unsigned(154,8) ,
9918	 => std_logic_vector(to_unsigned(152,8) ,
9919	 => std_logic_vector(to_unsigned(151,8) ,
9920	 => std_logic_vector(to_unsigned(152,8) ,
9921	 => std_logic_vector(to_unsigned(109,8) ,
9922	 => std_logic_vector(to_unsigned(107,8) ,
9923	 => std_logic_vector(to_unsigned(101,8) ,
9924	 => std_logic_vector(to_unsigned(100,8) ,
9925	 => std_logic_vector(to_unsigned(103,8) ,
9926	 => std_logic_vector(to_unsigned(99,8) ,
9927	 => std_logic_vector(to_unsigned(95,8) ,
9928	 => std_logic_vector(to_unsigned(104,8) ,
9929	 => std_logic_vector(to_unsigned(112,8) ,
9930	 => std_logic_vector(to_unsigned(101,8) ,
9931	 => std_logic_vector(to_unsigned(93,8) ,
9932	 => std_logic_vector(to_unsigned(92,8) ,
9933	 => std_logic_vector(to_unsigned(92,8) ,
9934	 => std_logic_vector(to_unsigned(95,8) ,
9935	 => std_logic_vector(to_unsigned(96,8) ,
9936	 => std_logic_vector(to_unsigned(97,8) ,
9937	 => std_logic_vector(to_unsigned(99,8) ,
9938	 => std_logic_vector(to_unsigned(95,8) ,
9939	 => std_logic_vector(to_unsigned(92,8) ,
9940	 => std_logic_vector(to_unsigned(93,8) ,
9941	 => std_logic_vector(to_unsigned(97,8) ,
9942	 => std_logic_vector(to_unsigned(97,8) ,
9943	 => std_logic_vector(to_unsigned(100,8) ,
9944	 => std_logic_vector(to_unsigned(96,8) ,
9945	 => std_logic_vector(to_unsigned(95,8) ,
9946	 => std_logic_vector(to_unsigned(96,8) ,
9947	 => std_logic_vector(to_unsigned(108,8) ,
9948	 => std_logic_vector(to_unsigned(114,8) ,
9949	 => std_logic_vector(to_unsigned(107,8) ,
9950	 => std_logic_vector(to_unsigned(107,8) ,
9951	 => std_logic_vector(to_unsigned(108,8) ,
9952	 => std_logic_vector(to_unsigned(107,8) ,
9953	 => std_logic_vector(to_unsigned(103,8) ,
9954	 => std_logic_vector(to_unsigned(100,8) ,
9955	 => std_logic_vector(to_unsigned(105,8) ,
9956	 => std_logic_vector(to_unsigned(103,8) ,
9957	 => std_logic_vector(to_unsigned(97,8) ,
9958	 => std_logic_vector(to_unsigned(100,8) ,
9959	 => std_logic_vector(to_unsigned(97,8) ,
9960	 => std_logic_vector(to_unsigned(100,8) ,
9961	 => std_logic_vector(to_unsigned(108,8) ,
9962	 => std_logic_vector(to_unsigned(114,8) ,
9963	 => std_logic_vector(to_unsigned(107,8) ,
9964	 => std_logic_vector(to_unsigned(107,8) ,
9965	 => std_logic_vector(to_unsigned(119,8) ,
9966	 => std_logic_vector(to_unsigned(118,8) ,
9967	 => std_logic_vector(to_unsigned(115,8) ,
9968	 => std_logic_vector(to_unsigned(119,8) ,
9969	 => std_logic_vector(to_unsigned(124,8) ,
9970	 => std_logic_vector(to_unsigned(121,8) ,
9971	 => std_logic_vector(to_unsigned(119,8) ,
9972	 => std_logic_vector(to_unsigned(124,8) ,
9973	 => std_logic_vector(to_unsigned(128,8) ,
9974	 => std_logic_vector(to_unsigned(124,8) ,
9975	 => std_logic_vector(to_unsigned(124,8) ,
9976	 => std_logic_vector(to_unsigned(128,8) ,
9977	 => std_logic_vector(to_unsigned(125,8) ,
9978	 => std_logic_vector(to_unsigned(128,8) ,
9979	 => std_logic_vector(to_unsigned(134,8) ,
9980	 => std_logic_vector(to_unsigned(136,8) ,
9981	 => std_logic_vector(to_unsigned(133,8) ,
9982	 => std_logic_vector(to_unsigned(138,8) ,
9983	 => std_logic_vector(to_unsigned(142,8) ,
9984	 => std_logic_vector(to_unsigned(139,8) ,
9985	 => std_logic_vector(to_unsigned(138,8) ,
9986	 => std_logic_vector(to_unsigned(131,8) ,
9987	 => std_logic_vector(to_unsigned(130,8) ,
9988	 => std_logic_vector(to_unsigned(136,8) ,
9989	 => std_logic_vector(to_unsigned(131,8) ,
9990	 => std_logic_vector(to_unsigned(133,8) ,
9991	 => std_logic_vector(to_unsigned(141,8) ,
9992	 => std_logic_vector(to_unsigned(141,8) ,
9993	 => std_logic_vector(to_unsigned(141,8) ,
9994	 => std_logic_vector(to_unsigned(146,8) ,
9995	 => std_logic_vector(to_unsigned(141,8) ,
9996	 => std_logic_vector(to_unsigned(141,8) ,
9997	 => std_logic_vector(to_unsigned(138,8) ,
9998	 => std_logic_vector(to_unsigned(134,8) ,
9999	 => std_logic_vector(to_unsigned(138,8) ,
10000	 => std_logic_vector(to_unsigned(136,8) ,
10001	 => std_logic_vector(to_unsigned(133,8) ,
10002	 => std_logic_vector(to_unsigned(131,8) ,
10003	 => std_logic_vector(to_unsigned(127,8) ,
10004	 => std_logic_vector(to_unsigned(127,8) ,
10005	 => std_logic_vector(to_unsigned(134,8) ,
10006	 => std_logic_vector(to_unsigned(133,8) ,
10007	 => std_logic_vector(to_unsigned(138,8) ,
10008	 => std_logic_vector(to_unsigned(138,8) ,
10009	 => std_logic_vector(to_unsigned(133,8) ,
10010	 => std_logic_vector(to_unsigned(134,8) ,
10011	 => std_logic_vector(to_unsigned(131,8) ,
10012	 => std_logic_vector(to_unsigned(134,8) ,
10013	 => std_logic_vector(to_unsigned(133,8) ,
10014	 => std_logic_vector(to_unsigned(122,8) ,
10015	 => std_logic_vector(to_unsigned(127,8) ,
10016	 => std_logic_vector(to_unsigned(124,8) ,
10017	 => std_logic_vector(to_unsigned(119,8) ,
10018	 => std_logic_vector(to_unsigned(122,8) ,
10019	 => std_logic_vector(to_unsigned(115,8) ,
10020	 => std_logic_vector(to_unsigned(109,8) ,
10021	 => std_logic_vector(to_unsigned(114,8) ,
10022	 => std_logic_vector(to_unsigned(104,8) ,
10023	 => std_logic_vector(to_unsigned(72,8) ,
10024	 => std_logic_vector(to_unsigned(88,8) ,
10025	 => std_logic_vector(to_unsigned(92,8) ,
10026	 => std_logic_vector(to_unsigned(72,8) ,
10027	 => std_logic_vector(to_unsigned(76,8) ,
10028	 => std_logic_vector(to_unsigned(67,8) ,
10029	 => std_logic_vector(to_unsigned(61,8) ,
10030	 => std_logic_vector(to_unsigned(66,8) ,
10031	 => std_logic_vector(to_unsigned(64,8) ,
10032	 => std_logic_vector(to_unsigned(65,8) ,
10033	 => std_logic_vector(to_unsigned(68,8) ,
10034	 => std_logic_vector(to_unsigned(72,8) ,
10035	 => std_logic_vector(to_unsigned(68,8) ,
10036	 => std_logic_vector(to_unsigned(66,8) ,
10037	 => std_logic_vector(to_unsigned(69,8) ,
10038	 => std_logic_vector(to_unsigned(80,8) ,
10039	 => std_logic_vector(to_unsigned(85,8) ,
10040	 => std_logic_vector(to_unsigned(85,8) ,
10041	 => std_logic_vector(to_unsigned(85,8) ,
10042	 => std_logic_vector(to_unsigned(96,8) ,
10043	 => std_logic_vector(to_unsigned(100,8) ,
10044	 => std_logic_vector(to_unsigned(97,8) ,
10045	 => std_logic_vector(to_unsigned(109,8) ,
10046	 => std_logic_vector(to_unsigned(114,8) ,
10047	 => std_logic_vector(to_unsigned(95,8) ,
10048	 => std_logic_vector(to_unsigned(96,8) ,
10049	 => std_logic_vector(to_unsigned(101,8) ,
10050	 => std_logic_vector(to_unsigned(100,8) ,
10051	 => std_logic_vector(to_unsigned(103,8) ,
10052	 => std_logic_vector(to_unsigned(100,8) ,
10053	 => std_logic_vector(to_unsigned(93,8) ,
10054	 => std_logic_vector(to_unsigned(96,8) ,
10055	 => std_logic_vector(to_unsigned(101,8) ,
10056	 => std_logic_vector(to_unsigned(104,8) ,
10057	 => std_logic_vector(to_unsigned(96,8) ,
10058	 => std_logic_vector(to_unsigned(97,8) ,
10059	 => std_logic_vector(to_unsigned(91,8) ,
10060	 => std_logic_vector(to_unsigned(100,8) ,
10061	 => std_logic_vector(to_unsigned(112,8) ,
10062	 => std_logic_vector(to_unsigned(99,8) ,
10063	 => std_logic_vector(to_unsigned(93,8) ,
10064	 => std_logic_vector(to_unsigned(114,8) ,
10065	 => std_logic_vector(to_unsigned(122,8) ,
10066	 => std_logic_vector(to_unsigned(119,8) ,
10067	 => std_logic_vector(to_unsigned(114,8) ,
10068	 => std_logic_vector(to_unsigned(101,8) ,
10069	 => std_logic_vector(to_unsigned(92,8) ,
10070	 => std_logic_vector(to_unsigned(84,8) ,
10071	 => std_logic_vector(to_unsigned(80,8) ,
10072	 => std_logic_vector(to_unsigned(82,8) ,
10073	 => std_logic_vector(to_unsigned(85,8) ,
10074	 => std_logic_vector(to_unsigned(92,8) ,
10075	 => std_logic_vector(to_unsigned(90,8) ,
10076	 => std_logic_vector(to_unsigned(81,8) ,
10077	 => std_logic_vector(to_unsigned(84,8) ,
10078	 => std_logic_vector(to_unsigned(81,8) ,
10079	 => std_logic_vector(to_unsigned(84,8) ,
10080	 => std_logic_vector(to_unsigned(93,8) ,
10081	 => std_logic_vector(to_unsigned(84,8) ,
10082	 => std_logic_vector(to_unsigned(76,8) ,
10083	 => std_logic_vector(to_unsigned(84,8) ,
10084	 => std_logic_vector(to_unsigned(91,8) ,
10085	 => std_logic_vector(to_unsigned(82,8) ,
10086	 => std_logic_vector(to_unsigned(80,8) ,
10087	 => std_logic_vector(to_unsigned(80,8) ,
10088	 => std_logic_vector(to_unsigned(78,8) ,
10089	 => std_logic_vector(to_unsigned(80,8) ,
10090	 => std_logic_vector(to_unsigned(81,8) ,
10091	 => std_logic_vector(to_unsigned(85,8) ,
10092	 => std_logic_vector(to_unsigned(88,8) ,
10093	 => std_logic_vector(to_unsigned(87,8) ,
10094	 => std_logic_vector(to_unsigned(85,8) ,
10095	 => std_logic_vector(to_unsigned(90,8) ,
10096	 => std_logic_vector(to_unsigned(93,8) ,
10097	 => std_logic_vector(to_unsigned(100,8) ,
10098	 => std_logic_vector(to_unsigned(96,8) ,
10099	 => std_logic_vector(to_unsigned(87,8) ,
10100	 => std_logic_vector(to_unsigned(95,8) ,
10101	 => std_logic_vector(to_unsigned(92,8) ,
10102	 => std_logic_vector(to_unsigned(82,8) ,
10103	 => std_logic_vector(to_unsigned(77,8) ,
10104	 => std_logic_vector(to_unsigned(91,8) ,
10105	 => std_logic_vector(to_unsigned(92,8) ,
10106	 => std_logic_vector(to_unsigned(92,8) ,
10107	 => std_logic_vector(to_unsigned(99,8) ,
10108	 => std_logic_vector(to_unsigned(97,8) ,
10109	 => std_logic_vector(to_unsigned(93,8) ,
10110	 => std_logic_vector(to_unsigned(96,8) ,
10111	 => std_logic_vector(to_unsigned(97,8) ,
10112	 => std_logic_vector(to_unsigned(104,8) ,
10113	 => std_logic_vector(to_unsigned(91,8) ,
10114	 => std_logic_vector(to_unsigned(80,8) ,
10115	 => std_logic_vector(to_unsigned(95,8) ,
10116	 => std_logic_vector(to_unsigned(101,8) ,
10117	 => std_logic_vector(to_unsigned(86,8) ,
10118	 => std_logic_vector(to_unsigned(86,8) ,
10119	 => std_logic_vector(to_unsigned(81,8) ,
10120	 => std_logic_vector(to_unsigned(79,8) ,
10121	 => std_logic_vector(to_unsigned(96,8) ,
10122	 => std_logic_vector(to_unsigned(88,8) ,
10123	 => std_logic_vector(to_unsigned(92,8) ,
10124	 => std_logic_vector(to_unsigned(90,8) ,
10125	 => std_logic_vector(to_unsigned(80,8) ,
10126	 => std_logic_vector(to_unsigned(81,8) ,
10127	 => std_logic_vector(to_unsigned(85,8) ,
10128	 => std_logic_vector(to_unsigned(85,8) ,
10129	 => std_logic_vector(to_unsigned(87,8) ,
10130	 => std_logic_vector(to_unsigned(86,8) ,
10131	 => std_logic_vector(to_unsigned(73,8) ,
10132	 => std_logic_vector(to_unsigned(65,8) ,
10133	 => std_logic_vector(to_unsigned(63,8) ,
10134	 => std_logic_vector(to_unsigned(62,8) ,
10135	 => std_logic_vector(to_unsigned(62,8) ,
10136	 => std_logic_vector(to_unsigned(65,8) ,
10137	 => std_logic_vector(to_unsigned(61,8) ,
10138	 => std_logic_vector(to_unsigned(68,8) ,
10139	 => std_logic_vector(to_unsigned(81,8) ,
10140	 => std_logic_vector(to_unsigned(72,8) ,
10141	 => std_logic_vector(to_unsigned(67,8) ,
10142	 => std_logic_vector(to_unsigned(85,8) ,
10143	 => std_logic_vector(to_unsigned(90,8) ,
10144	 => std_logic_vector(to_unsigned(84,8) ,
10145	 => std_logic_vector(to_unsigned(68,8) ,
10146	 => std_logic_vector(to_unsigned(81,8) ,
10147	 => std_logic_vector(to_unsigned(64,8) ,
10148	 => std_logic_vector(to_unsigned(53,8) ,
10149	 => std_logic_vector(to_unsigned(61,8) ,
10150	 => std_logic_vector(to_unsigned(70,8) ,
10151	 => std_logic_vector(to_unsigned(73,8) ,
10152	 => std_logic_vector(to_unsigned(80,8) ,
10153	 => std_logic_vector(to_unsigned(74,8) ,
10154	 => std_logic_vector(to_unsigned(65,8) ,
10155	 => std_logic_vector(to_unsigned(68,8) ,
10156	 => std_logic_vector(to_unsigned(54,8) ,
10157	 => std_logic_vector(to_unsigned(52,8) ,
10158	 => std_logic_vector(to_unsigned(62,8) ,
10159	 => std_logic_vector(to_unsigned(63,8) ,
10160	 => std_logic_vector(to_unsigned(67,8) ,
10161	 => std_logic_vector(to_unsigned(76,8) ,
10162	 => std_logic_vector(to_unsigned(18,8) ,
10163	 => std_logic_vector(to_unsigned(0,8) ,
10164	 => std_logic_vector(to_unsigned(0,8) ,
10165	 => std_logic_vector(to_unsigned(3,8) ,
10166	 => std_logic_vector(to_unsigned(51,8) ,
10167	 => std_logic_vector(to_unsigned(86,8) ,
10168	 => std_logic_vector(to_unsigned(82,8) ,
10169	 => std_logic_vector(to_unsigned(76,8) ,
10170	 => std_logic_vector(to_unsigned(97,8) ,
10171	 => std_logic_vector(to_unsigned(112,8) ,
10172	 => std_logic_vector(to_unsigned(99,8) ,
10173	 => std_logic_vector(to_unsigned(88,8) ,
10174	 => std_logic_vector(to_unsigned(81,8) ,
10175	 => std_logic_vector(to_unsigned(96,8) ,
10176	 => std_logic_vector(to_unsigned(80,8) ,
10177	 => std_logic_vector(to_unsigned(70,8) ,
10178	 => std_logic_vector(to_unsigned(78,8) ,
10179	 => std_logic_vector(to_unsigned(62,8) ,
10180	 => std_logic_vector(to_unsigned(59,8) ,
10181	 => std_logic_vector(to_unsigned(84,8) ,
10182	 => std_logic_vector(to_unsigned(104,8) ,
10183	 => std_logic_vector(to_unsigned(88,8) ,
10184	 => std_logic_vector(to_unsigned(69,8) ,
10185	 => std_logic_vector(to_unsigned(86,8) ,
10186	 => std_logic_vector(to_unsigned(92,8) ,
10187	 => std_logic_vector(to_unsigned(91,8) ,
10188	 => std_logic_vector(to_unsigned(93,8) ,
10189	 => std_logic_vector(to_unsigned(84,8) ,
10190	 => std_logic_vector(to_unsigned(71,8) ,
10191	 => std_logic_vector(to_unsigned(73,8) ,
10192	 => std_logic_vector(to_unsigned(73,8) ,
10193	 => std_logic_vector(to_unsigned(64,8) ,
10194	 => std_logic_vector(to_unsigned(63,8) ,
10195	 => std_logic_vector(to_unsigned(77,8) ,
10196	 => std_logic_vector(to_unsigned(81,8) ,
10197	 => std_logic_vector(to_unsigned(79,8) ,
10198	 => std_logic_vector(to_unsigned(79,8) ,
10199	 => std_logic_vector(to_unsigned(84,8) ,
10200	 => std_logic_vector(to_unsigned(82,8) ,
10201	 => std_logic_vector(to_unsigned(84,8) ,
10202	 => std_logic_vector(to_unsigned(86,8) ,
10203	 => std_logic_vector(to_unsigned(87,8) ,
10204	 => std_logic_vector(to_unsigned(90,8) ,
10205	 => std_logic_vector(to_unsigned(92,8) ,
10206	 => std_logic_vector(to_unsigned(96,8) ,
10207	 => std_logic_vector(to_unsigned(96,8) ,
10208	 => std_logic_vector(to_unsigned(92,8) ,
10209	 => std_logic_vector(to_unsigned(99,8) ,
10210	 => std_logic_vector(to_unsigned(108,8) ,
10211	 => std_logic_vector(to_unsigned(108,8) ,
10212	 => std_logic_vector(to_unsigned(105,8) ,
10213	 => std_logic_vector(to_unsigned(107,8) ,
10214	 => std_logic_vector(to_unsigned(109,8) ,
10215	 => std_logic_vector(to_unsigned(109,8) ,
10216	 => std_logic_vector(to_unsigned(105,8) ,
10217	 => std_logic_vector(to_unsigned(107,8) ,
10218	 => std_logic_vector(to_unsigned(111,8) ,
10219	 => std_logic_vector(to_unsigned(124,8) ,
10220	 => std_logic_vector(to_unsigned(131,8) ,
10221	 => std_logic_vector(to_unsigned(127,8) ,
10222	 => std_logic_vector(to_unsigned(128,8) ,
10223	 => std_logic_vector(to_unsigned(131,8) ,
10224	 => std_logic_vector(to_unsigned(136,8) ,
10225	 => std_logic_vector(to_unsigned(141,8) ,
10226	 => std_logic_vector(to_unsigned(139,8) ,
10227	 => std_logic_vector(to_unsigned(139,8) ,
10228	 => std_logic_vector(to_unsigned(141,8) ,
10229	 => std_logic_vector(to_unsigned(144,8) ,
10230	 => std_logic_vector(to_unsigned(147,8) ,
10231	 => std_logic_vector(to_unsigned(151,8) ,
10232	 => std_logic_vector(to_unsigned(157,8) ,
10233	 => std_logic_vector(to_unsigned(157,8) ,
10234	 => std_logic_vector(to_unsigned(154,8) ,
10235	 => std_logic_vector(to_unsigned(151,8) ,
10236	 => std_logic_vector(to_unsigned(154,8) ,
10237	 => std_logic_vector(to_unsigned(156,8) ,
10238	 => std_logic_vector(to_unsigned(152,8) ,
10239	 => std_logic_vector(to_unsigned(149,8) ,
10240	 => std_logic_vector(to_unsigned(149,8) ,
10241	 => std_logic_vector(to_unsigned(107,8) ,
10242	 => std_logic_vector(to_unsigned(104,8) ,
10243	 => std_logic_vector(to_unsigned(100,8) ,
10244	 => std_logic_vector(to_unsigned(101,8) ,
10245	 => std_logic_vector(to_unsigned(103,8) ,
10246	 => std_logic_vector(to_unsigned(101,8) ,
10247	 => std_logic_vector(to_unsigned(107,8) ,
10248	 => std_logic_vector(to_unsigned(114,8) ,
10249	 => std_logic_vector(to_unsigned(119,8) ,
10250	 => std_logic_vector(to_unsigned(111,8) ,
10251	 => std_logic_vector(to_unsigned(101,8) ,
10252	 => std_logic_vector(to_unsigned(97,8) ,
10253	 => std_logic_vector(to_unsigned(101,8) ,
10254	 => std_logic_vector(to_unsigned(104,8) ,
10255	 => std_logic_vector(to_unsigned(104,8) ,
10256	 => std_logic_vector(to_unsigned(115,8) ,
10257	 => std_logic_vector(to_unsigned(119,8) ,
10258	 => std_logic_vector(to_unsigned(105,8) ,
10259	 => std_logic_vector(to_unsigned(99,8) ,
10260	 => std_logic_vector(to_unsigned(100,8) ,
10261	 => std_logic_vector(to_unsigned(99,8) ,
10262	 => std_logic_vector(to_unsigned(97,8) ,
10263	 => std_logic_vector(to_unsigned(105,8) ,
10264	 => std_logic_vector(to_unsigned(111,8) ,
10265	 => std_logic_vector(to_unsigned(105,8) ,
10266	 => std_logic_vector(to_unsigned(104,8) ,
10267	 => std_logic_vector(to_unsigned(104,8) ,
10268	 => std_logic_vector(to_unsigned(108,8) ,
10269	 => std_logic_vector(to_unsigned(109,8) ,
10270	 => std_logic_vector(to_unsigned(115,8) ,
10271	 => std_logic_vector(to_unsigned(114,8) ,
10272	 => std_logic_vector(to_unsigned(112,8) ,
10273	 => std_logic_vector(to_unsigned(111,8) ,
10274	 => std_logic_vector(to_unsigned(111,8) ,
10275	 => std_logic_vector(to_unsigned(118,8) ,
10276	 => std_logic_vector(to_unsigned(114,8) ,
10277	 => std_logic_vector(to_unsigned(107,8) ,
10278	 => std_logic_vector(to_unsigned(115,8) ,
10279	 => std_logic_vector(to_unsigned(118,8) ,
10280	 => std_logic_vector(to_unsigned(116,8) ,
10281	 => std_logic_vector(to_unsigned(114,8) ,
10282	 => std_logic_vector(to_unsigned(112,8) ,
10283	 => std_logic_vector(to_unsigned(112,8) ,
10284	 => std_logic_vector(to_unsigned(115,8) ,
10285	 => std_logic_vector(to_unsigned(124,8) ,
10286	 => std_logic_vector(to_unsigned(119,8) ,
10287	 => std_logic_vector(to_unsigned(118,8) ,
10288	 => std_logic_vector(to_unsigned(124,8) ,
10289	 => std_logic_vector(to_unsigned(127,8) ,
10290	 => std_logic_vector(to_unsigned(124,8) ,
10291	 => std_logic_vector(to_unsigned(124,8) ,
10292	 => std_logic_vector(to_unsigned(124,8) ,
10293	 => std_logic_vector(to_unsigned(125,8) ,
10294	 => std_logic_vector(to_unsigned(124,8) ,
10295	 => std_logic_vector(to_unsigned(130,8) ,
10296	 => std_logic_vector(to_unsigned(138,8) ,
10297	 => std_logic_vector(to_unsigned(131,8) ,
10298	 => std_logic_vector(to_unsigned(133,8) ,
10299	 => std_logic_vector(to_unsigned(138,8) ,
10300	 => std_logic_vector(to_unsigned(142,8) ,
10301	 => std_logic_vector(to_unsigned(141,8) ,
10302	 => std_logic_vector(to_unsigned(141,8) ,
10303	 => std_logic_vector(to_unsigned(144,8) ,
10304	 => std_logic_vector(to_unsigned(138,8) ,
10305	 => std_logic_vector(to_unsigned(142,8) ,
10306	 => std_logic_vector(to_unsigned(136,8) ,
10307	 => std_logic_vector(to_unsigned(131,8) ,
10308	 => std_logic_vector(to_unsigned(138,8) ,
10309	 => std_logic_vector(to_unsigned(138,8) ,
10310	 => std_logic_vector(to_unsigned(139,8) ,
10311	 => std_logic_vector(to_unsigned(141,8) ,
10312	 => std_logic_vector(to_unsigned(139,8) ,
10313	 => std_logic_vector(to_unsigned(144,8) ,
10314	 => std_logic_vector(to_unsigned(147,8) ,
10315	 => std_logic_vector(to_unsigned(138,8) ,
10316	 => std_logic_vector(to_unsigned(141,8) ,
10317	 => std_logic_vector(to_unsigned(139,8) ,
10318	 => std_logic_vector(to_unsigned(134,8) ,
10319	 => std_logic_vector(to_unsigned(139,8) ,
10320	 => std_logic_vector(to_unsigned(136,8) ,
10321	 => std_logic_vector(to_unsigned(131,8) ,
10322	 => std_logic_vector(to_unsigned(130,8) ,
10323	 => std_logic_vector(to_unsigned(133,8) ,
10324	 => std_logic_vector(to_unsigned(134,8) ,
10325	 => std_logic_vector(to_unsigned(138,8) ,
10326	 => std_logic_vector(to_unsigned(134,8) ,
10327	 => std_logic_vector(to_unsigned(141,8) ,
10328	 => std_logic_vector(to_unsigned(142,8) ,
10329	 => std_logic_vector(to_unsigned(138,8) ,
10330	 => std_logic_vector(to_unsigned(141,8) ,
10331	 => std_logic_vector(to_unsigned(134,8) ,
10332	 => std_logic_vector(to_unsigned(131,8) ,
10333	 => std_logic_vector(to_unsigned(125,8) ,
10334	 => std_logic_vector(to_unsigned(107,8) ,
10335	 => std_logic_vector(to_unsigned(114,8) ,
10336	 => std_logic_vector(to_unsigned(109,8) ,
10337	 => std_logic_vector(to_unsigned(118,8) ,
10338	 => std_logic_vector(to_unsigned(124,8) ,
10339	 => std_logic_vector(to_unsigned(122,8) ,
10340	 => std_logic_vector(to_unsigned(115,8) ,
10341	 => std_logic_vector(to_unsigned(118,8) ,
10342	 => std_logic_vector(to_unsigned(108,8) ,
10343	 => std_logic_vector(to_unsigned(82,8) ,
10344	 => std_logic_vector(to_unsigned(85,8) ,
10345	 => std_logic_vector(to_unsigned(86,8) ,
10346	 => std_logic_vector(to_unsigned(70,8) ,
10347	 => std_logic_vector(to_unsigned(66,8) ,
10348	 => std_logic_vector(to_unsigned(66,8) ,
10349	 => std_logic_vector(to_unsigned(72,8) ,
10350	 => std_logic_vector(to_unsigned(76,8) ,
10351	 => std_logic_vector(to_unsigned(67,8) ,
10352	 => std_logic_vector(to_unsigned(66,8) ,
10353	 => std_logic_vector(to_unsigned(68,8) ,
10354	 => std_logic_vector(to_unsigned(74,8) ,
10355	 => std_logic_vector(to_unsigned(74,8) ,
10356	 => std_logic_vector(to_unsigned(78,8) ,
10357	 => std_logic_vector(to_unsigned(76,8) ,
10358	 => std_logic_vector(to_unsigned(81,8) ,
10359	 => std_logic_vector(to_unsigned(85,8) ,
10360	 => std_logic_vector(to_unsigned(81,8) ,
10361	 => std_logic_vector(to_unsigned(79,8) ,
10362	 => std_logic_vector(to_unsigned(90,8) ,
10363	 => std_logic_vector(to_unsigned(104,8) ,
10364	 => std_logic_vector(to_unsigned(103,8) ,
10365	 => std_logic_vector(to_unsigned(100,8) ,
10366	 => std_logic_vector(to_unsigned(105,8) ,
10367	 => std_logic_vector(to_unsigned(104,8) ,
10368	 => std_logic_vector(to_unsigned(97,8) ,
10369	 => std_logic_vector(to_unsigned(103,8) ,
10370	 => std_logic_vector(to_unsigned(109,8) ,
10371	 => std_logic_vector(to_unsigned(104,8) ,
10372	 => std_logic_vector(to_unsigned(101,8) ,
10373	 => std_logic_vector(to_unsigned(103,8) ,
10374	 => std_logic_vector(to_unsigned(101,8) ,
10375	 => std_logic_vector(to_unsigned(100,8) ,
10376	 => std_logic_vector(to_unsigned(105,8) ,
10377	 => std_logic_vector(to_unsigned(103,8) ,
10378	 => std_logic_vector(to_unsigned(107,8) ,
10379	 => std_logic_vector(to_unsigned(105,8) ,
10380	 => std_logic_vector(to_unsigned(105,8) ,
10381	 => std_logic_vector(to_unsigned(108,8) ,
10382	 => std_logic_vector(to_unsigned(101,8) ,
10383	 => std_logic_vector(to_unsigned(105,8) ,
10384	 => std_logic_vector(to_unsigned(109,8) ,
10385	 => std_logic_vector(to_unsigned(105,8) ,
10386	 => std_logic_vector(to_unsigned(95,8) ,
10387	 => std_logic_vector(to_unsigned(91,8) ,
10388	 => std_logic_vector(to_unsigned(87,8) ,
10389	 => std_logic_vector(to_unsigned(91,8) ,
10390	 => std_logic_vector(to_unsigned(82,8) ,
10391	 => std_logic_vector(to_unsigned(78,8) ,
10392	 => std_logic_vector(to_unsigned(85,8) ,
10393	 => std_logic_vector(to_unsigned(90,8) ,
10394	 => std_logic_vector(to_unsigned(91,8) ,
10395	 => std_logic_vector(to_unsigned(86,8) ,
10396	 => std_logic_vector(to_unsigned(77,8) ,
10397	 => std_logic_vector(to_unsigned(80,8) ,
10398	 => std_logic_vector(to_unsigned(79,8) ,
10399	 => std_logic_vector(to_unsigned(81,8) ,
10400	 => std_logic_vector(to_unsigned(91,8) ,
10401	 => std_logic_vector(to_unsigned(92,8) ,
10402	 => std_logic_vector(to_unsigned(80,8) ,
10403	 => std_logic_vector(to_unsigned(87,8) ,
10404	 => std_logic_vector(to_unsigned(77,8) ,
10405	 => std_logic_vector(to_unsigned(45,8) ,
10406	 => std_logic_vector(to_unsigned(72,8) ,
10407	 => std_logic_vector(to_unsigned(76,8) ,
10408	 => std_logic_vector(to_unsigned(73,8) ,
10409	 => std_logic_vector(to_unsigned(84,8) ,
10410	 => std_logic_vector(to_unsigned(84,8) ,
10411	 => std_logic_vector(to_unsigned(90,8) ,
10412	 => std_logic_vector(to_unsigned(85,8) ,
10413	 => std_logic_vector(to_unsigned(88,8) ,
10414	 => std_logic_vector(to_unsigned(97,8) ,
10415	 => std_logic_vector(to_unsigned(96,8) ,
10416	 => std_logic_vector(to_unsigned(95,8) ,
10417	 => std_logic_vector(to_unsigned(99,8) ,
10418	 => std_logic_vector(to_unsigned(85,8) ,
10419	 => std_logic_vector(to_unsigned(81,8) ,
10420	 => std_logic_vector(to_unsigned(87,8) ,
10421	 => std_logic_vector(to_unsigned(88,8) ,
10422	 => std_logic_vector(to_unsigned(82,8) ,
10423	 => std_logic_vector(to_unsigned(84,8) ,
10424	 => std_logic_vector(to_unsigned(99,8) ,
10425	 => std_logic_vector(to_unsigned(104,8) ,
10426	 => std_logic_vector(to_unsigned(93,8) ,
10427	 => std_logic_vector(to_unsigned(90,8) ,
10428	 => std_logic_vector(to_unsigned(96,8) ,
10429	 => std_logic_vector(to_unsigned(92,8) ,
10430	 => std_logic_vector(to_unsigned(90,8) ,
10431	 => std_logic_vector(to_unsigned(105,8) ,
10432	 => std_logic_vector(to_unsigned(130,8) ,
10433	 => std_logic_vector(to_unsigned(95,8) ,
10434	 => std_logic_vector(to_unsigned(78,8) ,
10435	 => std_logic_vector(to_unsigned(91,8) ,
10436	 => std_logic_vector(to_unsigned(90,8) ,
10437	 => std_logic_vector(to_unsigned(87,8) ,
10438	 => std_logic_vector(to_unsigned(90,8) ,
10439	 => std_logic_vector(to_unsigned(99,8) ,
10440	 => std_logic_vector(to_unsigned(97,8) ,
10441	 => std_logic_vector(to_unsigned(97,8) ,
10442	 => std_logic_vector(to_unsigned(100,8) ,
10443	 => std_logic_vector(to_unsigned(95,8) ,
10444	 => std_logic_vector(to_unsigned(88,8) ,
10445	 => std_logic_vector(to_unsigned(84,8) ,
10446	 => std_logic_vector(to_unsigned(84,8) ,
10447	 => std_logic_vector(to_unsigned(85,8) ,
10448	 => std_logic_vector(to_unsigned(86,8) ,
10449	 => std_logic_vector(to_unsigned(84,8) ,
10450	 => std_logic_vector(to_unsigned(79,8) ,
10451	 => std_logic_vector(to_unsigned(70,8) ,
10452	 => std_logic_vector(to_unsigned(72,8) ,
10453	 => std_logic_vector(to_unsigned(73,8) ,
10454	 => std_logic_vector(to_unsigned(65,8) ,
10455	 => std_logic_vector(to_unsigned(70,8) ,
10456	 => std_logic_vector(to_unsigned(72,8) ,
10457	 => std_logic_vector(to_unsigned(71,8) ,
10458	 => std_logic_vector(to_unsigned(90,8) ,
10459	 => std_logic_vector(to_unsigned(95,8) ,
10460	 => std_logic_vector(to_unsigned(72,8) ,
10461	 => std_logic_vector(to_unsigned(74,8) ,
10462	 => std_logic_vector(to_unsigned(91,8) ,
10463	 => std_logic_vector(to_unsigned(96,8) ,
10464	 => std_logic_vector(to_unsigned(79,8) ,
10465	 => std_logic_vector(to_unsigned(64,8) ,
10466	 => std_logic_vector(to_unsigned(72,8) ,
10467	 => std_logic_vector(to_unsigned(70,8) ,
10468	 => std_logic_vector(to_unsigned(69,8) ,
10469	 => std_logic_vector(to_unsigned(67,8) ,
10470	 => std_logic_vector(to_unsigned(65,8) ,
10471	 => std_logic_vector(to_unsigned(59,8) ,
10472	 => std_logic_vector(to_unsigned(82,8) ,
10473	 => std_logic_vector(to_unsigned(88,8) ,
10474	 => std_logic_vector(to_unsigned(76,8) ,
10475	 => std_logic_vector(to_unsigned(69,8) ,
10476	 => std_logic_vector(to_unsigned(57,8) ,
10477	 => std_logic_vector(to_unsigned(56,8) ,
10478	 => std_logic_vector(to_unsigned(68,8) ,
10479	 => std_logic_vector(to_unsigned(51,8) ,
10480	 => std_logic_vector(to_unsigned(53,8) ,
10481	 => std_logic_vector(to_unsigned(60,8) ,
10482	 => std_logic_vector(to_unsigned(24,8) ,
10483	 => std_logic_vector(to_unsigned(1,8) ,
10484	 => std_logic_vector(to_unsigned(0,8) ,
10485	 => std_logic_vector(to_unsigned(1,8) ,
10486	 => std_logic_vector(to_unsigned(35,8) ,
10487	 => std_logic_vector(to_unsigned(66,8) ,
10488	 => std_logic_vector(to_unsigned(56,8) ,
10489	 => std_logic_vector(to_unsigned(49,8) ,
10490	 => std_logic_vector(to_unsigned(84,8) ,
10491	 => std_logic_vector(to_unsigned(109,8) ,
10492	 => std_logic_vector(to_unsigned(95,8) ,
10493	 => std_logic_vector(to_unsigned(87,8) ,
10494	 => std_logic_vector(to_unsigned(82,8) ,
10495	 => std_logic_vector(to_unsigned(91,8) ,
10496	 => std_logic_vector(to_unsigned(74,8) ,
10497	 => std_logic_vector(to_unsigned(70,8) ,
10498	 => std_logic_vector(to_unsigned(80,8) ,
10499	 => std_logic_vector(to_unsigned(70,8) ,
10500	 => std_logic_vector(to_unsigned(82,8) ,
10501	 => std_logic_vector(to_unsigned(88,8) ,
10502	 => std_logic_vector(to_unsigned(101,8) ,
10503	 => std_logic_vector(to_unsigned(88,8) ,
10504	 => std_logic_vector(to_unsigned(82,8) ,
10505	 => std_logic_vector(to_unsigned(99,8) ,
10506	 => std_logic_vector(to_unsigned(97,8) ,
10507	 => std_logic_vector(to_unsigned(90,8) ,
10508	 => std_logic_vector(to_unsigned(93,8) ,
10509	 => std_logic_vector(to_unsigned(85,8) ,
10510	 => std_logic_vector(to_unsigned(62,8) ,
10511	 => std_logic_vector(to_unsigned(65,8) ,
10512	 => std_logic_vector(to_unsigned(65,8) ,
10513	 => std_logic_vector(to_unsigned(64,8) ,
10514	 => std_logic_vector(to_unsigned(65,8) ,
10515	 => std_logic_vector(to_unsigned(71,8) ,
10516	 => std_logic_vector(to_unsigned(74,8) ,
10517	 => std_logic_vector(to_unsigned(78,8) ,
10518	 => std_logic_vector(to_unsigned(79,8) ,
10519	 => std_logic_vector(to_unsigned(79,8) ,
10520	 => std_logic_vector(to_unsigned(77,8) ,
10521	 => std_logic_vector(to_unsigned(79,8) ,
10522	 => std_logic_vector(to_unsigned(85,8) ,
10523	 => std_logic_vector(to_unsigned(85,8) ,
10524	 => std_logic_vector(to_unsigned(87,8) ,
10525	 => std_logic_vector(to_unsigned(91,8) ,
10526	 => std_logic_vector(to_unsigned(95,8) ,
10527	 => std_logic_vector(to_unsigned(95,8) ,
10528	 => std_logic_vector(to_unsigned(90,8) ,
10529	 => std_logic_vector(to_unsigned(91,8) ,
10530	 => std_logic_vector(to_unsigned(95,8) ,
10531	 => std_logic_vector(to_unsigned(100,8) ,
10532	 => std_logic_vector(to_unsigned(99,8) ,
10533	 => std_logic_vector(to_unsigned(101,8) ,
10534	 => std_logic_vector(to_unsigned(105,8) ,
10535	 => std_logic_vector(to_unsigned(105,8) ,
10536	 => std_logic_vector(to_unsigned(99,8) ,
10537	 => std_logic_vector(to_unsigned(101,8) ,
10538	 => std_logic_vector(to_unsigned(111,8) ,
10539	 => std_logic_vector(to_unsigned(116,8) ,
10540	 => std_logic_vector(to_unsigned(121,8) ,
10541	 => std_logic_vector(to_unsigned(122,8) ,
10542	 => std_logic_vector(to_unsigned(130,8) ,
10543	 => std_logic_vector(to_unsigned(136,8) ,
10544	 => std_logic_vector(to_unsigned(134,8) ,
10545	 => std_logic_vector(to_unsigned(131,8) ,
10546	 => std_logic_vector(to_unsigned(134,8) ,
10547	 => std_logic_vector(to_unsigned(139,8) ,
10548	 => std_logic_vector(to_unsigned(136,8) ,
10549	 => std_logic_vector(to_unsigned(144,8) ,
10550	 => std_logic_vector(to_unsigned(154,8) ,
10551	 => std_logic_vector(to_unsigned(149,8) ,
10552	 => std_logic_vector(to_unsigned(152,8) ,
10553	 => std_logic_vector(to_unsigned(154,8) ,
10554	 => std_logic_vector(to_unsigned(149,8) ,
10555	 => std_logic_vector(to_unsigned(146,8) ,
10556	 => std_logic_vector(to_unsigned(149,8) ,
10557	 => std_logic_vector(to_unsigned(156,8) ,
10558	 => std_logic_vector(to_unsigned(149,8) ,
10559	 => std_logic_vector(to_unsigned(146,8) ,
10560	 => std_logic_vector(to_unsigned(146,8) ,
10561	 => std_logic_vector(to_unsigned(118,8) ,
10562	 => std_logic_vector(to_unsigned(114,8) ,
10563	 => std_logic_vector(to_unsigned(103,8) ,
10564	 => std_logic_vector(to_unsigned(104,8) ,
10565	 => std_logic_vector(to_unsigned(111,8) ,
10566	 => std_logic_vector(to_unsigned(112,8) ,
10567	 => std_logic_vector(to_unsigned(111,8) ,
10568	 => std_logic_vector(to_unsigned(116,8) ,
10569	 => std_logic_vector(to_unsigned(124,8) ,
10570	 => std_logic_vector(to_unsigned(121,8) ,
10571	 => std_logic_vector(to_unsigned(118,8) ,
10572	 => std_logic_vector(to_unsigned(116,8) ,
10573	 => std_logic_vector(to_unsigned(119,8) ,
10574	 => std_logic_vector(to_unsigned(122,8) ,
10575	 => std_logic_vector(to_unsigned(125,8) ,
10576	 => std_logic_vector(to_unsigned(127,8) ,
10577	 => std_logic_vector(to_unsigned(128,8) ,
10578	 => std_logic_vector(to_unsigned(114,8) ,
10579	 => std_logic_vector(to_unsigned(109,8) ,
10580	 => std_logic_vector(to_unsigned(109,8) ,
10581	 => std_logic_vector(to_unsigned(109,8) ,
10582	 => std_logic_vector(to_unsigned(109,8) ,
10583	 => std_logic_vector(to_unsigned(118,8) ,
10584	 => std_logic_vector(to_unsigned(127,8) ,
10585	 => std_logic_vector(to_unsigned(125,8) ,
10586	 => std_logic_vector(to_unsigned(121,8) ,
10587	 => std_logic_vector(to_unsigned(111,8) ,
10588	 => std_logic_vector(to_unsigned(112,8) ,
10589	 => std_logic_vector(to_unsigned(114,8) ,
10590	 => std_logic_vector(to_unsigned(112,8) ,
10591	 => std_logic_vector(to_unsigned(116,8) ,
10592	 => std_logic_vector(to_unsigned(109,8) ,
10593	 => std_logic_vector(to_unsigned(108,8) ,
10594	 => std_logic_vector(to_unsigned(115,8) ,
10595	 => std_logic_vector(to_unsigned(121,8) ,
10596	 => std_logic_vector(to_unsigned(115,8) ,
10597	 => std_logic_vector(to_unsigned(111,8) ,
10598	 => std_logic_vector(to_unsigned(114,8) ,
10599	 => std_logic_vector(to_unsigned(118,8) ,
10600	 => std_logic_vector(to_unsigned(118,8) ,
10601	 => std_logic_vector(to_unsigned(112,8) ,
10602	 => std_logic_vector(to_unsigned(116,8) ,
10603	 => std_logic_vector(to_unsigned(131,8) ,
10604	 => std_logic_vector(to_unsigned(130,8) ,
10605	 => std_logic_vector(to_unsigned(127,8) ,
10606	 => std_logic_vector(to_unsigned(127,8) ,
10607	 => std_logic_vector(to_unsigned(122,8) ,
10608	 => std_logic_vector(to_unsigned(121,8) ,
10609	 => std_logic_vector(to_unsigned(122,8) ,
10610	 => std_logic_vector(to_unsigned(130,8) ,
10611	 => std_logic_vector(to_unsigned(130,8) ,
10612	 => std_logic_vector(to_unsigned(122,8) ,
10613	 => std_logic_vector(to_unsigned(127,8) ,
10614	 => std_logic_vector(to_unsigned(125,8) ,
10615	 => std_logic_vector(to_unsigned(127,8) ,
10616	 => std_logic_vector(to_unsigned(131,8) ,
10617	 => std_logic_vector(to_unsigned(131,8) ,
10618	 => std_logic_vector(to_unsigned(141,8) ,
10619	 => std_logic_vector(to_unsigned(142,8) ,
10620	 => std_logic_vector(to_unsigned(144,8) ,
10621	 => std_logic_vector(to_unsigned(144,8) ,
10622	 => std_logic_vector(to_unsigned(138,8) ,
10623	 => std_logic_vector(to_unsigned(141,8) ,
10624	 => std_logic_vector(to_unsigned(146,8) ,
10625	 => std_logic_vector(to_unsigned(147,8) ,
10626	 => std_logic_vector(to_unsigned(139,8) ,
10627	 => std_logic_vector(to_unsigned(138,8) ,
10628	 => std_logic_vector(to_unsigned(142,8) ,
10629	 => std_logic_vector(to_unsigned(141,8) ,
10630	 => std_logic_vector(to_unsigned(142,8) ,
10631	 => std_logic_vector(to_unsigned(142,8) ,
10632	 => std_logic_vector(to_unsigned(138,8) ,
10633	 => std_logic_vector(to_unsigned(139,8) ,
10634	 => std_logic_vector(to_unsigned(136,8) ,
10635	 => std_logic_vector(to_unsigned(124,8) ,
10636	 => std_logic_vector(to_unsigned(133,8) ,
10637	 => std_logic_vector(to_unsigned(142,8) ,
10638	 => std_logic_vector(to_unsigned(138,8) ,
10639	 => std_logic_vector(to_unsigned(133,8) ,
10640	 => std_logic_vector(to_unsigned(133,8) ,
10641	 => std_logic_vector(to_unsigned(133,8) ,
10642	 => std_logic_vector(to_unsigned(133,8) ,
10643	 => std_logic_vector(to_unsigned(134,8) ,
10644	 => std_logic_vector(to_unsigned(133,8) ,
10645	 => std_logic_vector(to_unsigned(134,8) ,
10646	 => std_logic_vector(to_unsigned(138,8) ,
10647	 => std_logic_vector(to_unsigned(139,8) ,
10648	 => std_logic_vector(to_unsigned(138,8) ,
10649	 => std_logic_vector(to_unsigned(134,8) ,
10650	 => std_logic_vector(to_unsigned(141,8) ,
10651	 => std_logic_vector(to_unsigned(144,8) ,
10652	 => std_logic_vector(to_unsigned(138,8) ,
10653	 => std_logic_vector(to_unsigned(115,8) ,
10654	 => std_logic_vector(to_unsigned(97,8) ,
10655	 => std_logic_vector(to_unsigned(104,8) ,
10656	 => std_logic_vector(to_unsigned(99,8) ,
10657	 => std_logic_vector(to_unsigned(119,8) ,
10658	 => std_logic_vector(to_unsigned(131,8) ,
10659	 => std_logic_vector(to_unsigned(131,8) ,
10660	 => std_logic_vector(to_unsigned(124,8) ,
10661	 => std_logic_vector(to_unsigned(112,8) ,
10662	 => std_logic_vector(to_unsigned(105,8) ,
10663	 => std_logic_vector(to_unsigned(109,8) ,
10664	 => std_logic_vector(to_unsigned(105,8) ,
10665	 => std_logic_vector(to_unsigned(96,8) ,
10666	 => std_logic_vector(to_unsigned(91,8) ,
10667	 => std_logic_vector(to_unsigned(74,8) ,
10668	 => std_logic_vector(to_unsigned(73,8) ,
10669	 => std_logic_vector(to_unsigned(79,8) ,
10670	 => std_logic_vector(to_unsigned(77,8) ,
10671	 => std_logic_vector(to_unsigned(69,8) ,
10672	 => std_logic_vector(to_unsigned(62,8) ,
10673	 => std_logic_vector(to_unsigned(76,8) ,
10674	 => std_logic_vector(to_unsigned(78,8) ,
10675	 => std_logic_vector(to_unsigned(76,8) ,
10676	 => std_logic_vector(to_unsigned(86,8) ,
10677	 => std_logic_vector(to_unsigned(85,8) ,
10678	 => std_logic_vector(to_unsigned(85,8) ,
10679	 => std_logic_vector(to_unsigned(81,8) ,
10680	 => std_logic_vector(to_unsigned(84,8) ,
10681	 => std_logic_vector(to_unsigned(87,8) ,
10682	 => std_logic_vector(to_unsigned(87,8) ,
10683	 => std_logic_vector(to_unsigned(96,8) ,
10684	 => std_logic_vector(to_unsigned(115,8) ,
10685	 => std_logic_vector(to_unsigned(111,8) ,
10686	 => std_logic_vector(to_unsigned(100,8) ,
10687	 => std_logic_vector(to_unsigned(115,8) ,
10688	 => std_logic_vector(to_unsigned(109,8) ,
10689	 => std_logic_vector(to_unsigned(109,8) ,
10690	 => std_logic_vector(to_unsigned(119,8) ,
10691	 => std_logic_vector(to_unsigned(109,8) ,
10692	 => std_logic_vector(to_unsigned(103,8) ,
10693	 => std_logic_vector(to_unsigned(111,8) ,
10694	 => std_logic_vector(to_unsigned(108,8) ,
10695	 => std_logic_vector(to_unsigned(100,8) ,
10696	 => std_logic_vector(to_unsigned(92,8) ,
10697	 => std_logic_vector(to_unsigned(97,8) ,
10698	 => std_logic_vector(to_unsigned(104,8) ,
10699	 => std_logic_vector(to_unsigned(103,8) ,
10700	 => std_logic_vector(to_unsigned(99,8) ,
10701	 => std_logic_vector(to_unsigned(99,8) ,
10702	 => std_logic_vector(to_unsigned(103,8) ,
10703	 => std_logic_vector(to_unsigned(100,8) ,
10704	 => std_logic_vector(to_unsigned(97,8) ,
10705	 => std_logic_vector(to_unsigned(99,8) ,
10706	 => std_logic_vector(to_unsigned(91,8) ,
10707	 => std_logic_vector(to_unsigned(95,8) ,
10708	 => std_logic_vector(to_unsigned(96,8) ,
10709	 => std_logic_vector(to_unsigned(88,8) ,
10710	 => std_logic_vector(to_unsigned(81,8) ,
10711	 => std_logic_vector(to_unsigned(80,8) ,
10712	 => std_logic_vector(to_unsigned(87,8) ,
10713	 => std_logic_vector(to_unsigned(85,8) ,
10714	 => std_logic_vector(to_unsigned(88,8) ,
10715	 => std_logic_vector(to_unsigned(85,8) ,
10716	 => std_logic_vector(to_unsigned(86,8) ,
10717	 => std_logic_vector(to_unsigned(84,8) ,
10718	 => std_logic_vector(to_unsigned(79,8) ,
10719	 => std_logic_vector(to_unsigned(74,8) ,
10720	 => std_logic_vector(to_unsigned(82,8) ,
10721	 => std_logic_vector(to_unsigned(95,8) ,
10722	 => std_logic_vector(to_unsigned(77,8) ,
10723	 => std_logic_vector(to_unsigned(77,8) ,
10724	 => std_logic_vector(to_unsigned(70,8) ,
10725	 => std_logic_vector(to_unsigned(41,8) ,
10726	 => std_logic_vector(to_unsigned(62,8) ,
10727	 => std_logic_vector(to_unsigned(76,8) ,
10728	 => std_logic_vector(to_unsigned(76,8) ,
10729	 => std_logic_vector(to_unsigned(82,8) ,
10730	 => std_logic_vector(to_unsigned(82,8) ,
10731	 => std_logic_vector(to_unsigned(88,8) ,
10732	 => std_logic_vector(to_unsigned(85,8) ,
10733	 => std_logic_vector(to_unsigned(88,8) ,
10734	 => std_logic_vector(to_unsigned(96,8) ,
10735	 => std_logic_vector(to_unsigned(88,8) ,
10736	 => std_logic_vector(to_unsigned(79,8) ,
10737	 => std_logic_vector(to_unsigned(84,8) ,
10738	 => std_logic_vector(to_unsigned(84,8) ,
10739	 => std_logic_vector(to_unsigned(81,8) ,
10740	 => std_logic_vector(to_unsigned(77,8) ,
10741	 => std_logic_vector(to_unsigned(82,8) ,
10742	 => std_logic_vector(to_unsigned(85,8) ,
10743	 => std_logic_vector(to_unsigned(79,8) ,
10744	 => std_logic_vector(to_unsigned(87,8) ,
10745	 => std_logic_vector(to_unsigned(99,8) ,
10746	 => std_logic_vector(to_unsigned(95,8) ,
10747	 => std_logic_vector(to_unsigned(88,8) ,
10748	 => std_logic_vector(to_unsigned(100,8) ,
10749	 => std_logic_vector(to_unsigned(97,8) ,
10750	 => std_logic_vector(to_unsigned(91,8) ,
10751	 => std_logic_vector(to_unsigned(95,8) ,
10752	 => std_logic_vector(to_unsigned(125,8) ,
10753	 => std_logic_vector(to_unsigned(93,8) ,
10754	 => std_logic_vector(to_unsigned(74,8) ,
10755	 => std_logic_vector(to_unsigned(95,8) ,
10756	 => std_logic_vector(to_unsigned(90,8) ,
10757	 => std_logic_vector(to_unsigned(82,8) ,
10758	 => std_logic_vector(to_unsigned(88,8) ,
10759	 => std_logic_vector(to_unsigned(99,8) ,
10760	 => std_logic_vector(to_unsigned(107,8) ,
10761	 => std_logic_vector(to_unsigned(100,8) ,
10762	 => std_logic_vector(to_unsigned(92,8) ,
10763	 => std_logic_vector(to_unsigned(82,8) ,
10764	 => std_logic_vector(to_unsigned(78,8) ,
10765	 => std_logic_vector(to_unsigned(85,8) ,
10766	 => std_logic_vector(to_unsigned(86,8) ,
10767	 => std_logic_vector(to_unsigned(82,8) ,
10768	 => std_logic_vector(to_unsigned(80,8) ,
10769	 => std_logic_vector(to_unsigned(81,8) ,
10770	 => std_logic_vector(to_unsigned(85,8) ,
10771	 => std_logic_vector(to_unsigned(78,8) ,
10772	 => std_logic_vector(to_unsigned(76,8) ,
10773	 => std_logic_vector(to_unsigned(71,8) ,
10774	 => std_logic_vector(to_unsigned(64,8) ,
10775	 => std_logic_vector(to_unsigned(69,8) ,
10776	 => std_logic_vector(to_unsigned(74,8) ,
10777	 => std_logic_vector(to_unsigned(84,8) ,
10778	 => std_logic_vector(to_unsigned(90,8) ,
10779	 => std_logic_vector(to_unsigned(93,8) ,
10780	 => std_logic_vector(to_unsigned(82,8) ,
10781	 => std_logic_vector(to_unsigned(78,8) ,
10782	 => std_logic_vector(to_unsigned(87,8) ,
10783	 => std_logic_vector(to_unsigned(91,8) ,
10784	 => std_logic_vector(to_unsigned(81,8) ,
10785	 => std_logic_vector(to_unsigned(70,8) ,
10786	 => std_logic_vector(to_unsigned(76,8) ,
10787	 => std_logic_vector(to_unsigned(86,8) ,
10788	 => std_logic_vector(to_unsigned(80,8) ,
10789	 => std_logic_vector(to_unsigned(76,8) ,
10790	 => std_logic_vector(to_unsigned(74,8) ,
10791	 => std_logic_vector(to_unsigned(77,8) ,
10792	 => std_logic_vector(to_unsigned(81,8) ,
10793	 => std_logic_vector(to_unsigned(81,8) ,
10794	 => std_logic_vector(to_unsigned(78,8) ,
10795	 => std_logic_vector(to_unsigned(74,8) ,
10796	 => std_logic_vector(to_unsigned(62,8) ,
10797	 => std_logic_vector(to_unsigned(52,8) ,
10798	 => std_logic_vector(to_unsigned(52,8) ,
10799	 => std_logic_vector(to_unsigned(58,8) ,
10800	 => std_logic_vector(to_unsigned(61,8) ,
10801	 => std_logic_vector(to_unsigned(65,8) ,
10802	 => std_logic_vector(to_unsigned(49,8) ,
10803	 => std_logic_vector(to_unsigned(4,8) ,
10804	 => std_logic_vector(to_unsigned(0,8) ,
10805	 => std_logic_vector(to_unsigned(0,8) ,
10806	 => std_logic_vector(to_unsigned(17,8) ,
10807	 => std_logic_vector(to_unsigned(55,8) ,
10808	 => std_logic_vector(to_unsigned(50,8) ,
10809	 => std_logic_vector(to_unsigned(51,8) ,
10810	 => std_logic_vector(to_unsigned(82,8) ,
10811	 => std_logic_vector(to_unsigned(104,8) ,
10812	 => std_logic_vector(to_unsigned(101,8) ,
10813	 => std_logic_vector(to_unsigned(88,8) ,
10814	 => std_logic_vector(to_unsigned(77,8) ,
10815	 => std_logic_vector(to_unsigned(87,8) ,
10816	 => std_logic_vector(to_unsigned(84,8) ,
10817	 => std_logic_vector(to_unsigned(78,8) ,
10818	 => std_logic_vector(to_unsigned(74,8) ,
10819	 => std_logic_vector(to_unsigned(72,8) ,
10820	 => std_logic_vector(to_unsigned(82,8) ,
10821	 => std_logic_vector(to_unsigned(79,8) ,
10822	 => std_logic_vector(to_unsigned(85,8) ,
10823	 => std_logic_vector(to_unsigned(85,8) ,
10824	 => std_logic_vector(to_unsigned(84,8) ,
10825	 => std_logic_vector(to_unsigned(74,8) ,
10826	 => std_logic_vector(to_unsigned(69,8) ,
10827	 => std_logic_vector(to_unsigned(69,8) ,
10828	 => std_logic_vector(to_unsigned(66,8) ,
10829	 => std_logic_vector(to_unsigned(69,8) ,
10830	 => std_logic_vector(to_unsigned(58,8) ,
10831	 => std_logic_vector(to_unsigned(64,8) ,
10832	 => std_logic_vector(to_unsigned(64,8) ,
10833	 => std_logic_vector(to_unsigned(65,8) ,
10834	 => std_logic_vector(to_unsigned(72,8) ,
10835	 => std_logic_vector(to_unsigned(70,8) ,
10836	 => std_logic_vector(to_unsigned(70,8) ,
10837	 => std_logic_vector(to_unsigned(73,8) ,
10838	 => std_logic_vector(to_unsigned(77,8) ,
10839	 => std_logic_vector(to_unsigned(87,8) ,
10840	 => std_logic_vector(to_unsigned(97,8) ,
10841	 => std_logic_vector(to_unsigned(92,8) ,
10842	 => std_logic_vector(to_unsigned(90,8) ,
10843	 => std_logic_vector(to_unsigned(92,8) ,
10844	 => std_logic_vector(to_unsigned(96,8) ,
10845	 => std_logic_vector(to_unsigned(96,8) ,
10846	 => std_logic_vector(to_unsigned(99,8) ,
10847	 => std_logic_vector(to_unsigned(104,8) ,
10848	 => std_logic_vector(to_unsigned(107,8) ,
10849	 => std_logic_vector(to_unsigned(104,8) ,
10850	 => std_logic_vector(to_unsigned(103,8) ,
10851	 => std_logic_vector(to_unsigned(111,8) ,
10852	 => std_logic_vector(to_unsigned(114,8) ,
10853	 => std_logic_vector(to_unsigned(111,8) ,
10854	 => std_logic_vector(to_unsigned(115,8) ,
10855	 => std_logic_vector(to_unsigned(118,8) ,
10856	 => std_logic_vector(to_unsigned(105,8) ,
10857	 => std_logic_vector(to_unsigned(105,8) ,
10858	 => std_logic_vector(to_unsigned(122,8) ,
10859	 => std_logic_vector(to_unsigned(122,8) ,
10860	 => std_logic_vector(to_unsigned(128,8) ,
10861	 => std_logic_vector(to_unsigned(134,8) ,
10862	 => std_logic_vector(to_unsigned(138,8) ,
10863	 => std_logic_vector(to_unsigned(144,8) ,
10864	 => std_logic_vector(to_unsigned(147,8) ,
10865	 => std_logic_vector(to_unsigned(144,8) ,
10866	 => std_logic_vector(to_unsigned(142,8) ,
10867	 => std_logic_vector(to_unsigned(147,8) ,
10868	 => std_logic_vector(to_unsigned(151,8) ,
10869	 => std_logic_vector(to_unsigned(151,8) ,
10870	 => std_logic_vector(to_unsigned(156,8) ,
10871	 => std_logic_vector(to_unsigned(152,8) ,
10872	 => std_logic_vector(to_unsigned(154,8) ,
10873	 => std_logic_vector(to_unsigned(157,8) ,
10874	 => std_logic_vector(to_unsigned(154,8) ,
10875	 => std_logic_vector(to_unsigned(152,8) ,
10876	 => std_logic_vector(to_unsigned(156,8) ,
10877	 => std_logic_vector(to_unsigned(161,8) ,
10878	 => std_logic_vector(to_unsigned(157,8) ,
10879	 => std_logic_vector(to_unsigned(156,8) ,
10880	 => std_logic_vector(to_unsigned(156,8) ,
10881	 => std_logic_vector(to_unsigned(125,8) ,
10882	 => std_logic_vector(to_unsigned(119,8) ,
10883	 => std_logic_vector(to_unsigned(114,8) ,
10884	 => std_logic_vector(to_unsigned(116,8) ,
10885	 => std_logic_vector(to_unsigned(119,8) ,
10886	 => std_logic_vector(to_unsigned(124,8) ,
10887	 => std_logic_vector(to_unsigned(125,8) ,
10888	 => std_logic_vector(to_unsigned(130,8) ,
10889	 => std_logic_vector(to_unsigned(131,8) ,
10890	 => std_logic_vector(to_unsigned(127,8) ,
10891	 => std_logic_vector(to_unsigned(125,8) ,
10892	 => std_logic_vector(to_unsigned(128,8) ,
10893	 => std_logic_vector(to_unsigned(131,8) ,
10894	 => std_logic_vector(to_unsigned(134,8) ,
10895	 => std_logic_vector(to_unsigned(138,8) ,
10896	 => std_logic_vector(to_unsigned(136,8) ,
10897	 => std_logic_vector(to_unsigned(128,8) ,
10898	 => std_logic_vector(to_unsigned(122,8) ,
10899	 => std_logic_vector(to_unsigned(125,8) ,
10900	 => std_logic_vector(to_unsigned(124,8) ,
10901	 => std_logic_vector(to_unsigned(121,8) ,
10902	 => std_logic_vector(to_unsigned(128,8) ,
10903	 => std_logic_vector(to_unsigned(130,8) ,
10904	 => std_logic_vector(to_unsigned(133,8) ,
10905	 => std_logic_vector(to_unsigned(133,8) ,
10906	 => std_logic_vector(to_unsigned(130,8) ,
10907	 => std_logic_vector(to_unsigned(116,8) ,
10908	 => std_logic_vector(to_unsigned(108,8) ,
10909	 => std_logic_vector(to_unsigned(108,8) ,
10910	 => std_logic_vector(to_unsigned(104,8) ,
10911	 => std_logic_vector(to_unsigned(107,8) ,
10912	 => std_logic_vector(to_unsigned(108,8) ,
10913	 => std_logic_vector(to_unsigned(115,8) ,
10914	 => std_logic_vector(to_unsigned(121,8) ,
10915	 => std_logic_vector(to_unsigned(116,8) ,
10916	 => std_logic_vector(to_unsigned(118,8) ,
10917	 => std_logic_vector(to_unsigned(124,8) ,
10918	 => std_logic_vector(to_unsigned(118,8) ,
10919	 => std_logic_vector(to_unsigned(119,8) ,
10920	 => std_logic_vector(to_unsigned(118,8) ,
10921	 => std_logic_vector(to_unsigned(115,8) ,
10922	 => std_logic_vector(to_unsigned(124,8) ,
10923	 => std_logic_vector(to_unsigned(131,8) ,
10924	 => std_logic_vector(to_unsigned(130,8) ,
10925	 => std_logic_vector(to_unsigned(125,8) ,
10926	 => std_logic_vector(to_unsigned(127,8) ,
10927	 => std_logic_vector(to_unsigned(131,8) ,
10928	 => std_logic_vector(to_unsigned(134,8) ,
10929	 => std_logic_vector(to_unsigned(130,8) ,
10930	 => std_logic_vector(to_unsigned(130,8) ,
10931	 => std_logic_vector(to_unsigned(127,8) ,
10932	 => std_logic_vector(to_unsigned(125,8) ,
10933	 => std_logic_vector(to_unsigned(131,8) ,
10934	 => std_logic_vector(to_unsigned(133,8) ,
10935	 => std_logic_vector(to_unsigned(128,8) ,
10936	 => std_logic_vector(to_unsigned(130,8) ,
10937	 => std_logic_vector(to_unsigned(130,8) ,
10938	 => std_logic_vector(to_unsigned(141,8) ,
10939	 => std_logic_vector(to_unsigned(144,8) ,
10940	 => std_logic_vector(to_unsigned(142,8) ,
10941	 => std_logic_vector(to_unsigned(142,8) ,
10942	 => std_logic_vector(to_unsigned(134,8) ,
10943	 => std_logic_vector(to_unsigned(141,8) ,
10944	 => std_logic_vector(to_unsigned(151,8) ,
10945	 => std_logic_vector(to_unsigned(149,8) ,
10946	 => std_logic_vector(to_unsigned(144,8) ,
10947	 => std_logic_vector(to_unsigned(138,8) ,
10948	 => std_logic_vector(to_unsigned(139,8) ,
10949	 => std_logic_vector(to_unsigned(142,8) ,
10950	 => std_logic_vector(to_unsigned(139,8) ,
10951	 => std_logic_vector(to_unsigned(139,8) ,
10952	 => std_logic_vector(to_unsigned(138,8) ,
10953	 => std_logic_vector(to_unsigned(141,8) ,
10954	 => std_logic_vector(to_unsigned(130,8) ,
10955	 => std_logic_vector(to_unsigned(115,8) ,
10956	 => std_logic_vector(to_unsigned(130,8) ,
10957	 => std_logic_vector(to_unsigned(138,8) ,
10958	 => std_logic_vector(to_unsigned(134,8) ,
10959	 => std_logic_vector(to_unsigned(133,8) ,
10960	 => std_logic_vector(to_unsigned(134,8) ,
10961	 => std_logic_vector(to_unsigned(133,8) ,
10962	 => std_logic_vector(to_unsigned(131,8) ,
10963	 => std_logic_vector(to_unsigned(134,8) ,
10964	 => std_logic_vector(to_unsigned(133,8) ,
10965	 => std_logic_vector(to_unsigned(134,8) ,
10966	 => std_logic_vector(to_unsigned(139,8) ,
10967	 => std_logic_vector(to_unsigned(141,8) ,
10968	 => std_logic_vector(to_unsigned(136,8) ,
10969	 => std_logic_vector(to_unsigned(125,8) ,
10970	 => std_logic_vector(to_unsigned(138,8) ,
10971	 => std_logic_vector(to_unsigned(149,8) ,
10972	 => std_logic_vector(to_unsigned(136,8) ,
10973	 => std_logic_vector(to_unsigned(112,8) ,
10974	 => std_logic_vector(to_unsigned(97,8) ,
10975	 => std_logic_vector(to_unsigned(99,8) ,
10976	 => std_logic_vector(to_unsigned(100,8) ,
10977	 => std_logic_vector(to_unsigned(114,8) ,
10978	 => std_logic_vector(to_unsigned(131,8) ,
10979	 => std_logic_vector(to_unsigned(121,8) ,
10980	 => std_logic_vector(to_unsigned(101,8) ,
10981	 => std_logic_vector(to_unsigned(95,8) ,
10982	 => std_logic_vector(to_unsigned(99,8) ,
10983	 => std_logic_vector(to_unsigned(107,8) ,
10984	 => std_logic_vector(to_unsigned(116,8) ,
10985	 => std_logic_vector(to_unsigned(100,8) ,
10986	 => std_logic_vector(to_unsigned(88,8) ,
10987	 => std_logic_vector(to_unsigned(73,8) ,
10988	 => std_logic_vector(to_unsigned(77,8) ,
10989	 => std_logic_vector(to_unsigned(79,8) ,
10990	 => std_logic_vector(to_unsigned(72,8) ,
10991	 => std_logic_vector(to_unsigned(73,8) ,
10992	 => std_logic_vector(to_unsigned(73,8) ,
10993	 => std_logic_vector(to_unsigned(85,8) ,
10994	 => std_logic_vector(to_unsigned(80,8) ,
10995	 => std_logic_vector(to_unsigned(80,8) ,
10996	 => std_logic_vector(to_unsigned(85,8) ,
10997	 => std_logic_vector(to_unsigned(87,8) ,
10998	 => std_logic_vector(to_unsigned(90,8) ,
10999	 => std_logic_vector(to_unsigned(87,8) ,
11000	 => std_logic_vector(to_unsigned(93,8) ,
11001	 => std_logic_vector(to_unsigned(99,8) ,
11002	 => std_logic_vector(to_unsigned(88,8) ,
11003	 => std_logic_vector(to_unsigned(99,8) ,
11004	 => std_logic_vector(to_unsigned(130,8) ,
11005	 => std_logic_vector(to_unsigned(131,8) ,
11006	 => std_logic_vector(to_unsigned(107,8) ,
11007	 => std_logic_vector(to_unsigned(115,8) ,
11008	 => std_logic_vector(to_unsigned(119,8) ,
11009	 => std_logic_vector(to_unsigned(116,8) ,
11010	 => std_logic_vector(to_unsigned(115,8) ,
11011	 => std_logic_vector(to_unsigned(112,8) ,
11012	 => std_logic_vector(to_unsigned(105,8) ,
11013	 => std_logic_vector(to_unsigned(105,8) ,
11014	 => std_logic_vector(to_unsigned(100,8) ,
11015	 => std_logic_vector(to_unsigned(92,8) ,
11016	 => std_logic_vector(to_unsigned(85,8) ,
11017	 => std_logic_vector(to_unsigned(92,8) ,
11018	 => std_logic_vector(to_unsigned(96,8) ,
11019	 => std_logic_vector(to_unsigned(93,8) ,
11020	 => std_logic_vector(to_unsigned(92,8) ,
11021	 => std_logic_vector(to_unsigned(95,8) ,
11022	 => std_logic_vector(to_unsigned(99,8) ,
11023	 => std_logic_vector(to_unsigned(93,8) ,
11024	 => std_logic_vector(to_unsigned(104,8) ,
11025	 => std_logic_vector(to_unsigned(104,8) ,
11026	 => std_logic_vector(to_unsigned(100,8) ,
11027	 => std_logic_vector(to_unsigned(107,8) ,
11028	 => std_logic_vector(to_unsigned(104,8) ,
11029	 => std_logic_vector(to_unsigned(93,8) ,
11030	 => std_logic_vector(to_unsigned(87,8) ,
11031	 => std_logic_vector(to_unsigned(86,8) ,
11032	 => std_logic_vector(to_unsigned(86,8) ,
11033	 => std_logic_vector(to_unsigned(88,8) ,
11034	 => std_logic_vector(to_unsigned(85,8) ,
11035	 => std_logic_vector(to_unsigned(85,8) ,
11036	 => std_logic_vector(to_unsigned(81,8) ,
11037	 => std_logic_vector(to_unsigned(85,8) ,
11038	 => std_logic_vector(to_unsigned(86,8) ,
11039	 => std_logic_vector(to_unsigned(79,8) ,
11040	 => std_logic_vector(to_unsigned(77,8) ,
11041	 => std_logic_vector(to_unsigned(97,8) ,
11042	 => std_logic_vector(to_unsigned(88,8) ,
11043	 => std_logic_vector(to_unsigned(78,8) ,
11044	 => std_logic_vector(to_unsigned(58,8) ,
11045	 => std_logic_vector(to_unsigned(54,8) ,
11046	 => std_logic_vector(to_unsigned(73,8) ,
11047	 => std_logic_vector(to_unsigned(81,8) ,
11048	 => std_logic_vector(to_unsigned(78,8) ,
11049	 => std_logic_vector(to_unsigned(84,8) ,
11050	 => std_logic_vector(to_unsigned(80,8) ,
11051	 => std_logic_vector(to_unsigned(85,8) ,
11052	 => std_logic_vector(to_unsigned(88,8) ,
11053	 => std_logic_vector(to_unsigned(92,8) ,
11054	 => std_logic_vector(to_unsigned(91,8) ,
11055	 => std_logic_vector(to_unsigned(82,8) ,
11056	 => std_logic_vector(to_unsigned(77,8) ,
11057	 => std_logic_vector(to_unsigned(79,8) ,
11058	 => std_logic_vector(to_unsigned(85,8) ,
11059	 => std_logic_vector(to_unsigned(88,8) ,
11060	 => std_logic_vector(to_unsigned(70,8) ,
11061	 => std_logic_vector(to_unsigned(70,8) ,
11062	 => std_logic_vector(to_unsigned(81,8) ,
11063	 => std_logic_vector(to_unsigned(86,8) ,
11064	 => std_logic_vector(to_unsigned(95,8) ,
11065	 => std_logic_vector(to_unsigned(97,8) ,
11066	 => std_logic_vector(to_unsigned(99,8) ,
11067	 => std_logic_vector(to_unsigned(90,8) ,
11068	 => std_logic_vector(to_unsigned(103,8) ,
11069	 => std_logic_vector(to_unsigned(103,8) ,
11070	 => std_logic_vector(to_unsigned(81,8) ,
11071	 => std_logic_vector(to_unsigned(81,8) ,
11072	 => std_logic_vector(to_unsigned(131,8) ,
11073	 => std_logic_vector(to_unsigned(95,8) ,
11074	 => std_logic_vector(to_unsigned(70,8) ,
11075	 => std_logic_vector(to_unsigned(96,8) ,
11076	 => std_logic_vector(to_unsigned(88,8) ,
11077	 => std_logic_vector(to_unsigned(78,8) ,
11078	 => std_logic_vector(to_unsigned(85,8) ,
11079	 => std_logic_vector(to_unsigned(93,8) ,
11080	 => std_logic_vector(to_unsigned(103,8) ,
11081	 => std_logic_vector(to_unsigned(100,8) ,
11082	 => std_logic_vector(to_unsigned(96,8) ,
11083	 => std_logic_vector(to_unsigned(93,8) ,
11084	 => std_logic_vector(to_unsigned(78,8) ,
11085	 => std_logic_vector(to_unsigned(81,8) ,
11086	 => std_logic_vector(to_unsigned(81,8) ,
11087	 => std_logic_vector(to_unsigned(80,8) ,
11088	 => std_logic_vector(to_unsigned(74,8) ,
11089	 => std_logic_vector(to_unsigned(82,8) ,
11090	 => std_logic_vector(to_unsigned(92,8) ,
11091	 => std_logic_vector(to_unsigned(86,8) ,
11092	 => std_logic_vector(to_unsigned(78,8) ,
11093	 => std_logic_vector(to_unsigned(76,8) ,
11094	 => std_logic_vector(to_unsigned(76,8) ,
11095	 => std_logic_vector(to_unsigned(76,8) ,
11096	 => std_logic_vector(to_unsigned(84,8) ,
11097	 => std_logic_vector(to_unsigned(85,8) ,
11098	 => std_logic_vector(to_unsigned(80,8) ,
11099	 => std_logic_vector(to_unsigned(90,8) ,
11100	 => std_logic_vector(to_unsigned(85,8) ,
11101	 => std_logic_vector(to_unsigned(81,8) ,
11102	 => std_logic_vector(to_unsigned(90,8) ,
11103	 => std_logic_vector(to_unsigned(80,8) ,
11104	 => std_logic_vector(to_unsigned(84,8) ,
11105	 => std_logic_vector(to_unsigned(81,8) ,
11106	 => std_logic_vector(to_unsigned(79,8) ,
11107	 => std_logic_vector(to_unsigned(84,8) ,
11108	 => std_logic_vector(to_unsigned(70,8) ,
11109	 => std_logic_vector(to_unsigned(80,8) ,
11110	 => std_logic_vector(to_unsigned(85,8) ,
11111	 => std_logic_vector(to_unsigned(77,8) ,
11112	 => std_logic_vector(to_unsigned(77,8) ,
11113	 => std_logic_vector(to_unsigned(79,8) ,
11114	 => std_logic_vector(to_unsigned(84,8) ,
11115	 => std_logic_vector(to_unsigned(86,8) ,
11116	 => std_logic_vector(to_unsigned(76,8) ,
11117	 => std_logic_vector(to_unsigned(60,8) ,
11118	 => std_logic_vector(to_unsigned(59,8) ,
11119	 => std_logic_vector(to_unsigned(62,8) ,
11120	 => std_logic_vector(to_unsigned(54,8) ,
11121	 => std_logic_vector(to_unsigned(60,8) ,
11122	 => std_logic_vector(to_unsigned(57,8) ,
11123	 => std_logic_vector(to_unsigned(6,8) ,
11124	 => std_logic_vector(to_unsigned(0,8) ,
11125	 => std_logic_vector(to_unsigned(0,8) ,
11126	 => std_logic_vector(to_unsigned(8,8) ,
11127	 => std_logic_vector(to_unsigned(51,8) ,
11128	 => std_logic_vector(to_unsigned(52,8) ,
11129	 => std_logic_vector(to_unsigned(56,8) ,
11130	 => std_logic_vector(to_unsigned(87,8) ,
11131	 => std_logic_vector(to_unsigned(107,8) ,
11132	 => std_logic_vector(to_unsigned(103,8) ,
11133	 => std_logic_vector(to_unsigned(90,8) ,
11134	 => std_logic_vector(to_unsigned(84,8) ,
11135	 => std_logic_vector(to_unsigned(95,8) ,
11136	 => std_logic_vector(to_unsigned(92,8) ,
11137	 => std_logic_vector(to_unsigned(88,8) ,
11138	 => std_logic_vector(to_unsigned(76,8) ,
11139	 => std_logic_vector(to_unsigned(78,8) ,
11140	 => std_logic_vector(to_unsigned(86,8) ,
11141	 => std_logic_vector(to_unsigned(72,8) ,
11142	 => std_logic_vector(to_unsigned(62,8) ,
11143	 => std_logic_vector(to_unsigned(66,8) ,
11144	 => std_logic_vector(to_unsigned(56,8) ,
11145	 => std_logic_vector(to_unsigned(54,8) ,
11146	 => std_logic_vector(to_unsigned(57,8) ,
11147	 => std_logic_vector(to_unsigned(54,8) ,
11148	 => std_logic_vector(to_unsigned(58,8) ,
11149	 => std_logic_vector(to_unsigned(69,8) ,
11150	 => std_logic_vector(to_unsigned(70,8) ,
11151	 => std_logic_vector(to_unsigned(77,8) ,
11152	 => std_logic_vector(to_unsigned(72,8) ,
11153	 => std_logic_vector(to_unsigned(67,8) ,
11154	 => std_logic_vector(to_unsigned(70,8) ,
11155	 => std_logic_vector(to_unsigned(77,8) ,
11156	 => std_logic_vector(to_unsigned(70,8) ,
11157	 => std_logic_vector(to_unsigned(73,8) ,
11158	 => std_logic_vector(to_unsigned(78,8) ,
11159	 => std_logic_vector(to_unsigned(93,8) ,
11160	 => std_logic_vector(to_unsigned(100,8) ,
11161	 => std_logic_vector(to_unsigned(105,8) ,
11162	 => std_logic_vector(to_unsigned(108,8) ,
11163	 => std_logic_vector(to_unsigned(112,8) ,
11164	 => std_logic_vector(to_unsigned(107,8) ,
11165	 => std_logic_vector(to_unsigned(109,8) ,
11166	 => std_logic_vector(to_unsigned(127,8) ,
11167	 => std_logic_vector(to_unsigned(122,8) ,
11168	 => std_logic_vector(to_unsigned(124,8) ,
11169	 => std_logic_vector(to_unsigned(133,8) ,
11170	 => std_logic_vector(to_unsigned(127,8) ,
11171	 => std_logic_vector(to_unsigned(130,8) ,
11172	 => std_logic_vector(to_unsigned(133,8) ,
11173	 => std_logic_vector(to_unsigned(127,8) ,
11174	 => std_logic_vector(to_unsigned(136,8) ,
11175	 => std_logic_vector(to_unsigned(141,8) ,
11176	 => std_logic_vector(to_unsigned(138,8) ,
11177	 => std_logic_vector(to_unsigned(138,8) ,
11178	 => std_logic_vector(to_unsigned(147,8) ,
11179	 => std_logic_vector(to_unsigned(142,8) ,
11180	 => std_logic_vector(to_unsigned(149,8) ,
11181	 => std_logic_vector(to_unsigned(156,8) ,
11182	 => std_logic_vector(to_unsigned(151,8) ,
11183	 => std_logic_vector(to_unsigned(156,8) ,
11184	 => std_logic_vector(to_unsigned(159,8) ,
11185	 => std_logic_vector(to_unsigned(156,8) ,
11186	 => std_logic_vector(to_unsigned(157,8) ,
11187	 => std_logic_vector(to_unsigned(161,8) ,
11188	 => std_logic_vector(to_unsigned(159,8) ,
11189	 => std_logic_vector(to_unsigned(157,8) ,
11190	 => std_logic_vector(to_unsigned(159,8) ,
11191	 => std_logic_vector(to_unsigned(157,8) ,
11192	 => std_logic_vector(to_unsigned(156,8) ,
11193	 => std_logic_vector(to_unsigned(163,8) ,
11194	 => std_logic_vector(to_unsigned(161,8) ,
11195	 => std_logic_vector(to_unsigned(157,8) ,
11196	 => std_logic_vector(to_unsigned(157,8) ,
11197	 => std_logic_vector(to_unsigned(163,8) ,
11198	 => std_logic_vector(to_unsigned(163,8) ,
11199	 => std_logic_vector(to_unsigned(163,8) ,
11200	 => std_logic_vector(to_unsigned(164,8) ,
11201	 => std_logic_vector(to_unsigned(118,8) ,
11202	 => std_logic_vector(to_unsigned(115,8) ,
11203	 => std_logic_vector(to_unsigned(122,8) ,
11204	 => std_logic_vector(to_unsigned(130,8) ,
11205	 => std_logic_vector(to_unsigned(124,8) ,
11206	 => std_logic_vector(to_unsigned(130,8) ,
11207	 => std_logic_vector(to_unsigned(131,8) ,
11208	 => std_logic_vector(to_unsigned(130,8) ,
11209	 => std_logic_vector(to_unsigned(130,8) ,
11210	 => std_logic_vector(to_unsigned(119,8) ,
11211	 => std_logic_vector(to_unsigned(116,8) ,
11212	 => std_logic_vector(to_unsigned(127,8) ,
11213	 => std_logic_vector(to_unsigned(130,8) ,
11214	 => std_logic_vector(to_unsigned(136,8) ,
11215	 => std_logic_vector(to_unsigned(142,8) ,
11216	 => std_logic_vector(to_unsigned(138,8) ,
11217	 => std_logic_vector(to_unsigned(130,8) ,
11218	 => std_logic_vector(to_unsigned(130,8) ,
11219	 => std_logic_vector(to_unsigned(127,8) ,
11220	 => std_logic_vector(to_unsigned(130,8) ,
11221	 => std_logic_vector(to_unsigned(125,8) ,
11222	 => std_logic_vector(to_unsigned(136,8) ,
11223	 => std_logic_vector(to_unsigned(139,8) ,
11224	 => std_logic_vector(to_unsigned(138,8) ,
11225	 => std_logic_vector(to_unsigned(138,8) ,
11226	 => std_logic_vector(to_unsigned(139,8) ,
11227	 => std_logic_vector(to_unsigned(130,8) ,
11228	 => std_logic_vector(to_unsigned(118,8) ,
11229	 => std_logic_vector(to_unsigned(116,8) ,
11230	 => std_logic_vector(to_unsigned(112,8) ,
11231	 => std_logic_vector(to_unsigned(107,8) ,
11232	 => std_logic_vector(to_unsigned(111,8) ,
11233	 => std_logic_vector(to_unsigned(116,8) ,
11234	 => std_logic_vector(to_unsigned(122,8) ,
11235	 => std_logic_vector(to_unsigned(122,8) ,
11236	 => std_logic_vector(to_unsigned(124,8) ,
11237	 => std_logic_vector(to_unsigned(124,8) ,
11238	 => std_logic_vector(to_unsigned(121,8) ,
11239	 => std_logic_vector(to_unsigned(124,8) ,
11240	 => std_logic_vector(to_unsigned(121,8) ,
11241	 => std_logic_vector(to_unsigned(119,8) ,
11242	 => std_logic_vector(to_unsigned(124,8) ,
11243	 => std_logic_vector(to_unsigned(127,8) ,
11244	 => std_logic_vector(to_unsigned(128,8) ,
11245	 => std_logic_vector(to_unsigned(131,8) ,
11246	 => std_logic_vector(to_unsigned(127,8) ,
11247	 => std_logic_vector(to_unsigned(130,8) ,
11248	 => std_logic_vector(to_unsigned(138,8) ,
11249	 => std_logic_vector(to_unsigned(136,8) ,
11250	 => std_logic_vector(to_unsigned(138,8) ,
11251	 => std_logic_vector(to_unsigned(133,8) ,
11252	 => std_logic_vector(to_unsigned(130,8) ,
11253	 => std_logic_vector(to_unsigned(138,8) ,
11254	 => std_logic_vector(to_unsigned(138,8) ,
11255	 => std_logic_vector(to_unsigned(133,8) ,
11256	 => std_logic_vector(to_unsigned(136,8) ,
11257	 => std_logic_vector(to_unsigned(133,8) ,
11258	 => std_logic_vector(to_unsigned(142,8) ,
11259	 => std_logic_vector(to_unsigned(149,8) ,
11260	 => std_logic_vector(to_unsigned(152,8) ,
11261	 => std_logic_vector(to_unsigned(147,8) ,
11262	 => std_logic_vector(to_unsigned(144,8) ,
11263	 => std_logic_vector(to_unsigned(149,8) ,
11264	 => std_logic_vector(to_unsigned(146,8) ,
11265	 => std_logic_vector(to_unsigned(136,8) ,
11266	 => std_logic_vector(to_unsigned(146,8) ,
11267	 => std_logic_vector(to_unsigned(138,8) ,
11268	 => std_logic_vector(to_unsigned(134,8) ,
11269	 => std_logic_vector(to_unsigned(142,8) ,
11270	 => std_logic_vector(to_unsigned(139,8) ,
11271	 => std_logic_vector(to_unsigned(134,8) ,
11272	 => std_logic_vector(to_unsigned(139,8) ,
11273	 => std_logic_vector(to_unsigned(146,8) ,
11274	 => std_logic_vector(to_unsigned(128,8) ,
11275	 => std_logic_vector(to_unsigned(108,8) ,
11276	 => std_logic_vector(to_unsigned(124,8) ,
11277	 => std_logic_vector(to_unsigned(138,8) ,
11278	 => std_logic_vector(to_unsigned(134,8) ,
11279	 => std_logic_vector(to_unsigned(130,8) ,
11280	 => std_logic_vector(to_unsigned(134,8) ,
11281	 => std_logic_vector(to_unsigned(138,8) ,
11282	 => std_logic_vector(to_unsigned(133,8) ,
11283	 => std_logic_vector(to_unsigned(133,8) ,
11284	 => std_logic_vector(to_unsigned(133,8) ,
11285	 => std_logic_vector(to_unsigned(144,8) ,
11286	 => std_logic_vector(to_unsigned(142,8) ,
11287	 => std_logic_vector(to_unsigned(144,8) ,
11288	 => std_logic_vector(to_unsigned(141,8) ,
11289	 => std_logic_vector(to_unsigned(130,8) ,
11290	 => std_logic_vector(to_unsigned(142,8) ,
11291	 => std_logic_vector(to_unsigned(139,8) ,
11292	 => std_logic_vector(to_unsigned(125,8) ,
11293	 => std_logic_vector(to_unsigned(115,8) ,
11294	 => std_logic_vector(to_unsigned(104,8) ,
11295	 => std_logic_vector(to_unsigned(107,8) ,
11296	 => std_logic_vector(to_unsigned(109,8) ,
11297	 => std_logic_vector(to_unsigned(104,8) ,
11298	 => std_logic_vector(to_unsigned(124,8) ,
11299	 => std_logic_vector(to_unsigned(118,8) ,
11300	 => std_logic_vector(to_unsigned(104,8) ,
11301	 => std_logic_vector(to_unsigned(115,8) ,
11302	 => std_logic_vector(to_unsigned(112,8) ,
11303	 => std_logic_vector(to_unsigned(115,8) ,
11304	 => std_logic_vector(to_unsigned(118,8) ,
11305	 => std_logic_vector(to_unsigned(107,8) ,
11306	 => std_logic_vector(to_unsigned(93,8) ,
11307	 => std_logic_vector(to_unsigned(78,8) ,
11308	 => std_logic_vector(to_unsigned(80,8) ,
11309	 => std_logic_vector(to_unsigned(80,8) ,
11310	 => std_logic_vector(to_unsigned(84,8) ,
11311	 => std_logic_vector(to_unsigned(81,8) ,
11312	 => std_logic_vector(to_unsigned(85,8) ,
11313	 => std_logic_vector(to_unsigned(86,8) ,
11314	 => std_logic_vector(to_unsigned(80,8) ,
11315	 => std_logic_vector(to_unsigned(82,8) ,
11316	 => std_logic_vector(to_unsigned(90,8) ,
11317	 => std_logic_vector(to_unsigned(93,8) ,
11318	 => std_logic_vector(to_unsigned(96,8) ,
11319	 => std_logic_vector(to_unsigned(93,8) ,
11320	 => std_logic_vector(to_unsigned(101,8) ,
11321	 => std_logic_vector(to_unsigned(108,8) ,
11322	 => std_logic_vector(to_unsigned(96,8) ,
11323	 => std_logic_vector(to_unsigned(103,8) ,
11324	 => std_logic_vector(to_unsigned(131,8) ,
11325	 => std_logic_vector(to_unsigned(134,8) ,
11326	 => std_logic_vector(to_unsigned(109,8) ,
11327	 => std_logic_vector(to_unsigned(114,8) ,
11328	 => std_logic_vector(to_unsigned(128,8) ,
11329	 => std_logic_vector(to_unsigned(124,8) ,
11330	 => std_logic_vector(to_unsigned(121,8) ,
11331	 => std_logic_vector(to_unsigned(121,8) ,
11332	 => std_logic_vector(to_unsigned(116,8) ,
11333	 => std_logic_vector(to_unsigned(112,8) ,
11334	 => std_logic_vector(to_unsigned(107,8) ,
11335	 => std_logic_vector(to_unsigned(100,8) ,
11336	 => std_logic_vector(to_unsigned(92,8) ,
11337	 => std_logic_vector(to_unsigned(91,8) ,
11338	 => std_logic_vector(to_unsigned(92,8) ,
11339	 => std_logic_vector(to_unsigned(101,8) ,
11340	 => std_logic_vector(to_unsigned(100,8) ,
11341	 => std_logic_vector(to_unsigned(103,8) ,
11342	 => std_logic_vector(to_unsigned(97,8) ,
11343	 => std_logic_vector(to_unsigned(104,8) ,
11344	 => std_logic_vector(to_unsigned(111,8) ,
11345	 => std_logic_vector(to_unsigned(108,8) ,
11346	 => std_logic_vector(to_unsigned(101,8) ,
11347	 => std_logic_vector(to_unsigned(109,8) ,
11348	 => std_logic_vector(to_unsigned(97,8) ,
11349	 => std_logic_vector(to_unsigned(82,8) ,
11350	 => std_logic_vector(to_unsigned(92,8) ,
11351	 => std_logic_vector(to_unsigned(91,8) ,
11352	 => std_logic_vector(to_unsigned(78,8) ,
11353	 => std_logic_vector(to_unsigned(85,8) ,
11354	 => std_logic_vector(to_unsigned(81,8) ,
11355	 => std_logic_vector(to_unsigned(90,8) ,
11356	 => std_logic_vector(to_unsigned(92,8) ,
11357	 => std_logic_vector(to_unsigned(91,8) ,
11358	 => std_logic_vector(to_unsigned(82,8) ,
11359	 => std_logic_vector(to_unsigned(78,8) ,
11360	 => std_logic_vector(to_unsigned(84,8) ,
11361	 => std_logic_vector(to_unsigned(107,8) ,
11362	 => std_logic_vector(to_unsigned(96,8) ,
11363	 => std_logic_vector(to_unsigned(81,8) ,
11364	 => std_logic_vector(to_unsigned(68,8) ,
11365	 => std_logic_vector(to_unsigned(74,8) ,
11366	 => std_logic_vector(to_unsigned(91,8) ,
11367	 => std_logic_vector(to_unsigned(88,8) ,
11368	 => std_logic_vector(to_unsigned(82,8) ,
11369	 => std_logic_vector(to_unsigned(87,8) ,
11370	 => std_logic_vector(to_unsigned(87,8) ,
11371	 => std_logic_vector(to_unsigned(88,8) ,
11372	 => std_logic_vector(to_unsigned(93,8) ,
11373	 => std_logic_vector(to_unsigned(92,8) ,
11374	 => std_logic_vector(to_unsigned(80,8) ,
11375	 => std_logic_vector(to_unsigned(79,8) ,
11376	 => std_logic_vector(to_unsigned(86,8) ,
11377	 => std_logic_vector(to_unsigned(81,8) ,
11378	 => std_logic_vector(to_unsigned(79,8) ,
11379	 => std_logic_vector(to_unsigned(88,8) ,
11380	 => std_logic_vector(to_unsigned(67,8) ,
11381	 => std_logic_vector(to_unsigned(62,8) ,
11382	 => std_logic_vector(to_unsigned(81,8) ,
11383	 => std_logic_vector(to_unsigned(91,8) ,
11384	 => std_logic_vector(to_unsigned(95,8) ,
11385	 => std_logic_vector(to_unsigned(101,8) ,
11386	 => std_logic_vector(to_unsigned(100,8) ,
11387	 => std_logic_vector(to_unsigned(87,8) ,
11388	 => std_logic_vector(to_unsigned(91,8) ,
11389	 => std_logic_vector(to_unsigned(95,8) ,
11390	 => std_logic_vector(to_unsigned(86,8) ,
11391	 => std_logic_vector(to_unsigned(92,8) ,
11392	 => std_logic_vector(to_unsigned(139,8) ,
11393	 => std_logic_vector(to_unsigned(114,8) ,
11394	 => std_logic_vector(to_unsigned(81,8) ,
11395	 => std_logic_vector(to_unsigned(91,8) ,
11396	 => std_logic_vector(to_unsigned(91,8) ,
11397	 => std_logic_vector(to_unsigned(90,8) ,
11398	 => std_logic_vector(to_unsigned(93,8) ,
11399	 => std_logic_vector(to_unsigned(99,8) ,
11400	 => std_logic_vector(to_unsigned(100,8) ,
11401	 => std_logic_vector(to_unsigned(100,8) ,
11402	 => std_logic_vector(to_unsigned(105,8) ,
11403	 => std_logic_vector(to_unsigned(96,8) ,
11404	 => std_logic_vector(to_unsigned(74,8) ,
11405	 => std_logic_vector(to_unsigned(86,8) ,
11406	 => std_logic_vector(to_unsigned(93,8) ,
11407	 => std_logic_vector(to_unsigned(84,8) ,
11408	 => std_logic_vector(to_unsigned(82,8) ,
11409	 => std_logic_vector(to_unsigned(92,8) ,
11410	 => std_logic_vector(to_unsigned(88,8) ,
11411	 => std_logic_vector(to_unsigned(90,8) ,
11412	 => std_logic_vector(to_unsigned(86,8) ,
11413	 => std_logic_vector(to_unsigned(81,8) ,
11414	 => std_logic_vector(to_unsigned(82,8) ,
11415	 => std_logic_vector(to_unsigned(87,8) ,
11416	 => std_logic_vector(to_unsigned(91,8) ,
11417	 => std_logic_vector(to_unsigned(86,8) ,
11418	 => std_logic_vector(to_unsigned(88,8) ,
11419	 => std_logic_vector(to_unsigned(90,8) ,
11420	 => std_logic_vector(to_unsigned(86,8) ,
11421	 => std_logic_vector(to_unsigned(87,8) ,
11422	 => std_logic_vector(to_unsigned(74,8) ,
11423	 => std_logic_vector(to_unsigned(71,8) ,
11424	 => std_logic_vector(to_unsigned(69,8) ,
11425	 => std_logic_vector(to_unsigned(74,8) ,
11426	 => std_logic_vector(to_unsigned(72,8) ,
11427	 => std_logic_vector(to_unsigned(68,8) ,
11428	 => std_logic_vector(to_unsigned(63,8) ,
11429	 => std_logic_vector(to_unsigned(67,8) ,
11430	 => std_logic_vector(to_unsigned(77,8) ,
11431	 => std_logic_vector(to_unsigned(65,8) ,
11432	 => std_logic_vector(to_unsigned(68,8) ,
11433	 => std_logic_vector(to_unsigned(87,8) ,
11434	 => std_logic_vector(to_unsigned(91,8) ,
11435	 => std_logic_vector(to_unsigned(81,8) ,
11436	 => std_logic_vector(to_unsigned(82,8) ,
11437	 => std_logic_vector(to_unsigned(70,8) ,
11438	 => std_logic_vector(to_unsigned(74,8) ,
11439	 => std_logic_vector(to_unsigned(60,8) ,
11440	 => std_logic_vector(to_unsigned(46,8) ,
11441	 => std_logic_vector(to_unsigned(50,8) ,
11442	 => std_logic_vector(to_unsigned(57,8) ,
11443	 => std_logic_vector(to_unsigned(17,8) ,
11444	 => std_logic_vector(to_unsigned(0,8) ,
11445	 => std_logic_vector(to_unsigned(0,8) ,
11446	 => std_logic_vector(to_unsigned(2,8) ,
11447	 => std_logic_vector(to_unsigned(37,8) ,
11448	 => std_logic_vector(to_unsigned(53,8) ,
11449	 => std_logic_vector(to_unsigned(51,8) ,
11450	 => std_logic_vector(to_unsigned(82,8) ,
11451	 => std_logic_vector(to_unsigned(104,8) ,
11452	 => std_logic_vector(to_unsigned(92,8) ,
11453	 => std_logic_vector(to_unsigned(77,8) ,
11454	 => std_logic_vector(to_unsigned(73,8) ,
11455	 => std_logic_vector(to_unsigned(95,8) ,
11456	 => std_logic_vector(to_unsigned(84,8) ,
11457	 => std_logic_vector(to_unsigned(68,8) ,
11458	 => std_logic_vector(to_unsigned(54,8) ,
11459	 => std_logic_vector(to_unsigned(55,8) ,
11460	 => std_logic_vector(to_unsigned(71,8) ,
11461	 => std_logic_vector(to_unsigned(52,8) ,
11462	 => std_logic_vector(to_unsigned(44,8) ,
11463	 => std_logic_vector(to_unsigned(51,8) ,
11464	 => std_logic_vector(to_unsigned(48,8) ,
11465	 => std_logic_vector(to_unsigned(55,8) ,
11466	 => std_logic_vector(to_unsigned(61,8) ,
11467	 => std_logic_vector(to_unsigned(57,8) ,
11468	 => std_logic_vector(to_unsigned(67,8) ,
11469	 => std_logic_vector(to_unsigned(76,8) ,
11470	 => std_logic_vector(to_unsigned(79,8) ,
11471	 => std_logic_vector(to_unsigned(72,8) ,
11472	 => std_logic_vector(to_unsigned(63,8) ,
11473	 => std_logic_vector(to_unsigned(58,8) ,
11474	 => std_logic_vector(to_unsigned(61,8) ,
11475	 => std_logic_vector(to_unsigned(68,8) ,
11476	 => std_logic_vector(to_unsigned(69,8) ,
11477	 => std_logic_vector(to_unsigned(65,8) ,
11478	 => std_logic_vector(to_unsigned(67,8) ,
11479	 => std_logic_vector(to_unsigned(76,8) ,
11480	 => std_logic_vector(to_unsigned(80,8) ,
11481	 => std_logic_vector(to_unsigned(91,8) ,
11482	 => std_logic_vector(to_unsigned(100,8) ,
11483	 => std_logic_vector(to_unsigned(114,8) ,
11484	 => std_logic_vector(to_unsigned(122,8) ,
11485	 => std_logic_vector(to_unsigned(109,8) ,
11486	 => std_logic_vector(to_unsigned(105,8) ,
11487	 => std_logic_vector(to_unsigned(97,8) ,
11488	 => std_logic_vector(to_unsigned(104,8) ,
11489	 => std_logic_vector(to_unsigned(127,8) ,
11490	 => std_logic_vector(to_unsigned(134,8) ,
11491	 => std_logic_vector(to_unsigned(144,8) ,
11492	 => std_logic_vector(to_unsigned(149,8) ,
11493	 => std_logic_vector(to_unsigned(147,8) ,
11494	 => std_logic_vector(to_unsigned(141,8) ,
11495	 => std_logic_vector(to_unsigned(142,8) ,
11496	 => std_logic_vector(to_unsigned(152,8) ,
11497	 => std_logic_vector(to_unsigned(146,8) ,
11498	 => std_logic_vector(to_unsigned(154,8) ,
11499	 => std_logic_vector(to_unsigned(157,8) ,
11500	 => std_logic_vector(to_unsigned(156,8) ,
11501	 => std_logic_vector(to_unsigned(159,8) ,
11502	 => std_logic_vector(to_unsigned(161,8) ,
11503	 => std_logic_vector(to_unsigned(161,8) ,
11504	 => std_logic_vector(to_unsigned(161,8) ,
11505	 => std_logic_vector(to_unsigned(157,8) ,
11506	 => std_logic_vector(to_unsigned(159,8) ,
11507	 => std_logic_vector(to_unsigned(164,8) ,
11508	 => std_logic_vector(to_unsigned(163,8) ,
11509	 => std_logic_vector(to_unsigned(159,8) ,
11510	 => std_logic_vector(to_unsigned(163,8) ,
11511	 => std_logic_vector(to_unsigned(163,8) ,
11512	 => std_logic_vector(to_unsigned(163,8) ,
11513	 => std_logic_vector(to_unsigned(168,8) ,
11514	 => std_logic_vector(to_unsigned(168,8) ,
11515	 => std_logic_vector(to_unsigned(163,8) ,
11516	 => std_logic_vector(to_unsigned(161,8) ,
11517	 => std_logic_vector(to_unsigned(166,8) ,
11518	 => std_logic_vector(to_unsigned(164,8) ,
11519	 => std_logic_vector(to_unsigned(164,8) ,
11520	 => std_logic_vector(to_unsigned(164,8) ,
11521	 => std_logic_vector(to_unsigned(116,8) ,
11522	 => std_logic_vector(to_unsigned(124,8) ,
11523	 => std_logic_vector(to_unsigned(127,8) ,
11524	 => std_logic_vector(to_unsigned(130,8) ,
11525	 => std_logic_vector(to_unsigned(134,8) ,
11526	 => std_logic_vector(to_unsigned(136,8) ,
11527	 => std_logic_vector(to_unsigned(138,8) ,
11528	 => std_logic_vector(to_unsigned(131,8) ,
11529	 => std_logic_vector(to_unsigned(130,8) ,
11530	 => std_logic_vector(to_unsigned(112,8) ,
11531	 => std_logic_vector(to_unsigned(111,8) ,
11532	 => std_logic_vector(to_unsigned(131,8) ,
11533	 => std_logic_vector(to_unsigned(134,8) ,
11534	 => std_logic_vector(to_unsigned(133,8) ,
11535	 => std_logic_vector(to_unsigned(134,8) ,
11536	 => std_logic_vector(to_unsigned(136,8) ,
11537	 => std_logic_vector(to_unsigned(133,8) ,
11538	 => std_logic_vector(to_unsigned(134,8) ,
11539	 => std_logic_vector(to_unsigned(128,8) ,
11540	 => std_logic_vector(to_unsigned(133,8) ,
11541	 => std_logic_vector(to_unsigned(133,8) ,
11542	 => std_logic_vector(to_unsigned(134,8) ,
11543	 => std_logic_vector(to_unsigned(144,8) ,
11544	 => std_logic_vector(to_unsigned(139,8) ,
11545	 => std_logic_vector(to_unsigned(138,8) ,
11546	 => std_logic_vector(to_unsigned(139,8) ,
11547	 => std_logic_vector(to_unsigned(139,8) ,
11548	 => std_logic_vector(to_unsigned(139,8) ,
11549	 => std_logic_vector(to_unsigned(125,8) ,
11550	 => std_logic_vector(to_unsigned(103,8) ,
11551	 => std_logic_vector(to_unsigned(100,8) ,
11552	 => std_logic_vector(to_unsigned(103,8) ,
11553	 => std_logic_vector(to_unsigned(97,8) ,
11554	 => std_logic_vector(to_unsigned(111,8) ,
11555	 => std_logic_vector(to_unsigned(127,8) ,
11556	 => std_logic_vector(to_unsigned(122,8) ,
11557	 => std_logic_vector(to_unsigned(121,8) ,
11558	 => std_logic_vector(to_unsigned(122,8) ,
11559	 => std_logic_vector(to_unsigned(127,8) ,
11560	 => std_logic_vector(to_unsigned(125,8) ,
11561	 => std_logic_vector(to_unsigned(128,8) ,
11562	 => std_logic_vector(to_unsigned(127,8) ,
11563	 => std_logic_vector(to_unsigned(130,8) ,
11564	 => std_logic_vector(to_unsigned(136,8) ,
11565	 => std_logic_vector(to_unsigned(141,8) ,
11566	 => std_logic_vector(to_unsigned(139,8) ,
11567	 => std_logic_vector(to_unsigned(134,8) ,
11568	 => std_logic_vector(to_unsigned(138,8) ,
11569	 => std_logic_vector(to_unsigned(131,8) ,
11570	 => std_logic_vector(to_unsigned(130,8) ,
11571	 => std_logic_vector(to_unsigned(138,8) ,
11572	 => std_logic_vector(to_unsigned(134,8) ,
11573	 => std_logic_vector(to_unsigned(142,8) ,
11574	 => std_logic_vector(to_unsigned(141,8) ,
11575	 => std_logic_vector(to_unsigned(134,8) ,
11576	 => std_logic_vector(to_unsigned(139,8) ,
11577	 => std_logic_vector(to_unsigned(138,8) ,
11578	 => std_logic_vector(to_unsigned(144,8) ,
11579	 => std_logic_vector(to_unsigned(149,8) ,
11580	 => std_logic_vector(to_unsigned(151,8) ,
11581	 => std_logic_vector(to_unsigned(146,8) ,
11582	 => std_logic_vector(to_unsigned(146,8) ,
11583	 => std_logic_vector(to_unsigned(147,8) ,
11584	 => std_logic_vector(to_unsigned(133,8) ,
11585	 => std_logic_vector(to_unsigned(116,8) ,
11586	 => std_logic_vector(to_unsigned(139,8) ,
11587	 => std_logic_vector(to_unsigned(134,8) ,
11588	 => std_logic_vector(to_unsigned(134,8) ,
11589	 => std_logic_vector(to_unsigned(133,8) ,
11590	 => std_logic_vector(to_unsigned(122,8) ,
11591	 => std_logic_vector(to_unsigned(128,8) ,
11592	 => std_logic_vector(to_unsigned(138,8) ,
11593	 => std_logic_vector(to_unsigned(139,8) ,
11594	 => std_logic_vector(to_unsigned(125,8) ,
11595	 => std_logic_vector(to_unsigned(108,8) ,
11596	 => std_logic_vector(to_unsigned(114,8) ,
11597	 => std_logic_vector(to_unsigned(130,8) ,
11598	 => std_logic_vector(to_unsigned(125,8) ,
11599	 => std_logic_vector(to_unsigned(124,8) ,
11600	 => std_logic_vector(to_unsigned(128,8) ,
11601	 => std_logic_vector(to_unsigned(134,8) ,
11602	 => std_logic_vector(to_unsigned(136,8) ,
11603	 => std_logic_vector(to_unsigned(128,8) ,
11604	 => std_logic_vector(to_unsigned(133,8) ,
11605	 => std_logic_vector(to_unsigned(142,8) ,
11606	 => std_logic_vector(to_unsigned(136,8) ,
11607	 => std_logic_vector(to_unsigned(144,8) ,
11608	 => std_logic_vector(to_unsigned(154,8) ,
11609	 => std_logic_vector(to_unsigned(151,8) ,
11610	 => std_logic_vector(to_unsigned(156,8) ,
11611	 => std_logic_vector(to_unsigned(131,8) ,
11612	 => std_logic_vector(to_unsigned(118,8) ,
11613	 => std_logic_vector(to_unsigned(124,8) ,
11614	 => std_logic_vector(to_unsigned(116,8) ,
11615	 => std_logic_vector(to_unsigned(116,8) ,
11616	 => std_logic_vector(to_unsigned(121,8) ,
11617	 => std_logic_vector(to_unsigned(114,8) ,
11618	 => std_logic_vector(to_unsigned(119,8) ,
11619	 => std_logic_vector(to_unsigned(121,8) ,
11620	 => std_logic_vector(to_unsigned(122,8) ,
11621	 => std_logic_vector(to_unsigned(134,8) ,
11622	 => std_logic_vector(to_unsigned(131,8) ,
11623	 => std_logic_vector(to_unsigned(125,8) ,
11624	 => std_logic_vector(to_unsigned(114,8) ,
11625	 => std_logic_vector(to_unsigned(107,8) ,
11626	 => std_logic_vector(to_unsigned(99,8) ,
11627	 => std_logic_vector(to_unsigned(84,8) ,
11628	 => std_logic_vector(to_unsigned(84,8) ,
11629	 => std_logic_vector(to_unsigned(92,8) ,
11630	 => std_logic_vector(to_unsigned(88,8) ,
11631	 => std_logic_vector(to_unsigned(76,8) ,
11632	 => std_logic_vector(to_unsigned(88,8) ,
11633	 => std_logic_vector(to_unsigned(96,8) ,
11634	 => std_logic_vector(to_unsigned(88,8) ,
11635	 => std_logic_vector(to_unsigned(97,8) ,
11636	 => std_logic_vector(to_unsigned(100,8) ,
11637	 => std_logic_vector(to_unsigned(101,8) ,
11638	 => std_logic_vector(to_unsigned(108,8) ,
11639	 => std_logic_vector(to_unsigned(101,8) ,
11640	 => std_logic_vector(to_unsigned(99,8) ,
11641	 => std_logic_vector(to_unsigned(115,8) ,
11642	 => std_logic_vector(to_unsigned(107,8) ,
11643	 => std_logic_vector(to_unsigned(107,8) ,
11644	 => std_logic_vector(to_unsigned(127,8) ,
11645	 => std_logic_vector(to_unsigned(125,8) ,
11646	 => std_logic_vector(to_unsigned(111,8) ,
11647	 => std_logic_vector(to_unsigned(119,8) ,
11648	 => std_logic_vector(to_unsigned(125,8) ,
11649	 => std_logic_vector(to_unsigned(118,8) ,
11650	 => std_logic_vector(to_unsigned(122,8) ,
11651	 => std_logic_vector(to_unsigned(122,8) ,
11652	 => std_logic_vector(to_unsigned(119,8) ,
11653	 => std_logic_vector(to_unsigned(111,8) ,
11654	 => std_logic_vector(to_unsigned(111,8) ,
11655	 => std_logic_vector(to_unsigned(101,8) ,
11656	 => std_logic_vector(to_unsigned(91,8) ,
11657	 => std_logic_vector(to_unsigned(86,8) ,
11658	 => std_logic_vector(to_unsigned(88,8) ,
11659	 => std_logic_vector(to_unsigned(109,8) ,
11660	 => std_logic_vector(to_unsigned(115,8) ,
11661	 => std_logic_vector(to_unsigned(115,8) ,
11662	 => std_logic_vector(to_unsigned(107,8) ,
11663	 => std_logic_vector(to_unsigned(99,8) ,
11664	 => std_logic_vector(to_unsigned(107,8) ,
11665	 => std_logic_vector(to_unsigned(100,8) ,
11666	 => std_logic_vector(to_unsigned(84,8) ,
11667	 => std_logic_vector(to_unsigned(97,8) ,
11668	 => std_logic_vector(to_unsigned(100,8) ,
11669	 => std_logic_vector(to_unsigned(88,8) ,
11670	 => std_logic_vector(to_unsigned(107,8) ,
11671	 => std_logic_vector(to_unsigned(121,8) ,
11672	 => std_logic_vector(to_unsigned(85,8) ,
11673	 => std_logic_vector(to_unsigned(79,8) ,
11674	 => std_logic_vector(to_unsigned(80,8) ,
11675	 => std_logic_vector(to_unsigned(78,8) ,
11676	 => std_logic_vector(to_unsigned(95,8) ,
11677	 => std_logic_vector(to_unsigned(97,8) ,
11678	 => std_logic_vector(to_unsigned(87,8) ,
11679	 => std_logic_vector(to_unsigned(84,8) ,
11680	 => std_logic_vector(to_unsigned(87,8) ,
11681	 => std_logic_vector(to_unsigned(101,8) ,
11682	 => std_logic_vector(to_unsigned(93,8) ,
11683	 => std_logic_vector(to_unsigned(74,8) ,
11684	 => std_logic_vector(to_unsigned(71,8) ,
11685	 => std_logic_vector(to_unsigned(68,8) ,
11686	 => std_logic_vector(to_unsigned(73,8) ,
11687	 => std_logic_vector(to_unsigned(82,8) ,
11688	 => std_logic_vector(to_unsigned(85,8) ,
11689	 => std_logic_vector(to_unsigned(84,8) ,
11690	 => std_logic_vector(to_unsigned(86,8) ,
11691	 => std_logic_vector(to_unsigned(87,8) ,
11692	 => std_logic_vector(to_unsigned(93,8) ,
11693	 => std_logic_vector(to_unsigned(96,8) ,
11694	 => std_logic_vector(to_unsigned(73,8) ,
11695	 => std_logic_vector(to_unsigned(70,8) ,
11696	 => std_logic_vector(to_unsigned(85,8) ,
11697	 => std_logic_vector(to_unsigned(76,8) ,
11698	 => std_logic_vector(to_unsigned(74,8) ,
11699	 => std_logic_vector(to_unsigned(88,8) ,
11700	 => std_logic_vector(to_unsigned(68,8) ,
11701	 => std_logic_vector(to_unsigned(62,8) ,
11702	 => std_logic_vector(to_unsigned(78,8) ,
11703	 => std_logic_vector(to_unsigned(92,8) ,
11704	 => std_logic_vector(to_unsigned(88,8) ,
11705	 => std_logic_vector(to_unsigned(103,8) ,
11706	 => std_logic_vector(to_unsigned(91,8) ,
11707	 => std_logic_vector(to_unsigned(78,8) ,
11708	 => std_logic_vector(to_unsigned(73,8) ,
11709	 => std_logic_vector(to_unsigned(78,8) ,
11710	 => std_logic_vector(to_unsigned(76,8) ,
11711	 => std_logic_vector(to_unsigned(85,8) ,
11712	 => std_logic_vector(to_unsigned(115,8) ,
11713	 => std_logic_vector(to_unsigned(109,8) ,
11714	 => std_logic_vector(to_unsigned(93,8) ,
11715	 => std_logic_vector(to_unsigned(99,8) ,
11716	 => std_logic_vector(to_unsigned(101,8) ,
11717	 => std_logic_vector(to_unsigned(99,8) ,
11718	 => std_logic_vector(to_unsigned(100,8) ,
11719	 => std_logic_vector(to_unsigned(111,8) ,
11720	 => std_logic_vector(to_unsigned(105,8) ,
11721	 => std_logic_vector(to_unsigned(107,8) ,
11722	 => std_logic_vector(to_unsigned(107,8) ,
11723	 => std_logic_vector(to_unsigned(84,8) ,
11724	 => std_logic_vector(to_unsigned(70,8) ,
11725	 => std_logic_vector(to_unsigned(93,8) ,
11726	 => std_logic_vector(to_unsigned(119,8) ,
11727	 => std_logic_vector(to_unsigned(107,8) ,
11728	 => std_logic_vector(to_unsigned(112,8) ,
11729	 => std_logic_vector(to_unsigned(111,8) ,
11730	 => std_logic_vector(to_unsigned(82,8) ,
11731	 => std_logic_vector(to_unsigned(79,8) ,
11732	 => std_logic_vector(to_unsigned(80,8) ,
11733	 => std_logic_vector(to_unsigned(76,8) ,
11734	 => std_logic_vector(to_unsigned(77,8) ,
11735	 => std_logic_vector(to_unsigned(87,8) ,
11736	 => std_logic_vector(to_unsigned(91,8) ,
11737	 => std_logic_vector(to_unsigned(96,8) ,
11738	 => std_logic_vector(to_unsigned(96,8) ,
11739	 => std_logic_vector(to_unsigned(86,8) ,
11740	 => std_logic_vector(to_unsigned(87,8) ,
11741	 => std_logic_vector(to_unsigned(87,8) ,
11742	 => std_logic_vector(to_unsigned(62,8) ,
11743	 => std_logic_vector(to_unsigned(65,8) ,
11744	 => std_logic_vector(to_unsigned(72,8) ,
11745	 => std_logic_vector(to_unsigned(65,8) ,
11746	 => std_logic_vector(to_unsigned(69,8) ,
11747	 => std_logic_vector(to_unsigned(74,8) ,
11748	 => std_logic_vector(to_unsigned(72,8) ,
11749	 => std_logic_vector(to_unsigned(67,8) ,
11750	 => std_logic_vector(to_unsigned(62,8) ,
11751	 => std_logic_vector(to_unsigned(69,8) ,
11752	 => std_logic_vector(to_unsigned(68,8) ,
11753	 => std_logic_vector(to_unsigned(76,8) ,
11754	 => std_logic_vector(to_unsigned(87,8) ,
11755	 => std_logic_vector(to_unsigned(77,8) ,
11756	 => std_logic_vector(to_unsigned(76,8) ,
11757	 => std_logic_vector(to_unsigned(61,8) ,
11758	 => std_logic_vector(to_unsigned(64,8) ,
11759	 => std_logic_vector(to_unsigned(58,8) ,
11760	 => std_logic_vector(to_unsigned(48,8) ,
11761	 => std_logic_vector(to_unsigned(53,8) ,
11762	 => std_logic_vector(to_unsigned(56,8) ,
11763	 => std_logic_vector(to_unsigned(40,8) ,
11764	 => std_logic_vector(to_unsigned(2,8) ,
11765	 => std_logic_vector(to_unsigned(0,8) ,
11766	 => std_logic_vector(to_unsigned(0,8) ,
11767	 => std_logic_vector(to_unsigned(25,8) ,
11768	 => std_logic_vector(to_unsigned(60,8) ,
11769	 => std_logic_vector(to_unsigned(52,8) ,
11770	 => std_logic_vector(to_unsigned(82,8) ,
11771	 => std_logic_vector(to_unsigned(97,8) ,
11772	 => std_logic_vector(to_unsigned(90,8) ,
11773	 => std_logic_vector(to_unsigned(81,8) ,
11774	 => std_logic_vector(to_unsigned(73,8) ,
11775	 => std_logic_vector(to_unsigned(73,8) ,
11776	 => std_logic_vector(to_unsigned(54,8) ,
11777	 => std_logic_vector(to_unsigned(44,8) ,
11778	 => std_logic_vector(to_unsigned(37,8) ,
11779	 => std_logic_vector(to_unsigned(41,8) ,
11780	 => std_logic_vector(to_unsigned(47,8) ,
11781	 => std_logic_vector(to_unsigned(41,8) ,
11782	 => std_logic_vector(to_unsigned(45,8) ,
11783	 => std_logic_vector(to_unsigned(46,8) ,
11784	 => std_logic_vector(to_unsigned(45,8) ,
11785	 => std_logic_vector(to_unsigned(46,8) ,
11786	 => std_logic_vector(to_unsigned(51,8) ,
11787	 => std_logic_vector(to_unsigned(55,8) ,
11788	 => std_logic_vector(to_unsigned(56,8) ,
11789	 => std_logic_vector(to_unsigned(72,8) ,
11790	 => std_logic_vector(to_unsigned(76,8) ,
11791	 => std_logic_vector(to_unsigned(61,8) ,
11792	 => std_logic_vector(to_unsigned(51,8) ,
11793	 => std_logic_vector(to_unsigned(53,8) ,
11794	 => std_logic_vector(to_unsigned(54,8) ,
11795	 => std_logic_vector(to_unsigned(58,8) ,
11796	 => std_logic_vector(to_unsigned(69,8) ,
11797	 => std_logic_vector(to_unsigned(68,8) ,
11798	 => std_logic_vector(to_unsigned(67,8) ,
11799	 => std_logic_vector(to_unsigned(65,8) ,
11800	 => std_logic_vector(to_unsigned(70,8) ,
11801	 => std_logic_vector(to_unsigned(85,8) ,
11802	 => std_logic_vector(to_unsigned(86,8) ,
11803	 => std_logic_vector(to_unsigned(96,8) ,
11804	 => std_logic_vector(to_unsigned(107,8) ,
11805	 => std_logic_vector(to_unsigned(82,8) ,
11806	 => std_logic_vector(to_unsigned(72,8) ,
11807	 => std_logic_vector(to_unsigned(72,8) ,
11808	 => std_logic_vector(to_unsigned(79,8) ,
11809	 => std_logic_vector(to_unsigned(91,8) ,
11810	 => std_logic_vector(to_unsigned(101,8) ,
11811	 => std_logic_vector(to_unsigned(112,8) ,
11812	 => std_logic_vector(to_unsigned(122,8) ,
11813	 => std_logic_vector(to_unsigned(131,8) ,
11814	 => std_logic_vector(to_unsigned(105,8) ,
11815	 => std_logic_vector(to_unsigned(125,8) ,
11816	 => std_logic_vector(to_unsigned(139,8) ,
11817	 => std_logic_vector(to_unsigned(109,8) ,
11818	 => std_logic_vector(to_unsigned(130,8) ,
11819	 => std_logic_vector(to_unsigned(149,8) ,
11820	 => std_logic_vector(to_unsigned(134,8) ,
11821	 => std_logic_vector(to_unsigned(149,8) ,
11822	 => std_logic_vector(to_unsigned(156,8) ,
11823	 => std_logic_vector(to_unsigned(157,8) ,
11824	 => std_logic_vector(to_unsigned(157,8) ,
11825	 => std_logic_vector(to_unsigned(161,8) ,
11826	 => std_logic_vector(to_unsigned(164,8) ,
11827	 => std_logic_vector(to_unsigned(159,8) ,
11828	 => std_logic_vector(to_unsigned(152,8) ,
11829	 => std_logic_vector(to_unsigned(151,8) ,
11830	 => std_logic_vector(to_unsigned(164,8) ,
11831	 => std_logic_vector(to_unsigned(161,8) ,
11832	 => std_logic_vector(to_unsigned(152,8) ,
11833	 => std_logic_vector(to_unsigned(156,8) ,
11834	 => std_logic_vector(to_unsigned(157,8) ,
11835	 => std_logic_vector(to_unsigned(159,8) ,
11836	 => std_logic_vector(to_unsigned(163,8) ,
11837	 => std_logic_vector(to_unsigned(161,8) ,
11838	 => std_logic_vector(to_unsigned(157,8) ,
11839	 => std_logic_vector(to_unsigned(159,8) ,
11840	 => std_logic_vector(to_unsigned(161,8) ,
11841	 => std_logic_vector(to_unsigned(127,8) ,
11842	 => std_logic_vector(to_unsigned(130,8) ,
11843	 => std_logic_vector(to_unsigned(128,8) ,
11844	 => std_logic_vector(to_unsigned(134,8) ,
11845	 => std_logic_vector(to_unsigned(139,8) ,
11846	 => std_logic_vector(to_unsigned(138,8) ,
11847	 => std_logic_vector(to_unsigned(138,8) ,
11848	 => std_logic_vector(to_unsigned(134,8) ,
11849	 => std_logic_vector(to_unsigned(138,8) ,
11850	 => std_logic_vector(to_unsigned(133,8) ,
11851	 => std_logic_vector(to_unsigned(128,8) ,
11852	 => std_logic_vector(to_unsigned(136,8) ,
11853	 => std_logic_vector(to_unsigned(144,8) ,
11854	 => std_logic_vector(to_unsigned(139,8) ,
11855	 => std_logic_vector(to_unsigned(136,8) ,
11856	 => std_logic_vector(to_unsigned(139,8) ,
11857	 => std_logic_vector(to_unsigned(141,8) ,
11858	 => std_logic_vector(to_unsigned(139,8) ,
11859	 => std_logic_vector(to_unsigned(136,8) ,
11860	 => std_logic_vector(to_unsigned(144,8) ,
11861	 => std_logic_vector(to_unsigned(146,8) ,
11862	 => std_logic_vector(to_unsigned(139,8) ,
11863	 => std_logic_vector(to_unsigned(151,8) ,
11864	 => std_logic_vector(to_unsigned(146,8) ,
11865	 => std_logic_vector(to_unsigned(144,8) ,
11866	 => std_logic_vector(to_unsigned(139,8) ,
11867	 => std_logic_vector(to_unsigned(134,8) ,
11868	 => std_logic_vector(to_unsigned(138,8) ,
11869	 => std_logic_vector(to_unsigned(116,8) ,
11870	 => std_logic_vector(to_unsigned(90,8) ,
11871	 => std_logic_vector(to_unsigned(97,8) ,
11872	 => std_logic_vector(to_unsigned(92,8) ,
11873	 => std_logic_vector(to_unsigned(87,8) ,
11874	 => std_logic_vector(to_unsigned(97,8) ,
11875	 => std_logic_vector(to_unsigned(116,8) ,
11876	 => std_logic_vector(to_unsigned(124,8) ,
11877	 => std_logic_vector(to_unsigned(111,8) ,
11878	 => std_logic_vector(to_unsigned(116,8) ,
11879	 => std_logic_vector(to_unsigned(131,8) ,
11880	 => std_logic_vector(to_unsigned(127,8) ,
11881	 => std_logic_vector(to_unsigned(133,8) ,
11882	 => std_logic_vector(to_unsigned(130,8) ,
11883	 => std_logic_vector(to_unsigned(131,8) ,
11884	 => std_logic_vector(to_unsigned(141,8) ,
11885	 => std_logic_vector(to_unsigned(136,8) ,
11886	 => std_logic_vector(to_unsigned(133,8) ,
11887	 => std_logic_vector(to_unsigned(128,8) ,
11888	 => std_logic_vector(to_unsigned(127,8) ,
11889	 => std_logic_vector(to_unsigned(114,8) ,
11890	 => std_logic_vector(to_unsigned(109,8) ,
11891	 => std_logic_vector(to_unsigned(136,8) ,
11892	 => std_logic_vector(to_unsigned(136,8) ,
11893	 => std_logic_vector(to_unsigned(144,8) ,
11894	 => std_logic_vector(to_unsigned(146,8) ,
11895	 => std_logic_vector(to_unsigned(139,8) ,
11896	 => std_logic_vector(to_unsigned(142,8) ,
11897	 => std_logic_vector(to_unsigned(144,8) ,
11898	 => std_logic_vector(to_unsigned(149,8) ,
11899	 => std_logic_vector(to_unsigned(152,8) ,
11900	 => std_logic_vector(to_unsigned(154,8) ,
11901	 => std_logic_vector(to_unsigned(136,8) ,
11902	 => std_logic_vector(to_unsigned(128,8) ,
11903	 => std_logic_vector(to_unsigned(139,8) ,
11904	 => std_logic_vector(to_unsigned(122,8) ,
11905	 => std_logic_vector(to_unsigned(118,8) ,
11906	 => std_logic_vector(to_unsigned(127,8) ,
11907	 => std_logic_vector(to_unsigned(115,8) ,
11908	 => std_logic_vector(to_unsigned(114,8) ,
11909	 => std_logic_vector(to_unsigned(121,8) ,
11910	 => std_logic_vector(to_unsigned(109,8) ,
11911	 => std_logic_vector(to_unsigned(108,8) ,
11912	 => std_logic_vector(to_unsigned(122,8) ,
11913	 => std_logic_vector(to_unsigned(127,8) ,
11914	 => std_logic_vector(to_unsigned(116,8) ,
11915	 => std_logic_vector(to_unsigned(109,8) ,
11916	 => std_logic_vector(to_unsigned(115,8) ,
11917	 => std_logic_vector(to_unsigned(118,8) ,
11918	 => std_logic_vector(to_unsigned(119,8) ,
11919	 => std_logic_vector(to_unsigned(130,8) ,
11920	 => std_logic_vector(to_unsigned(116,8) ,
11921	 => std_logic_vector(to_unsigned(125,8) ,
11922	 => std_logic_vector(to_unsigned(130,8) ,
11923	 => std_logic_vector(to_unsigned(114,8) ,
11924	 => std_logic_vector(to_unsigned(119,8) ,
11925	 => std_logic_vector(to_unsigned(124,8) ,
11926	 => std_logic_vector(to_unsigned(125,8) ,
11927	 => std_logic_vector(to_unsigned(141,8) ,
11928	 => std_logic_vector(to_unsigned(159,8) ,
11929	 => std_logic_vector(to_unsigned(147,8) ,
11930	 => std_logic_vector(to_unsigned(141,8) ,
11931	 => std_logic_vector(to_unsigned(128,8) ,
11932	 => std_logic_vector(to_unsigned(124,8) ,
11933	 => std_logic_vector(to_unsigned(124,8) ,
11934	 => std_logic_vector(to_unsigned(121,8) ,
11935	 => std_logic_vector(to_unsigned(122,8) ,
11936	 => std_logic_vector(to_unsigned(122,8) ,
11937	 => std_logic_vector(to_unsigned(122,8) ,
11938	 => std_logic_vector(to_unsigned(128,8) ,
11939	 => std_logic_vector(to_unsigned(125,8) ,
11940	 => std_logic_vector(to_unsigned(115,8) ,
11941	 => std_logic_vector(to_unsigned(119,8) ,
11942	 => std_logic_vector(to_unsigned(134,8) ,
11943	 => std_logic_vector(to_unsigned(130,8) ,
11944	 => std_logic_vector(to_unsigned(114,8) ,
11945	 => std_logic_vector(to_unsigned(103,8) ,
11946	 => std_logic_vector(to_unsigned(93,8) ,
11947	 => std_logic_vector(to_unsigned(85,8) ,
11948	 => std_logic_vector(to_unsigned(88,8) ,
11949	 => std_logic_vector(to_unsigned(105,8) ,
11950	 => std_logic_vector(to_unsigned(85,8) ,
11951	 => std_logic_vector(to_unsigned(82,8) ,
11952	 => std_logic_vector(to_unsigned(101,8) ,
11953	 => std_logic_vector(to_unsigned(112,8) ,
11954	 => std_logic_vector(to_unsigned(111,8) ,
11955	 => std_logic_vector(to_unsigned(112,8) ,
11956	 => std_logic_vector(to_unsigned(109,8) ,
11957	 => std_logic_vector(to_unsigned(112,8) ,
11958	 => std_logic_vector(to_unsigned(111,8) ,
11959	 => std_logic_vector(to_unsigned(103,8) ,
11960	 => std_logic_vector(to_unsigned(100,8) ,
11961	 => std_logic_vector(to_unsigned(109,8) ,
11962	 => std_logic_vector(to_unsigned(100,8) ,
11963	 => std_logic_vector(to_unsigned(103,8) ,
11964	 => std_logic_vector(to_unsigned(133,8) ,
11965	 => std_logic_vector(to_unsigned(124,8) ,
11966	 => std_logic_vector(to_unsigned(108,8) ,
11967	 => std_logic_vector(to_unsigned(116,8) ,
11968	 => std_logic_vector(to_unsigned(116,8) ,
11969	 => std_logic_vector(to_unsigned(114,8) ,
11970	 => std_logic_vector(to_unsigned(118,8) ,
11971	 => std_logic_vector(to_unsigned(121,8) ,
11972	 => std_logic_vector(to_unsigned(109,8) ,
11973	 => std_logic_vector(to_unsigned(92,8) ,
11974	 => std_logic_vector(to_unsigned(95,8) ,
11975	 => std_logic_vector(to_unsigned(92,8) ,
11976	 => std_logic_vector(to_unsigned(90,8) ,
11977	 => std_logic_vector(to_unsigned(88,8) ,
11978	 => std_logic_vector(to_unsigned(100,8) ,
11979	 => std_logic_vector(to_unsigned(118,8) ,
11980	 => std_logic_vector(to_unsigned(118,8) ,
11981	 => std_logic_vector(to_unsigned(115,8) ,
11982	 => std_logic_vector(to_unsigned(97,8) ,
11983	 => std_logic_vector(to_unsigned(90,8) ,
11984	 => std_logic_vector(to_unsigned(103,8) ,
11985	 => std_logic_vector(to_unsigned(103,8) ,
11986	 => std_logic_vector(to_unsigned(104,8) ,
11987	 => std_logic_vector(to_unsigned(105,8) ,
11988	 => std_logic_vector(to_unsigned(93,8) ,
11989	 => std_logic_vector(to_unsigned(95,8) ,
11990	 => std_logic_vector(to_unsigned(103,8) ,
11991	 => std_logic_vector(to_unsigned(108,8) ,
11992	 => std_logic_vector(to_unsigned(91,8) ,
11993	 => std_logic_vector(to_unsigned(87,8) ,
11994	 => std_logic_vector(to_unsigned(88,8) ,
11995	 => std_logic_vector(to_unsigned(82,8) ,
11996	 => std_logic_vector(to_unsigned(88,8) ,
11997	 => std_logic_vector(to_unsigned(96,8) ,
11998	 => std_logic_vector(to_unsigned(109,8) ,
11999	 => std_logic_vector(to_unsigned(87,8) ,
12000	 => std_logic_vector(to_unsigned(78,8) ,
12001	 => std_logic_vector(to_unsigned(91,8) ,
12002	 => std_logic_vector(to_unsigned(90,8) ,
12003	 => std_logic_vector(to_unsigned(73,8) ,
12004	 => std_logic_vector(to_unsigned(69,8) ,
12005	 => std_logic_vector(to_unsigned(63,8) ,
12006	 => std_logic_vector(to_unsigned(64,8) ,
12007	 => std_logic_vector(to_unsigned(79,8) ,
12008	 => std_logic_vector(to_unsigned(82,8) ,
12009	 => std_logic_vector(to_unsigned(79,8) ,
12010	 => std_logic_vector(to_unsigned(87,8) ,
12011	 => std_logic_vector(to_unsigned(84,8) ,
12012	 => std_logic_vector(to_unsigned(80,8) ,
12013	 => std_logic_vector(to_unsigned(97,8) ,
12014	 => std_logic_vector(to_unsigned(79,8) ,
12015	 => std_logic_vector(to_unsigned(71,8) ,
12016	 => std_logic_vector(to_unsigned(86,8) ,
12017	 => std_logic_vector(to_unsigned(79,8) ,
12018	 => std_logic_vector(to_unsigned(74,8) ,
12019	 => std_logic_vector(to_unsigned(86,8) ,
12020	 => std_logic_vector(to_unsigned(70,8) ,
12021	 => std_logic_vector(to_unsigned(66,8) ,
12022	 => std_logic_vector(to_unsigned(86,8) ,
12023	 => std_logic_vector(to_unsigned(103,8) ,
12024	 => std_logic_vector(to_unsigned(86,8) ,
12025	 => std_logic_vector(to_unsigned(84,8) ,
12026	 => std_logic_vector(to_unsigned(80,8) ,
12027	 => std_logic_vector(to_unsigned(77,8) ,
12028	 => std_logic_vector(to_unsigned(73,8) ,
12029	 => std_logic_vector(to_unsigned(77,8) ,
12030	 => std_logic_vector(to_unsigned(81,8) ,
12031	 => std_logic_vector(to_unsigned(77,8) ,
12032	 => std_logic_vector(to_unsigned(78,8) ,
12033	 => std_logic_vector(to_unsigned(91,8) ,
12034	 => std_logic_vector(to_unsigned(103,8) ,
12035	 => std_logic_vector(to_unsigned(99,8) ,
12036	 => std_logic_vector(to_unsigned(105,8) ,
12037	 => std_logic_vector(to_unsigned(105,8) ,
12038	 => std_logic_vector(to_unsigned(99,8) ,
12039	 => std_logic_vector(to_unsigned(112,8) ,
12040	 => std_logic_vector(to_unsigned(111,8) ,
12041	 => std_logic_vector(to_unsigned(108,8) ,
12042	 => std_logic_vector(to_unsigned(105,8) ,
12043	 => std_logic_vector(to_unsigned(76,8) ,
12044	 => std_logic_vector(to_unsigned(71,8) ,
12045	 => std_logic_vector(to_unsigned(92,8) ,
12046	 => std_logic_vector(to_unsigned(109,8) ,
12047	 => std_logic_vector(to_unsigned(109,8) ,
12048	 => std_logic_vector(to_unsigned(115,8) ,
12049	 => std_logic_vector(to_unsigned(108,8) ,
12050	 => std_logic_vector(to_unsigned(81,8) ,
12051	 => std_logic_vector(to_unsigned(78,8) ,
12052	 => std_logic_vector(to_unsigned(78,8) ,
12053	 => std_logic_vector(to_unsigned(76,8) ,
12054	 => std_logic_vector(to_unsigned(77,8) ,
12055	 => std_logic_vector(to_unsigned(86,8) ,
12056	 => std_logic_vector(to_unsigned(93,8) ,
12057	 => std_logic_vector(to_unsigned(101,8) ,
12058	 => std_logic_vector(to_unsigned(97,8) ,
12059	 => std_logic_vector(to_unsigned(97,8) ,
12060	 => std_logic_vector(to_unsigned(92,8) ,
12061	 => std_logic_vector(to_unsigned(92,8) ,
12062	 => std_logic_vector(to_unsigned(76,8) ,
12063	 => std_logic_vector(to_unsigned(80,8) ,
12064	 => std_logic_vector(to_unsigned(79,8) ,
12065	 => std_logic_vector(to_unsigned(71,8) ,
12066	 => std_logic_vector(to_unsigned(76,8) ,
12067	 => std_logic_vector(to_unsigned(76,8) ,
12068	 => std_logic_vector(to_unsigned(72,8) ,
12069	 => std_logic_vector(to_unsigned(68,8) ,
12070	 => std_logic_vector(to_unsigned(67,8) ,
12071	 => std_logic_vector(to_unsigned(76,8) ,
12072	 => std_logic_vector(to_unsigned(76,8) ,
12073	 => std_logic_vector(to_unsigned(84,8) ,
12074	 => std_logic_vector(to_unsigned(87,8) ,
12075	 => std_logic_vector(to_unsigned(76,8) ,
12076	 => std_logic_vector(to_unsigned(80,8) ,
12077	 => std_logic_vector(to_unsigned(67,8) ,
12078	 => std_logic_vector(to_unsigned(57,8) ,
12079	 => std_logic_vector(to_unsigned(52,8) ,
12080	 => std_logic_vector(to_unsigned(46,8) ,
12081	 => std_logic_vector(to_unsigned(55,8) ,
12082	 => std_logic_vector(to_unsigned(54,8) ,
12083	 => std_logic_vector(to_unsigned(53,8) ,
12084	 => std_logic_vector(to_unsigned(6,8) ,
12085	 => std_logic_vector(to_unsigned(0,8) ,
12086	 => std_logic_vector(to_unsigned(0,8) ,
12087	 => std_logic_vector(to_unsigned(16,8) ,
12088	 => std_logic_vector(to_unsigned(64,8) ,
12089	 => std_logic_vector(to_unsigned(62,8) ,
12090	 => std_logic_vector(to_unsigned(91,8) ,
12091	 => std_logic_vector(to_unsigned(97,8) ,
12092	 => std_logic_vector(to_unsigned(80,8) ,
12093	 => std_logic_vector(to_unsigned(76,8) ,
12094	 => std_logic_vector(to_unsigned(68,8) ,
12095	 => std_logic_vector(to_unsigned(51,8) ,
12096	 => std_logic_vector(to_unsigned(43,8) ,
12097	 => std_logic_vector(to_unsigned(44,8) ,
12098	 => std_logic_vector(to_unsigned(44,8) ,
12099	 => std_logic_vector(to_unsigned(47,8) ,
12100	 => std_logic_vector(to_unsigned(45,8) ,
12101	 => std_logic_vector(to_unsigned(40,8) ,
12102	 => std_logic_vector(to_unsigned(48,8) ,
12103	 => std_logic_vector(to_unsigned(47,8) ,
12104	 => std_logic_vector(to_unsigned(51,8) ,
12105	 => std_logic_vector(to_unsigned(52,8) ,
12106	 => std_logic_vector(to_unsigned(50,8) ,
12107	 => std_logic_vector(to_unsigned(49,8) ,
12108	 => std_logic_vector(to_unsigned(47,8) ,
12109	 => std_logic_vector(to_unsigned(63,8) ,
12110	 => std_logic_vector(to_unsigned(65,8) ,
12111	 => std_logic_vector(to_unsigned(57,8) ,
12112	 => std_logic_vector(to_unsigned(56,8) ,
12113	 => std_logic_vector(to_unsigned(56,8) ,
12114	 => std_logic_vector(to_unsigned(55,8) ,
12115	 => std_logic_vector(to_unsigned(59,8) ,
12116	 => std_logic_vector(to_unsigned(63,8) ,
12117	 => std_logic_vector(to_unsigned(62,8) ,
12118	 => std_logic_vector(to_unsigned(72,8) ,
12119	 => std_logic_vector(to_unsigned(72,8) ,
12120	 => std_logic_vector(to_unsigned(69,8) ,
12121	 => std_logic_vector(to_unsigned(78,8) ,
12122	 => std_logic_vector(to_unsigned(82,8) ,
12123	 => std_logic_vector(to_unsigned(91,8) ,
12124	 => std_logic_vector(to_unsigned(86,8) ,
12125	 => std_logic_vector(to_unsigned(73,8) ,
12126	 => std_logic_vector(to_unsigned(76,8) ,
12127	 => std_logic_vector(to_unsigned(78,8) ,
12128	 => std_logic_vector(to_unsigned(78,8) ,
12129	 => std_logic_vector(to_unsigned(78,8) ,
12130	 => std_logic_vector(to_unsigned(81,8) ,
12131	 => std_logic_vector(to_unsigned(84,8) ,
12132	 => std_logic_vector(to_unsigned(87,8) ,
12133	 => std_logic_vector(to_unsigned(97,8) ,
12134	 => std_logic_vector(to_unsigned(92,8) ,
12135	 => std_logic_vector(to_unsigned(105,8) ,
12136	 => std_logic_vector(to_unsigned(100,8) ,
12137	 => std_logic_vector(to_unsigned(85,8) ,
12138	 => std_logic_vector(to_unsigned(99,8) ,
12139	 => std_logic_vector(to_unsigned(114,8) ,
12140	 => std_logic_vector(to_unsigned(108,8) ,
12141	 => std_logic_vector(to_unsigned(122,8) ,
12142	 => std_logic_vector(to_unsigned(124,8) ,
12143	 => std_logic_vector(to_unsigned(128,8) ,
12144	 => std_logic_vector(to_unsigned(130,8) ,
12145	 => std_logic_vector(to_unsigned(142,8) ,
12146	 => std_logic_vector(to_unsigned(163,8) ,
12147	 => std_logic_vector(to_unsigned(157,8) ,
12148	 => std_logic_vector(to_unsigned(136,8) ,
12149	 => std_logic_vector(to_unsigned(149,8) ,
12150	 => std_logic_vector(to_unsigned(166,8) ,
12151	 => std_logic_vector(to_unsigned(151,8) ,
12152	 => std_logic_vector(to_unsigned(127,8) ,
12153	 => std_logic_vector(to_unsigned(131,8) ,
12154	 => std_logic_vector(to_unsigned(139,8) ,
12155	 => std_logic_vector(to_unsigned(144,8) ,
12156	 => std_logic_vector(to_unsigned(161,8) ,
12157	 => std_logic_vector(to_unsigned(159,8) ,
12158	 => std_logic_vector(to_unsigned(144,8) ,
12159	 => std_logic_vector(to_unsigned(144,8) ,
12160	 => std_logic_vector(to_unsigned(149,8) ,
12161	 => std_logic_vector(to_unsigned(134,8) ,
12162	 => std_logic_vector(to_unsigned(133,8) ,
12163	 => std_logic_vector(to_unsigned(138,8) ,
12164	 => std_logic_vector(to_unsigned(138,8) ,
12165	 => std_logic_vector(to_unsigned(139,8) ,
12166	 => std_logic_vector(to_unsigned(141,8) ,
12167	 => std_logic_vector(to_unsigned(139,8) ,
12168	 => std_logic_vector(to_unsigned(139,8) ,
12169	 => std_logic_vector(to_unsigned(133,8) ,
12170	 => std_logic_vector(to_unsigned(142,8) ,
12171	 => std_logic_vector(to_unsigned(142,8) ,
12172	 => std_logic_vector(to_unsigned(138,8) ,
12173	 => std_logic_vector(to_unsigned(149,8) ,
12174	 => std_logic_vector(to_unsigned(152,8) ,
12175	 => std_logic_vector(to_unsigned(147,8) ,
12176	 => std_logic_vector(to_unsigned(146,8) ,
12177	 => std_logic_vector(to_unsigned(147,8) ,
12178	 => std_logic_vector(to_unsigned(149,8) ,
12179	 => std_logic_vector(to_unsigned(151,8) ,
12180	 => std_logic_vector(to_unsigned(151,8) ,
12181	 => std_logic_vector(to_unsigned(147,8) ,
12182	 => std_logic_vector(to_unsigned(147,8) ,
12183	 => std_logic_vector(to_unsigned(156,8) ,
12184	 => std_logic_vector(to_unsigned(154,8) ,
12185	 => std_logic_vector(to_unsigned(154,8) ,
12186	 => std_logic_vector(to_unsigned(151,8) ,
12187	 => std_logic_vector(to_unsigned(144,8) ,
12188	 => std_logic_vector(to_unsigned(141,8) ,
12189	 => std_logic_vector(to_unsigned(114,8) ,
12190	 => std_logic_vector(to_unsigned(97,8) ,
12191	 => std_logic_vector(to_unsigned(104,8) ,
12192	 => std_logic_vector(to_unsigned(95,8) ,
12193	 => std_logic_vector(to_unsigned(96,8) ,
12194	 => std_logic_vector(to_unsigned(91,8) ,
12195	 => std_logic_vector(to_unsigned(105,8) ,
12196	 => std_logic_vector(to_unsigned(133,8) ,
12197	 => std_logic_vector(to_unsigned(104,8) ,
12198	 => std_logic_vector(to_unsigned(109,8) ,
12199	 => std_logic_vector(to_unsigned(131,8) ,
12200	 => std_logic_vector(to_unsigned(128,8) ,
12201	 => std_logic_vector(to_unsigned(133,8) ,
12202	 => std_logic_vector(to_unsigned(134,8) ,
12203	 => std_logic_vector(to_unsigned(127,8) ,
12204	 => std_logic_vector(to_unsigned(124,8) ,
12205	 => std_logic_vector(to_unsigned(116,8) ,
12206	 => std_logic_vector(to_unsigned(116,8) ,
12207	 => std_logic_vector(to_unsigned(116,8) ,
12208	 => std_logic_vector(to_unsigned(114,8) ,
12209	 => std_logic_vector(to_unsigned(112,8) ,
12210	 => std_logic_vector(to_unsigned(118,8) ,
12211	 => std_logic_vector(to_unsigned(131,8) ,
12212	 => std_logic_vector(to_unsigned(139,8) ,
12213	 => std_logic_vector(to_unsigned(127,8) ,
12214	 => std_logic_vector(to_unsigned(119,8) ,
12215	 => std_logic_vector(to_unsigned(138,8) ,
12216	 => std_logic_vector(to_unsigned(152,8) ,
12217	 => std_logic_vector(to_unsigned(147,8) ,
12218	 => std_logic_vector(to_unsigned(154,8) ,
12219	 => std_logic_vector(to_unsigned(151,8) ,
12220	 => std_logic_vector(to_unsigned(147,8) ,
12221	 => std_logic_vector(to_unsigned(139,8) ,
12222	 => std_logic_vector(to_unsigned(121,8) ,
12223	 => std_logic_vector(to_unsigned(127,8) ,
12224	 => std_logic_vector(to_unsigned(124,8) ,
12225	 => std_logic_vector(to_unsigned(130,8) ,
12226	 => std_logic_vector(to_unsigned(125,8) ,
12227	 => std_logic_vector(to_unsigned(115,8) ,
12228	 => std_logic_vector(to_unsigned(115,8) ,
12229	 => std_logic_vector(to_unsigned(112,8) ,
12230	 => std_logic_vector(to_unsigned(116,8) ,
12231	 => std_logic_vector(to_unsigned(122,8) ,
12232	 => std_logic_vector(to_unsigned(116,8) ,
12233	 => std_logic_vector(to_unsigned(124,8) ,
12234	 => std_logic_vector(to_unsigned(138,8) ,
12235	 => std_logic_vector(to_unsigned(139,8) ,
12236	 => std_logic_vector(to_unsigned(125,8) ,
12237	 => std_logic_vector(to_unsigned(114,8) ,
12238	 => std_logic_vector(to_unsigned(124,8) ,
12239	 => std_logic_vector(to_unsigned(131,8) ,
12240	 => std_logic_vector(to_unsigned(128,8) ,
12241	 => std_logic_vector(to_unsigned(141,8) ,
12242	 => std_logic_vector(to_unsigned(130,8) ,
12243	 => std_logic_vector(to_unsigned(116,8) ,
12244	 => std_logic_vector(to_unsigned(127,8) ,
12245	 => std_logic_vector(to_unsigned(134,8) ,
12246	 => std_logic_vector(to_unsigned(133,8) ,
12247	 => std_logic_vector(to_unsigned(128,8) ,
12248	 => std_logic_vector(to_unsigned(125,8) ,
12249	 => std_logic_vector(to_unsigned(121,8) ,
12250	 => std_logic_vector(to_unsigned(125,8) ,
12251	 => std_logic_vector(to_unsigned(127,8) ,
12252	 => std_logic_vector(to_unsigned(133,8) ,
12253	 => std_logic_vector(to_unsigned(130,8) ,
12254	 => std_logic_vector(to_unsigned(130,8) ,
12255	 => std_logic_vector(to_unsigned(125,8) ,
12256	 => std_logic_vector(to_unsigned(122,8) ,
12257	 => std_logic_vector(to_unsigned(121,8) ,
12258	 => std_logic_vector(to_unsigned(125,8) ,
12259	 => std_logic_vector(to_unsigned(131,8) ,
12260	 => std_logic_vector(to_unsigned(130,8) ,
12261	 => std_logic_vector(to_unsigned(127,8) ,
12262	 => std_logic_vector(to_unsigned(130,8) ,
12263	 => std_logic_vector(to_unsigned(130,8) ,
12264	 => std_logic_vector(to_unsigned(119,8) ,
12265	 => std_logic_vector(to_unsigned(104,8) ,
12266	 => std_logic_vector(to_unsigned(101,8) ,
12267	 => std_logic_vector(to_unsigned(90,8) ,
12268	 => std_logic_vector(to_unsigned(87,8) ,
12269	 => std_logic_vector(to_unsigned(95,8) ,
12270	 => std_logic_vector(to_unsigned(82,8) ,
12271	 => std_logic_vector(to_unsigned(90,8) ,
12272	 => std_logic_vector(to_unsigned(97,8) ,
12273	 => std_logic_vector(to_unsigned(108,8) ,
12274	 => std_logic_vector(to_unsigned(111,8) ,
12275	 => std_logic_vector(to_unsigned(121,8) ,
12276	 => std_logic_vector(to_unsigned(130,8) ,
12277	 => std_logic_vector(to_unsigned(116,8) ,
12278	 => std_logic_vector(to_unsigned(99,8) ,
12279	 => std_logic_vector(to_unsigned(95,8) ,
12280	 => std_logic_vector(to_unsigned(99,8) ,
12281	 => std_logic_vector(to_unsigned(108,8) ,
12282	 => std_logic_vector(to_unsigned(107,8) ,
12283	 => std_logic_vector(to_unsigned(109,8) ,
12284	 => std_logic_vector(to_unsigned(131,8) ,
12285	 => std_logic_vector(to_unsigned(127,8) ,
12286	 => std_logic_vector(to_unsigned(118,8) ,
12287	 => std_logic_vector(to_unsigned(115,8) ,
12288	 => std_logic_vector(to_unsigned(109,8) ,
12289	 => std_logic_vector(to_unsigned(109,8) ,
12290	 => std_logic_vector(to_unsigned(118,8) ,
12291	 => std_logic_vector(to_unsigned(125,8) ,
12292	 => std_logic_vector(to_unsigned(115,8) ,
12293	 => std_logic_vector(to_unsigned(99,8) ,
12294	 => std_logic_vector(to_unsigned(96,8) ,
12295	 => std_logic_vector(to_unsigned(93,8) ,
12296	 => std_logic_vector(to_unsigned(91,8) ,
12297	 => std_logic_vector(to_unsigned(99,8) ,
12298	 => std_logic_vector(to_unsigned(107,8) ,
12299	 => std_logic_vector(to_unsigned(116,8) ,
12300	 => std_logic_vector(to_unsigned(122,8) ,
12301	 => std_logic_vector(to_unsigned(119,8) ,
12302	 => std_logic_vector(to_unsigned(96,8) ,
12303	 => std_logic_vector(to_unsigned(87,8) ,
12304	 => std_logic_vector(to_unsigned(111,8) ,
12305	 => std_logic_vector(to_unsigned(109,8) ,
12306	 => std_logic_vector(to_unsigned(112,8) ,
12307	 => std_logic_vector(to_unsigned(115,8) ,
12308	 => std_logic_vector(to_unsigned(95,8) ,
12309	 => std_logic_vector(to_unsigned(91,8) ,
12310	 => std_logic_vector(to_unsigned(93,8) ,
12311	 => std_logic_vector(to_unsigned(88,8) ,
12312	 => std_logic_vector(to_unsigned(91,8) ,
12313	 => std_logic_vector(to_unsigned(101,8) ,
12314	 => std_logic_vector(to_unsigned(92,8) ,
12315	 => std_logic_vector(to_unsigned(91,8) ,
12316	 => std_logic_vector(to_unsigned(103,8) ,
12317	 => std_logic_vector(to_unsigned(103,8) ,
12318	 => std_logic_vector(to_unsigned(114,8) ,
12319	 => std_logic_vector(to_unsigned(85,8) ,
12320	 => std_logic_vector(to_unsigned(72,8) ,
12321	 => std_logic_vector(to_unsigned(88,8) ,
12322	 => std_logic_vector(to_unsigned(91,8) ,
12323	 => std_logic_vector(to_unsigned(72,8) ,
12324	 => std_logic_vector(to_unsigned(74,8) ,
12325	 => std_logic_vector(to_unsigned(76,8) ,
12326	 => std_logic_vector(to_unsigned(73,8) ,
12327	 => std_logic_vector(to_unsigned(82,8) ,
12328	 => std_logic_vector(to_unsigned(90,8) ,
12329	 => std_logic_vector(to_unsigned(92,8) ,
12330	 => std_logic_vector(to_unsigned(93,8) ,
12331	 => std_logic_vector(to_unsigned(82,8) ,
12332	 => std_logic_vector(to_unsigned(70,8) ,
12333	 => std_logic_vector(to_unsigned(90,8) ,
12334	 => std_logic_vector(to_unsigned(81,8) ,
12335	 => std_logic_vector(to_unsigned(72,8) ,
12336	 => std_logic_vector(to_unsigned(87,8) ,
12337	 => std_logic_vector(to_unsigned(84,8) ,
12338	 => std_logic_vector(to_unsigned(78,8) ,
12339	 => std_logic_vector(to_unsigned(81,8) ,
12340	 => std_logic_vector(to_unsigned(65,8) ,
12341	 => std_logic_vector(to_unsigned(67,8) ,
12342	 => std_logic_vector(to_unsigned(86,8) ,
12343	 => std_logic_vector(to_unsigned(92,8) ,
12344	 => std_logic_vector(to_unsigned(76,8) ,
12345	 => std_logic_vector(to_unsigned(71,8) ,
12346	 => std_logic_vector(to_unsigned(77,8) ,
12347	 => std_logic_vector(to_unsigned(77,8) ,
12348	 => std_logic_vector(to_unsigned(77,8) ,
12349	 => std_logic_vector(to_unsigned(72,8) ,
12350	 => std_logic_vector(to_unsigned(82,8) ,
12351	 => std_logic_vector(to_unsigned(72,8) ,
12352	 => std_logic_vector(to_unsigned(64,8) ,
12353	 => std_logic_vector(to_unsigned(73,8) ,
12354	 => std_logic_vector(to_unsigned(95,8) ,
12355	 => std_logic_vector(to_unsigned(95,8) ,
12356	 => std_logic_vector(to_unsigned(103,8) ,
12357	 => std_logic_vector(to_unsigned(105,8) ,
12358	 => std_logic_vector(to_unsigned(100,8) ,
12359	 => std_logic_vector(to_unsigned(112,8) ,
12360	 => std_logic_vector(to_unsigned(114,8) ,
12361	 => std_logic_vector(to_unsigned(114,8) ,
12362	 => std_logic_vector(to_unsigned(107,8) ,
12363	 => std_logic_vector(to_unsigned(73,8) ,
12364	 => std_logic_vector(to_unsigned(66,8) ,
12365	 => std_logic_vector(to_unsigned(90,8) ,
12366	 => std_logic_vector(to_unsigned(104,8) ,
12367	 => std_logic_vector(to_unsigned(105,8) ,
12368	 => std_logic_vector(to_unsigned(119,8) ,
12369	 => std_logic_vector(to_unsigned(100,8) ,
12370	 => std_logic_vector(to_unsigned(70,8) ,
12371	 => std_logic_vector(to_unsigned(74,8) ,
12372	 => std_logic_vector(to_unsigned(77,8) ,
12373	 => std_logic_vector(to_unsigned(70,8) ,
12374	 => std_logic_vector(to_unsigned(76,8) ,
12375	 => std_logic_vector(to_unsigned(95,8) ,
12376	 => std_logic_vector(to_unsigned(111,8) ,
12377	 => std_logic_vector(to_unsigned(105,8) ,
12378	 => std_logic_vector(to_unsigned(107,8) ,
12379	 => std_logic_vector(to_unsigned(104,8) ,
12380	 => std_logic_vector(to_unsigned(91,8) ,
12381	 => std_logic_vector(to_unsigned(93,8) ,
12382	 => std_logic_vector(to_unsigned(87,8) ,
12383	 => std_logic_vector(to_unsigned(92,8) ,
12384	 => std_logic_vector(to_unsigned(80,8) ,
12385	 => std_logic_vector(to_unsigned(77,8) ,
12386	 => std_logic_vector(to_unsigned(73,8) ,
12387	 => std_logic_vector(to_unsigned(74,8) ,
12388	 => std_logic_vector(to_unsigned(78,8) ,
12389	 => std_logic_vector(to_unsigned(72,8) ,
12390	 => std_logic_vector(to_unsigned(74,8) ,
12391	 => std_logic_vector(to_unsigned(72,8) ,
12392	 => std_logic_vector(to_unsigned(73,8) ,
12393	 => std_logic_vector(to_unsigned(80,8) ,
12394	 => std_logic_vector(to_unsigned(82,8) ,
12395	 => std_logic_vector(to_unsigned(85,8) ,
12396	 => std_logic_vector(to_unsigned(85,8) ,
12397	 => std_logic_vector(to_unsigned(73,8) ,
12398	 => std_logic_vector(to_unsigned(65,8) ,
12399	 => std_logic_vector(to_unsigned(54,8) ,
12400	 => std_logic_vector(to_unsigned(49,8) ,
12401	 => std_logic_vector(to_unsigned(62,8) ,
12402	 => std_logic_vector(to_unsigned(55,8) ,
12403	 => std_logic_vector(to_unsigned(70,8) ,
12404	 => std_logic_vector(to_unsigned(30,8) ,
12405	 => std_logic_vector(to_unsigned(1,8) ,
12406	 => std_logic_vector(to_unsigned(0,8) ,
12407	 => std_logic_vector(to_unsigned(5,8) ,
12408	 => std_logic_vector(to_unsigned(45,8) ,
12409	 => std_logic_vector(to_unsigned(49,8) ,
12410	 => std_logic_vector(to_unsigned(61,8) ,
12411	 => std_logic_vector(to_unsigned(63,8) ,
12412	 => std_logic_vector(to_unsigned(47,8) ,
12413	 => std_logic_vector(to_unsigned(45,8) ,
12414	 => std_logic_vector(to_unsigned(51,8) ,
12415	 => std_logic_vector(to_unsigned(49,8) ,
12416	 => std_logic_vector(to_unsigned(45,8) ,
12417	 => std_logic_vector(to_unsigned(47,8) ,
12418	 => std_logic_vector(to_unsigned(49,8) ,
12419	 => std_logic_vector(to_unsigned(43,8) ,
12420	 => std_logic_vector(to_unsigned(41,8) ,
12421	 => std_logic_vector(to_unsigned(44,8) ,
12422	 => std_logic_vector(to_unsigned(47,8) ,
12423	 => std_logic_vector(to_unsigned(46,8) ,
12424	 => std_logic_vector(to_unsigned(52,8) ,
12425	 => std_logic_vector(to_unsigned(58,8) ,
12426	 => std_logic_vector(to_unsigned(52,8) ,
12427	 => std_logic_vector(to_unsigned(50,8) ,
12428	 => std_logic_vector(to_unsigned(54,8) ,
12429	 => std_logic_vector(to_unsigned(54,8) ,
12430	 => std_logic_vector(to_unsigned(51,8) ,
12431	 => std_logic_vector(to_unsigned(50,8) ,
12432	 => std_logic_vector(to_unsigned(51,8) ,
12433	 => std_logic_vector(to_unsigned(62,8) ,
12434	 => std_logic_vector(to_unsigned(61,8) ,
12435	 => std_logic_vector(to_unsigned(63,8) ,
12436	 => std_logic_vector(to_unsigned(70,8) ,
12437	 => std_logic_vector(to_unsigned(76,8) ,
12438	 => std_logic_vector(to_unsigned(77,8) ,
12439	 => std_logic_vector(to_unsigned(80,8) ,
12440	 => std_logic_vector(to_unsigned(81,8) ,
12441	 => std_logic_vector(to_unsigned(78,8) ,
12442	 => std_logic_vector(to_unsigned(82,8) ,
12443	 => std_logic_vector(to_unsigned(87,8) ,
12444	 => std_logic_vector(to_unsigned(90,8) ,
12445	 => std_logic_vector(to_unsigned(79,8) ,
12446	 => std_logic_vector(to_unsigned(77,8) ,
12447	 => std_logic_vector(to_unsigned(81,8) ,
12448	 => std_logic_vector(to_unsigned(79,8) ,
12449	 => std_logic_vector(to_unsigned(73,8) ,
12450	 => std_logic_vector(to_unsigned(82,8) ,
12451	 => std_logic_vector(to_unsigned(92,8) ,
12452	 => std_logic_vector(to_unsigned(82,8) ,
12453	 => std_logic_vector(to_unsigned(90,8) ,
12454	 => std_logic_vector(to_unsigned(95,8) ,
12455	 => std_logic_vector(to_unsigned(91,8) ,
12456	 => std_logic_vector(to_unsigned(91,8) ,
12457	 => std_logic_vector(to_unsigned(99,8) ,
12458	 => std_logic_vector(to_unsigned(105,8) ,
12459	 => std_logic_vector(to_unsigned(108,8) ,
12460	 => std_logic_vector(to_unsigned(114,8) ,
12461	 => std_logic_vector(to_unsigned(109,8) ,
12462	 => std_logic_vector(to_unsigned(116,8) ,
12463	 => std_logic_vector(to_unsigned(127,8) ,
12464	 => std_logic_vector(to_unsigned(115,8) ,
12465	 => std_logic_vector(to_unsigned(125,8) ,
12466	 => std_logic_vector(to_unsigned(144,8) ,
12467	 => std_logic_vector(to_unsigned(147,8) ,
12468	 => std_logic_vector(to_unsigned(142,8) ,
12469	 => std_logic_vector(to_unsigned(144,8) ,
12470	 => std_logic_vector(to_unsigned(154,8) ,
12471	 => std_logic_vector(to_unsigned(139,8) ,
12472	 => std_logic_vector(to_unsigned(119,8) ,
12473	 => std_logic_vector(to_unsigned(119,8) ,
12474	 => std_logic_vector(to_unsigned(124,8) ,
12475	 => std_logic_vector(to_unsigned(133,8) ,
12476	 => std_logic_vector(to_unsigned(147,8) ,
12477	 => std_logic_vector(to_unsigned(144,8) ,
12478	 => std_logic_vector(to_unsigned(144,8) ,
12479	 => std_logic_vector(to_unsigned(147,8) ,
12480	 => std_logic_vector(to_unsigned(146,8) ,
12481	 => std_logic_vector(to_unsigned(136,8) ,
12482	 => std_logic_vector(to_unsigned(138,8) ,
12483	 => std_logic_vector(to_unsigned(144,8) ,
12484	 => std_logic_vector(to_unsigned(138,8) ,
12485	 => std_logic_vector(to_unsigned(141,8) ,
12486	 => std_logic_vector(to_unsigned(146,8) ,
12487	 => std_logic_vector(to_unsigned(142,8) ,
12488	 => std_logic_vector(to_unsigned(149,8) ,
12489	 => std_logic_vector(to_unsigned(122,8) ,
12490	 => std_logic_vector(to_unsigned(130,8) ,
12491	 => std_logic_vector(to_unsigned(151,8) ,
12492	 => std_logic_vector(to_unsigned(147,8) ,
12493	 => std_logic_vector(to_unsigned(151,8) ,
12494	 => std_logic_vector(to_unsigned(156,8) ,
12495	 => std_logic_vector(to_unsigned(156,8) ,
12496	 => std_logic_vector(to_unsigned(151,8) ,
12497	 => std_logic_vector(to_unsigned(151,8) ,
12498	 => std_logic_vector(to_unsigned(152,8) ,
12499	 => std_logic_vector(to_unsigned(157,8) ,
12500	 => std_logic_vector(to_unsigned(154,8) ,
12501	 => std_logic_vector(to_unsigned(151,8) ,
12502	 => std_logic_vector(to_unsigned(152,8) ,
12503	 => std_logic_vector(to_unsigned(156,8) ,
12504	 => std_logic_vector(to_unsigned(154,8) ,
12505	 => std_logic_vector(to_unsigned(152,8) ,
12506	 => std_logic_vector(to_unsigned(151,8) ,
12507	 => std_logic_vector(to_unsigned(156,8) ,
12508	 => std_logic_vector(to_unsigned(149,8) ,
12509	 => std_logic_vector(to_unsigned(128,8) ,
12510	 => std_logic_vector(to_unsigned(115,8) ,
12511	 => std_logic_vector(to_unsigned(107,8) ,
12512	 => std_logic_vector(to_unsigned(103,8) ,
12513	 => std_logic_vector(to_unsigned(112,8) ,
12514	 => std_logic_vector(to_unsigned(104,8) ,
12515	 => std_logic_vector(to_unsigned(108,8) ,
12516	 => std_logic_vector(to_unsigned(121,8) ,
12517	 => std_logic_vector(to_unsigned(105,8) ,
12518	 => std_logic_vector(to_unsigned(116,8) ,
12519	 => std_logic_vector(to_unsigned(139,8) ,
12520	 => std_logic_vector(to_unsigned(136,8) ,
12521	 => std_logic_vector(to_unsigned(136,8) ,
12522	 => std_logic_vector(to_unsigned(138,8) ,
12523	 => std_logic_vector(to_unsigned(119,8) ,
12524	 => std_logic_vector(to_unsigned(112,8) ,
12525	 => std_logic_vector(to_unsigned(116,8) ,
12526	 => std_logic_vector(to_unsigned(116,8) ,
12527	 => std_logic_vector(to_unsigned(116,8) ,
12528	 => std_logic_vector(to_unsigned(109,8) ,
12529	 => std_logic_vector(to_unsigned(119,8) ,
12530	 => std_logic_vector(to_unsigned(130,8) ,
12531	 => std_logic_vector(to_unsigned(124,8) ,
12532	 => std_logic_vector(to_unsigned(124,8) ,
12533	 => std_logic_vector(to_unsigned(107,8) ,
12534	 => std_logic_vector(to_unsigned(99,8) ,
12535	 => std_logic_vector(to_unsigned(128,8) ,
12536	 => std_logic_vector(to_unsigned(141,8) ,
12537	 => std_logic_vector(to_unsigned(128,8) ,
12538	 => std_logic_vector(to_unsigned(130,8) ,
12539	 => std_logic_vector(to_unsigned(133,8) ,
12540	 => std_logic_vector(to_unsigned(138,8) ,
12541	 => std_logic_vector(to_unsigned(133,8) ,
12542	 => std_logic_vector(to_unsigned(119,8) ,
12543	 => std_logic_vector(to_unsigned(128,8) ,
12544	 => std_logic_vector(to_unsigned(138,8) ,
12545	 => std_logic_vector(to_unsigned(134,8) ,
12546	 => std_logic_vector(to_unsigned(134,8) ,
12547	 => std_logic_vector(to_unsigned(139,8) ,
12548	 => std_logic_vector(to_unsigned(133,8) ,
12549	 => std_logic_vector(to_unsigned(114,8) ,
12550	 => std_logic_vector(to_unsigned(127,8) ,
12551	 => std_logic_vector(to_unsigned(147,8) ,
12552	 => std_logic_vector(to_unsigned(144,8) ,
12553	 => std_logic_vector(to_unsigned(134,8) ,
12554	 => std_logic_vector(to_unsigned(139,8) ,
12555	 => std_logic_vector(to_unsigned(146,8) ,
12556	 => std_logic_vector(to_unsigned(139,8) ,
12557	 => std_logic_vector(to_unsigned(139,8) ,
12558	 => std_logic_vector(to_unsigned(136,8) ,
12559	 => std_logic_vector(to_unsigned(144,8) ,
12560	 => std_logic_vector(to_unsigned(146,8) ,
12561	 => std_logic_vector(to_unsigned(144,8) ,
12562	 => std_logic_vector(to_unsigned(136,8) ,
12563	 => std_logic_vector(to_unsigned(139,8) ,
12564	 => std_logic_vector(to_unsigned(144,8) ,
12565	 => std_logic_vector(to_unsigned(154,8) ,
12566	 => std_logic_vector(to_unsigned(134,8) ,
12567	 => std_logic_vector(to_unsigned(122,8) ,
12568	 => std_logic_vector(to_unsigned(118,8) ,
12569	 => std_logic_vector(to_unsigned(130,8) ,
12570	 => std_logic_vector(to_unsigned(142,8) ,
12571	 => std_logic_vector(to_unsigned(142,8) ,
12572	 => std_logic_vector(to_unsigned(139,8) ,
12573	 => std_logic_vector(to_unsigned(139,8) ,
12574	 => std_logic_vector(to_unsigned(136,8) ,
12575	 => std_logic_vector(to_unsigned(131,8) ,
12576	 => std_logic_vector(to_unsigned(130,8) ,
12577	 => std_logic_vector(to_unsigned(128,8) ,
12578	 => std_logic_vector(to_unsigned(130,8) ,
12579	 => std_logic_vector(to_unsigned(128,8) ,
12580	 => std_logic_vector(to_unsigned(131,8) ,
12581	 => std_logic_vector(to_unsigned(146,8) ,
12582	 => std_logic_vector(to_unsigned(142,8) ,
12583	 => std_logic_vector(to_unsigned(134,8) ,
12584	 => std_logic_vector(to_unsigned(125,8) ,
12585	 => std_logic_vector(to_unsigned(116,8) ,
12586	 => std_logic_vector(to_unsigned(108,8) ,
12587	 => std_logic_vector(to_unsigned(96,8) ,
12588	 => std_logic_vector(to_unsigned(97,8) ,
12589	 => std_logic_vector(to_unsigned(103,8) ,
12590	 => std_logic_vector(to_unsigned(97,8) ,
12591	 => std_logic_vector(to_unsigned(96,8) ,
12592	 => std_logic_vector(to_unsigned(99,8) ,
12593	 => std_logic_vector(to_unsigned(100,8) ,
12594	 => std_logic_vector(to_unsigned(103,8) ,
12595	 => std_logic_vector(to_unsigned(115,8) ,
12596	 => std_logic_vector(to_unsigned(130,8) ,
12597	 => std_logic_vector(to_unsigned(118,8) ,
12598	 => std_logic_vector(to_unsigned(101,8) ,
12599	 => std_logic_vector(to_unsigned(107,8) ,
12600	 => std_logic_vector(to_unsigned(112,8) ,
12601	 => std_logic_vector(to_unsigned(124,8) ,
12602	 => std_logic_vector(to_unsigned(127,8) ,
12603	 => std_logic_vector(to_unsigned(127,8) ,
12604	 => std_logic_vector(to_unsigned(130,8) ,
12605	 => std_logic_vector(to_unsigned(131,8) ,
12606	 => std_logic_vector(to_unsigned(127,8) ,
12607	 => std_logic_vector(to_unsigned(119,8) ,
12608	 => std_logic_vector(to_unsigned(115,8) ,
12609	 => std_logic_vector(to_unsigned(112,8) ,
12610	 => std_logic_vector(to_unsigned(115,8) ,
12611	 => std_logic_vector(to_unsigned(119,8) ,
12612	 => std_logic_vector(to_unsigned(109,8) ,
12613	 => std_logic_vector(to_unsigned(96,8) ,
12614	 => std_logic_vector(to_unsigned(100,8) ,
12615	 => std_logic_vector(to_unsigned(93,8) ,
12616	 => std_logic_vector(to_unsigned(96,8) ,
12617	 => std_logic_vector(to_unsigned(100,8) ,
12618	 => std_logic_vector(to_unsigned(107,8) ,
12619	 => std_logic_vector(to_unsigned(118,8) ,
12620	 => std_logic_vector(to_unsigned(114,8) ,
12621	 => std_logic_vector(to_unsigned(118,8) ,
12622	 => std_logic_vector(to_unsigned(103,8) ,
12623	 => std_logic_vector(to_unsigned(91,8) ,
12624	 => std_logic_vector(to_unsigned(108,8) ,
12625	 => std_logic_vector(to_unsigned(111,8) ,
12626	 => std_logic_vector(to_unsigned(114,8) ,
12627	 => std_logic_vector(to_unsigned(114,8) ,
12628	 => std_logic_vector(to_unsigned(109,8) ,
12629	 => std_logic_vector(to_unsigned(107,8) ,
12630	 => std_logic_vector(to_unsigned(100,8) ,
12631	 => std_logic_vector(to_unsigned(91,8) ,
12632	 => std_logic_vector(to_unsigned(91,8) ,
12633	 => std_logic_vector(to_unsigned(100,8) ,
12634	 => std_logic_vector(to_unsigned(88,8) ,
12635	 => std_logic_vector(to_unsigned(80,8) ,
12636	 => std_logic_vector(to_unsigned(101,8) ,
12637	 => std_logic_vector(to_unsigned(103,8) ,
12638	 => std_logic_vector(to_unsigned(114,8) ,
12639	 => std_logic_vector(to_unsigned(92,8) ,
12640	 => std_logic_vector(to_unsigned(74,8) ,
12641	 => std_logic_vector(to_unsigned(95,8) ,
12642	 => std_logic_vector(to_unsigned(95,8) ,
12643	 => std_logic_vector(to_unsigned(63,8) ,
12644	 => std_logic_vector(to_unsigned(74,8) ,
12645	 => std_logic_vector(to_unsigned(74,8) ,
12646	 => std_logic_vector(to_unsigned(68,8) ,
12647	 => std_logic_vector(to_unsigned(82,8) ,
12648	 => std_logic_vector(to_unsigned(95,8) ,
12649	 => std_logic_vector(to_unsigned(93,8) ,
12650	 => std_logic_vector(to_unsigned(91,8) ,
12651	 => std_logic_vector(to_unsigned(86,8) ,
12652	 => std_logic_vector(to_unsigned(73,8) ,
12653	 => std_logic_vector(to_unsigned(74,8) ,
12654	 => std_logic_vector(to_unsigned(76,8) ,
12655	 => std_logic_vector(to_unsigned(73,8) ,
12656	 => std_logic_vector(to_unsigned(79,8) ,
12657	 => std_logic_vector(to_unsigned(77,8) ,
12658	 => std_logic_vector(to_unsigned(87,8) ,
12659	 => std_logic_vector(to_unsigned(88,8) ,
12660	 => std_logic_vector(to_unsigned(65,8) ,
12661	 => std_logic_vector(to_unsigned(69,8) ,
12662	 => std_logic_vector(to_unsigned(88,8) ,
12663	 => std_logic_vector(to_unsigned(103,8) ,
12664	 => std_logic_vector(to_unsigned(97,8) ,
12665	 => std_logic_vector(to_unsigned(86,8) ,
12666	 => std_logic_vector(to_unsigned(88,8) ,
12667	 => std_logic_vector(to_unsigned(82,8) ,
12668	 => std_logic_vector(to_unsigned(76,8) ,
12669	 => std_logic_vector(to_unsigned(74,8) ,
12670	 => std_logic_vector(to_unsigned(86,8) ,
12671	 => std_logic_vector(to_unsigned(71,8) ,
12672	 => std_logic_vector(to_unsigned(63,8) ,
12673	 => std_logic_vector(to_unsigned(64,8) ,
12674	 => std_logic_vector(to_unsigned(79,8) ,
12675	 => std_logic_vector(to_unsigned(95,8) ,
12676	 => std_logic_vector(to_unsigned(101,8) ,
12677	 => std_logic_vector(to_unsigned(105,8) ,
12678	 => std_logic_vector(to_unsigned(112,8) ,
12679	 => std_logic_vector(to_unsigned(119,8) ,
12680	 => std_logic_vector(to_unsigned(109,8) ,
12681	 => std_logic_vector(to_unsigned(119,8) ,
12682	 => std_logic_vector(to_unsigned(118,8) ,
12683	 => std_logic_vector(to_unsigned(88,8) ,
12684	 => std_logic_vector(to_unsigned(78,8) ,
12685	 => std_logic_vector(to_unsigned(101,8) ,
12686	 => std_logic_vector(to_unsigned(101,8) ,
12687	 => std_logic_vector(to_unsigned(97,8) ,
12688	 => std_logic_vector(to_unsigned(115,8) ,
12689	 => std_logic_vector(to_unsigned(100,8) ,
12690	 => std_logic_vector(to_unsigned(79,8) ,
12691	 => std_logic_vector(to_unsigned(92,8) ,
12692	 => std_logic_vector(to_unsigned(85,8) ,
12693	 => std_logic_vector(to_unsigned(74,8) ,
12694	 => std_logic_vector(to_unsigned(84,8) ,
12695	 => std_logic_vector(to_unsigned(99,8) ,
12696	 => std_logic_vector(to_unsigned(114,8) ,
12697	 => std_logic_vector(to_unsigned(108,8) ,
12698	 => std_logic_vector(to_unsigned(100,8) ,
12699	 => std_logic_vector(to_unsigned(96,8) ,
12700	 => std_logic_vector(to_unsigned(88,8) ,
12701	 => std_logic_vector(to_unsigned(85,8) ,
12702	 => std_logic_vector(to_unsigned(87,8) ,
12703	 => std_logic_vector(to_unsigned(86,8) ,
12704	 => std_logic_vector(to_unsigned(84,8) ,
12705	 => std_logic_vector(to_unsigned(90,8) ,
12706	 => std_logic_vector(to_unsigned(90,8) ,
12707	 => std_logic_vector(to_unsigned(80,8) ,
12708	 => std_logic_vector(to_unsigned(73,8) ,
12709	 => std_logic_vector(to_unsigned(79,8) ,
12710	 => std_logic_vector(to_unsigned(79,8) ,
12711	 => std_logic_vector(to_unsigned(80,8) ,
12712	 => std_logic_vector(to_unsigned(84,8) ,
12713	 => std_logic_vector(to_unsigned(90,8) ,
12714	 => std_logic_vector(to_unsigned(84,8) ,
12715	 => std_logic_vector(to_unsigned(85,8) ,
12716	 => std_logic_vector(to_unsigned(79,8) ,
12717	 => std_logic_vector(to_unsigned(73,8) ,
12718	 => std_logic_vector(to_unsigned(77,8) ,
12719	 => std_logic_vector(to_unsigned(64,8) ,
12720	 => std_logic_vector(to_unsigned(58,8) ,
12721	 => std_logic_vector(to_unsigned(76,8) ,
12722	 => std_logic_vector(to_unsigned(73,8) ,
12723	 => std_logic_vector(to_unsigned(91,8) ,
12724	 => std_logic_vector(to_unsigned(58,8) ,
12725	 => std_logic_vector(to_unsigned(2,8) ,
12726	 => std_logic_vector(to_unsigned(0,8) ,
12727	 => std_logic_vector(to_unsigned(1,8) ,
12728	 => std_logic_vector(to_unsigned(27,8) ,
12729	 => std_logic_vector(to_unsigned(51,8) ,
12730	 => std_logic_vector(to_unsigned(44,8) ,
12731	 => std_logic_vector(to_unsigned(48,8) ,
12732	 => std_logic_vector(to_unsigned(48,8) ,
12733	 => std_logic_vector(to_unsigned(37,8) ,
12734	 => std_logic_vector(to_unsigned(43,8) ,
12735	 => std_logic_vector(to_unsigned(60,8) ,
12736	 => std_logic_vector(to_unsigned(61,8) ,
12737	 => std_logic_vector(to_unsigned(42,8) ,
12738	 => std_logic_vector(to_unsigned(44,8) ,
12739	 => std_logic_vector(to_unsigned(44,8) ,
12740	 => std_logic_vector(to_unsigned(44,8) ,
12741	 => std_logic_vector(to_unsigned(46,8) ,
12742	 => std_logic_vector(to_unsigned(49,8) ,
12743	 => std_logic_vector(to_unsigned(49,8) ,
12744	 => std_logic_vector(to_unsigned(53,8) ,
12745	 => std_logic_vector(to_unsigned(58,8) ,
12746	 => std_logic_vector(to_unsigned(55,8) ,
12747	 => std_logic_vector(to_unsigned(54,8) ,
12748	 => std_logic_vector(to_unsigned(56,8) ,
12749	 => std_logic_vector(to_unsigned(57,8) ,
12750	 => std_logic_vector(to_unsigned(54,8) ,
12751	 => std_logic_vector(to_unsigned(59,8) ,
12752	 => std_logic_vector(to_unsigned(59,8) ,
12753	 => std_logic_vector(to_unsigned(62,8) ,
12754	 => std_logic_vector(to_unsigned(61,8) ,
12755	 => std_logic_vector(to_unsigned(61,8) ,
12756	 => std_logic_vector(to_unsigned(67,8) ,
12757	 => std_logic_vector(to_unsigned(77,8) ,
12758	 => std_logic_vector(to_unsigned(68,8) ,
12759	 => std_logic_vector(to_unsigned(68,8) ,
12760	 => std_logic_vector(to_unsigned(79,8) ,
12761	 => std_logic_vector(to_unsigned(79,8) ,
12762	 => std_logic_vector(to_unsigned(82,8) ,
12763	 => std_logic_vector(to_unsigned(70,8) ,
12764	 => std_logic_vector(to_unsigned(82,8) ,
12765	 => std_logic_vector(to_unsigned(95,8) ,
12766	 => std_logic_vector(to_unsigned(78,8) ,
12767	 => std_logic_vector(to_unsigned(77,8) ,
12768	 => std_logic_vector(to_unsigned(88,8) ,
12769	 => std_logic_vector(to_unsigned(84,8) ,
12770	 => std_logic_vector(to_unsigned(81,8) ,
12771	 => std_logic_vector(to_unsigned(85,8) ,
12772	 => std_logic_vector(to_unsigned(86,8) ,
12773	 => std_logic_vector(to_unsigned(88,8) ,
12774	 => std_logic_vector(to_unsigned(95,8) ,
12775	 => std_logic_vector(to_unsigned(103,8) ,
12776	 => std_logic_vector(to_unsigned(111,8) ,
12777	 => std_logic_vector(to_unsigned(114,8) ,
12778	 => std_logic_vector(to_unsigned(115,8) ,
12779	 => std_logic_vector(to_unsigned(124,8) ,
12780	 => std_logic_vector(to_unsigned(130,8) ,
12781	 => std_logic_vector(to_unsigned(128,8) ,
12782	 => std_logic_vector(to_unsigned(139,8) ,
12783	 => std_logic_vector(to_unsigned(142,8) ,
12784	 => std_logic_vector(to_unsigned(136,8) ,
12785	 => std_logic_vector(to_unsigned(147,8) ,
12786	 => std_logic_vector(to_unsigned(144,8) ,
12787	 => std_logic_vector(to_unsigned(147,8) ,
12788	 => std_logic_vector(to_unsigned(151,8) ,
12789	 => std_logic_vector(to_unsigned(149,8) ,
12790	 => std_logic_vector(to_unsigned(149,8) ,
12791	 => std_logic_vector(to_unsigned(147,8) ,
12792	 => std_logic_vector(to_unsigned(141,8) ,
12793	 => std_logic_vector(to_unsigned(130,8) ,
12794	 => std_logic_vector(to_unsigned(130,8) ,
12795	 => std_logic_vector(to_unsigned(138,8) ,
12796	 => std_logic_vector(to_unsigned(146,8) ,
12797	 => std_logic_vector(to_unsigned(136,8) ,
12798	 => std_logic_vector(to_unsigned(142,8) ,
12799	 => std_logic_vector(to_unsigned(149,8) ,
12800	 => std_logic_vector(to_unsigned(151,8) ,
12801	 => std_logic_vector(to_unsigned(142,8) ,
12802	 => std_logic_vector(to_unsigned(144,8) ,
12803	 => std_logic_vector(to_unsigned(146,8) ,
12804	 => std_logic_vector(to_unsigned(146,8) ,
12805	 => std_logic_vector(to_unsigned(144,8) ,
12806	 => std_logic_vector(to_unsigned(146,8) ,
12807	 => std_logic_vector(to_unsigned(147,8) ,
12808	 => std_logic_vector(to_unsigned(151,8) ,
12809	 => std_logic_vector(to_unsigned(142,8) ,
12810	 => std_logic_vector(to_unsigned(141,8) ,
12811	 => std_logic_vector(to_unsigned(147,8) ,
12812	 => std_logic_vector(to_unsigned(151,8) ,
12813	 => std_logic_vector(to_unsigned(156,8) ,
12814	 => std_logic_vector(to_unsigned(154,8) ,
12815	 => std_logic_vector(to_unsigned(156,8) ,
12816	 => std_logic_vector(to_unsigned(152,8) ,
12817	 => std_logic_vector(to_unsigned(152,8) ,
12818	 => std_logic_vector(to_unsigned(151,8) ,
12819	 => std_logic_vector(to_unsigned(156,8) ,
12820	 => std_logic_vector(to_unsigned(156,8) ,
12821	 => std_logic_vector(to_unsigned(154,8) ,
12822	 => std_logic_vector(to_unsigned(157,8) ,
12823	 => std_logic_vector(to_unsigned(159,8) ,
12824	 => std_logic_vector(to_unsigned(157,8) ,
12825	 => std_logic_vector(to_unsigned(156,8) ,
12826	 => std_logic_vector(to_unsigned(156,8) ,
12827	 => std_logic_vector(to_unsigned(159,8) ,
12828	 => std_logic_vector(to_unsigned(152,8) ,
12829	 => std_logic_vector(to_unsigned(125,8) ,
12830	 => std_logic_vector(to_unsigned(114,8) ,
12831	 => std_logic_vector(to_unsigned(116,8) ,
12832	 => std_logic_vector(to_unsigned(114,8) ,
12833	 => std_logic_vector(to_unsigned(114,8) ,
12834	 => std_logic_vector(to_unsigned(119,8) ,
12835	 => std_logic_vector(to_unsigned(116,8) ,
12836	 => std_logic_vector(to_unsigned(108,8) ,
12837	 => std_logic_vector(to_unsigned(108,8) ,
12838	 => std_logic_vector(to_unsigned(109,8) ,
12839	 => std_logic_vector(to_unsigned(136,8) ,
12840	 => std_logic_vector(to_unsigned(147,8) ,
12841	 => std_logic_vector(to_unsigned(139,8) ,
12842	 => std_logic_vector(to_unsigned(138,8) ,
12843	 => std_logic_vector(to_unsigned(119,8) ,
12844	 => std_logic_vector(to_unsigned(122,8) ,
12845	 => std_logic_vector(to_unsigned(133,8) ,
12846	 => std_logic_vector(to_unsigned(124,8) ,
12847	 => std_logic_vector(to_unsigned(116,8) ,
12848	 => std_logic_vector(to_unsigned(115,8) ,
12849	 => std_logic_vector(to_unsigned(130,8) ,
12850	 => std_logic_vector(to_unsigned(134,8) ,
12851	 => std_logic_vector(to_unsigned(128,8) ,
12852	 => std_logic_vector(to_unsigned(109,8) ,
12853	 => std_logic_vector(to_unsigned(104,8) ,
12854	 => std_logic_vector(to_unsigned(109,8) ,
12855	 => std_logic_vector(to_unsigned(136,8) ,
12856	 => std_logic_vector(to_unsigned(142,8) ,
12857	 => std_logic_vector(to_unsigned(136,8) ,
12858	 => std_logic_vector(to_unsigned(133,8) ,
12859	 => std_logic_vector(to_unsigned(141,8) ,
12860	 => std_logic_vector(to_unsigned(149,8) ,
12861	 => std_logic_vector(to_unsigned(141,8) ,
12862	 => std_logic_vector(to_unsigned(136,8) ,
12863	 => std_logic_vector(to_unsigned(141,8) ,
12864	 => std_logic_vector(to_unsigned(138,8) ,
12865	 => std_logic_vector(to_unsigned(134,8) ,
12866	 => std_logic_vector(to_unsigned(136,8) ,
12867	 => std_logic_vector(to_unsigned(142,8) ,
12868	 => std_logic_vector(to_unsigned(133,8) ,
12869	 => std_logic_vector(to_unsigned(112,8) ,
12870	 => std_logic_vector(to_unsigned(125,8) ,
12871	 => std_logic_vector(to_unsigned(136,8) ,
12872	 => std_logic_vector(to_unsigned(149,8) ,
12873	 => std_logic_vector(to_unsigned(139,8) ,
12874	 => std_logic_vector(to_unsigned(130,8) ,
12875	 => std_logic_vector(to_unsigned(128,8) ,
12876	 => std_logic_vector(to_unsigned(134,8) ,
12877	 => std_logic_vector(to_unsigned(136,8) ,
12878	 => std_logic_vector(to_unsigned(139,8) ,
12879	 => std_logic_vector(to_unsigned(139,8) ,
12880	 => std_logic_vector(to_unsigned(136,8) ,
12881	 => std_logic_vector(to_unsigned(131,8) ,
12882	 => std_logic_vector(to_unsigned(136,8) ,
12883	 => std_logic_vector(to_unsigned(146,8) ,
12884	 => std_logic_vector(to_unsigned(144,8) ,
12885	 => std_logic_vector(to_unsigned(152,8) ,
12886	 => std_logic_vector(to_unsigned(142,8) ,
12887	 => std_logic_vector(to_unsigned(127,8) ,
12888	 => std_logic_vector(to_unsigned(144,8) ,
12889	 => std_logic_vector(to_unsigned(147,8) ,
12890	 => std_logic_vector(to_unsigned(154,8) ,
12891	 => std_logic_vector(to_unsigned(151,8) ,
12892	 => std_logic_vector(to_unsigned(139,8) ,
12893	 => std_logic_vector(to_unsigned(141,8) ,
12894	 => std_logic_vector(to_unsigned(139,8) ,
12895	 => std_logic_vector(to_unsigned(134,8) ,
12896	 => std_logic_vector(to_unsigned(136,8) ,
12897	 => std_logic_vector(to_unsigned(141,8) ,
12898	 => std_logic_vector(to_unsigned(138,8) ,
12899	 => std_logic_vector(to_unsigned(133,8) ,
12900	 => std_logic_vector(to_unsigned(138,8) ,
12901	 => std_logic_vector(to_unsigned(149,8) ,
12902	 => std_logic_vector(to_unsigned(152,8) ,
12903	 => std_logic_vector(to_unsigned(139,8) ,
12904	 => std_logic_vector(to_unsigned(124,8) ,
12905	 => std_logic_vector(to_unsigned(115,8) ,
12906	 => std_logic_vector(to_unsigned(108,8) ,
12907	 => std_logic_vector(to_unsigned(100,8) ,
12908	 => std_logic_vector(to_unsigned(107,8) ,
12909	 => std_logic_vector(to_unsigned(127,8) ,
12910	 => std_logic_vector(to_unsigned(116,8) ,
12911	 => std_logic_vector(to_unsigned(103,8) ,
12912	 => std_logic_vector(to_unsigned(111,8) ,
12913	 => std_logic_vector(to_unsigned(119,8) ,
12914	 => std_logic_vector(to_unsigned(121,8) ,
12915	 => std_logic_vector(to_unsigned(114,8) ,
12916	 => std_logic_vector(to_unsigned(116,8) ,
12917	 => std_logic_vector(to_unsigned(119,8) ,
12918	 => std_logic_vector(to_unsigned(114,8) ,
12919	 => std_logic_vector(to_unsigned(115,8) ,
12920	 => std_logic_vector(to_unsigned(124,8) ,
12921	 => std_logic_vector(to_unsigned(127,8) ,
12922	 => std_logic_vector(to_unsigned(127,8) ,
12923	 => std_logic_vector(to_unsigned(130,8) ,
12924	 => std_logic_vector(to_unsigned(141,8) ,
12925	 => std_logic_vector(to_unsigned(149,8) ,
12926	 => std_logic_vector(to_unsigned(125,8) ,
12927	 => std_logic_vector(to_unsigned(112,8) ,
12928	 => std_logic_vector(to_unsigned(116,8) ,
12929	 => std_logic_vector(to_unsigned(108,8) ,
12930	 => std_logic_vector(to_unsigned(114,8) ,
12931	 => std_logic_vector(to_unsigned(115,8) ,
12932	 => std_logic_vector(to_unsigned(100,8) ,
12933	 => std_logic_vector(to_unsigned(90,8) ,
12934	 => std_logic_vector(to_unsigned(96,8) ,
12935	 => std_logic_vector(to_unsigned(96,8) ,
12936	 => std_logic_vector(to_unsigned(100,8) ,
12937	 => std_logic_vector(to_unsigned(95,8) ,
12938	 => std_logic_vector(to_unsigned(115,8) ,
12939	 => std_logic_vector(to_unsigned(128,8) ,
12940	 => std_logic_vector(to_unsigned(115,8) ,
12941	 => std_logic_vector(to_unsigned(118,8) ,
12942	 => std_logic_vector(to_unsigned(99,8) ,
12943	 => std_logic_vector(to_unsigned(90,8) ,
12944	 => std_logic_vector(to_unsigned(107,8) ,
12945	 => std_logic_vector(to_unsigned(112,8) ,
12946	 => std_logic_vector(to_unsigned(114,8) ,
12947	 => std_logic_vector(to_unsigned(115,8) ,
12948	 => std_logic_vector(to_unsigned(109,8) ,
12949	 => std_logic_vector(to_unsigned(111,8) ,
12950	 => std_logic_vector(to_unsigned(111,8) ,
12951	 => std_logic_vector(to_unsigned(104,8) ,
12952	 => std_logic_vector(to_unsigned(90,8) ,
12953	 => std_logic_vector(to_unsigned(84,8) ,
12954	 => std_logic_vector(to_unsigned(85,8) ,
12955	 => std_logic_vector(to_unsigned(72,8) ,
12956	 => std_logic_vector(to_unsigned(92,8) ,
12957	 => std_logic_vector(to_unsigned(103,8) ,
12958	 => std_logic_vector(to_unsigned(108,8) ,
12959	 => std_logic_vector(to_unsigned(87,8) ,
12960	 => std_logic_vector(to_unsigned(73,8) ,
12961	 => std_logic_vector(to_unsigned(99,8) ,
12962	 => std_logic_vector(to_unsigned(96,8) ,
12963	 => std_logic_vector(to_unsigned(70,8) ,
12964	 => std_logic_vector(to_unsigned(86,8) ,
12965	 => std_logic_vector(to_unsigned(88,8) ,
12966	 => std_logic_vector(to_unsigned(87,8) ,
12967	 => std_logic_vector(to_unsigned(95,8) ,
12968	 => std_logic_vector(to_unsigned(101,8) ,
12969	 => std_logic_vector(to_unsigned(97,8) ,
12970	 => std_logic_vector(to_unsigned(84,8) ,
12971	 => std_logic_vector(to_unsigned(90,8) ,
12972	 => std_logic_vector(to_unsigned(104,8) ,
12973	 => std_logic_vector(to_unsigned(93,8) ,
12974	 => std_logic_vector(to_unsigned(79,8) ,
12975	 => std_logic_vector(to_unsigned(74,8) ,
12976	 => std_logic_vector(to_unsigned(78,8) ,
12977	 => std_logic_vector(to_unsigned(84,8) ,
12978	 => std_logic_vector(to_unsigned(86,8) ,
12979	 => std_logic_vector(to_unsigned(84,8) ,
12980	 => std_logic_vector(to_unsigned(67,8) ,
12981	 => std_logic_vector(to_unsigned(69,8) ,
12982	 => std_logic_vector(to_unsigned(93,8) ,
12983	 => std_logic_vector(to_unsigned(112,8) ,
12984	 => std_logic_vector(to_unsigned(114,8) ,
12985	 => std_logic_vector(to_unsigned(105,8) ,
12986	 => std_logic_vector(to_unsigned(108,8) ,
12987	 => std_logic_vector(to_unsigned(100,8) ,
12988	 => std_logic_vector(to_unsigned(90,8) ,
12989	 => std_logic_vector(to_unsigned(91,8) ,
12990	 => std_logic_vector(to_unsigned(104,8) ,
12991	 => std_logic_vector(to_unsigned(86,8) ,
12992	 => std_logic_vector(to_unsigned(74,8) ,
12993	 => std_logic_vector(to_unsigned(90,8) ,
12994	 => std_logic_vector(to_unsigned(84,8) ,
12995	 => std_logic_vector(to_unsigned(92,8) ,
12996	 => std_logic_vector(to_unsigned(97,8) ,
12997	 => std_logic_vector(to_unsigned(86,8) ,
12998	 => std_logic_vector(to_unsigned(97,8) ,
12999	 => std_logic_vector(to_unsigned(118,8) ,
13000	 => std_logic_vector(to_unsigned(114,8) ,
13001	 => std_logic_vector(to_unsigned(112,8) ,
13002	 => std_logic_vector(to_unsigned(112,8) ,
13003	 => std_logic_vector(to_unsigned(101,8) ,
13004	 => std_logic_vector(to_unsigned(92,8) ,
13005	 => std_logic_vector(to_unsigned(109,8) ,
13006	 => std_logic_vector(to_unsigned(101,8) ,
13007	 => std_logic_vector(to_unsigned(90,8) ,
13008	 => std_logic_vector(to_unsigned(105,8) ,
13009	 => std_logic_vector(to_unsigned(93,8) ,
13010	 => std_logic_vector(to_unsigned(93,8) ,
13011	 => std_logic_vector(to_unsigned(108,8) ,
13012	 => std_logic_vector(to_unsigned(99,8) ,
13013	 => std_logic_vector(to_unsigned(87,8) ,
13014	 => std_logic_vector(to_unsigned(91,8) ,
13015	 => std_logic_vector(to_unsigned(86,8) ,
13016	 => std_logic_vector(to_unsigned(97,8) ,
13017	 => std_logic_vector(to_unsigned(104,8) ,
13018	 => std_logic_vector(to_unsigned(101,8) ,
13019	 => std_logic_vector(to_unsigned(118,8) ,
13020	 => std_logic_vector(to_unsigned(114,8) ,
13021	 => std_logic_vector(to_unsigned(108,8) ,
13022	 => std_logic_vector(to_unsigned(100,8) ,
13023	 => std_logic_vector(to_unsigned(99,8) ,
13024	 => std_logic_vector(to_unsigned(97,8) ,
13025	 => std_logic_vector(to_unsigned(86,8) ,
13026	 => std_logic_vector(to_unsigned(93,8) ,
13027	 => std_logic_vector(to_unsigned(87,8) ,
13028	 => std_logic_vector(to_unsigned(79,8) ,
13029	 => std_logic_vector(to_unsigned(81,8) ,
13030	 => std_logic_vector(to_unsigned(84,8) ,
13031	 => std_logic_vector(to_unsigned(87,8) ,
13032	 => std_logic_vector(to_unsigned(87,8) ,
13033	 => std_logic_vector(to_unsigned(96,8) ,
13034	 => std_logic_vector(to_unsigned(92,8) ,
13035	 => std_logic_vector(to_unsigned(85,8) ,
13036	 => std_logic_vector(to_unsigned(79,8) ,
13037	 => std_logic_vector(to_unsigned(73,8) ,
13038	 => std_logic_vector(to_unsigned(76,8) ,
13039	 => std_logic_vector(to_unsigned(66,8) ,
13040	 => std_logic_vector(to_unsigned(72,8) ,
13041	 => std_logic_vector(to_unsigned(84,8) ,
13042	 => std_logic_vector(to_unsigned(80,8) ,
13043	 => std_logic_vector(to_unsigned(90,8) ,
13044	 => std_logic_vector(to_unsigned(45,8) ,
13045	 => std_logic_vector(to_unsigned(3,8) ,
13046	 => std_logic_vector(to_unsigned(0,8) ,
13047	 => std_logic_vector(to_unsigned(0,8) ,
13048	 => std_logic_vector(to_unsigned(16,8) ,
13049	 => std_logic_vector(to_unsigned(61,8) ,
13050	 => std_logic_vector(to_unsigned(47,8) ,
13051	 => std_logic_vector(to_unsigned(51,8) ,
13052	 => std_logic_vector(to_unsigned(47,8) ,
13053	 => std_logic_vector(to_unsigned(42,8) ,
13054	 => std_logic_vector(to_unsigned(41,8) ,
13055	 => std_logic_vector(to_unsigned(64,8) ,
13056	 => std_logic_vector(to_unsigned(67,8) ,
13057	 => std_logic_vector(to_unsigned(46,8) ,
13058	 => std_logic_vector(to_unsigned(41,8) ,
13059	 => std_logic_vector(to_unsigned(53,8) ,
13060	 => std_logic_vector(to_unsigned(54,8) ,
13061	 => std_logic_vector(to_unsigned(51,8) ,
13062	 => std_logic_vector(to_unsigned(51,8) ,
13063	 => std_logic_vector(to_unsigned(57,8) ,
13064	 => std_logic_vector(to_unsigned(82,8) ,
13065	 => std_logic_vector(to_unsigned(85,8) ,
13066	 => std_logic_vector(to_unsigned(64,8) ,
13067	 => std_logic_vector(to_unsigned(56,8) ,
13068	 => std_logic_vector(to_unsigned(56,8) ,
13069	 => std_logic_vector(to_unsigned(60,8) ,
13070	 => std_logic_vector(to_unsigned(62,8) ,
13071	 => std_logic_vector(to_unsigned(68,8) ,
13072	 => std_logic_vector(to_unsigned(71,8) ,
13073	 => std_logic_vector(to_unsigned(61,8) ,
13074	 => std_logic_vector(to_unsigned(56,8) ,
13075	 => std_logic_vector(to_unsigned(52,8) ,
13076	 => std_logic_vector(to_unsigned(56,8) ,
13077	 => std_logic_vector(to_unsigned(57,8) ,
13078	 => std_logic_vector(to_unsigned(56,8) ,
13079	 => std_logic_vector(to_unsigned(61,8) ,
13080	 => std_logic_vector(to_unsigned(67,8) ,
13081	 => std_logic_vector(to_unsigned(77,8) ,
13082	 => std_logic_vector(to_unsigned(78,8) ,
13083	 => std_logic_vector(to_unsigned(66,8) ,
13084	 => std_logic_vector(to_unsigned(79,8) ,
13085	 => std_logic_vector(to_unsigned(101,8) ,
13086	 => std_logic_vector(to_unsigned(90,8) ,
13087	 => std_logic_vector(to_unsigned(81,8) ,
13088	 => std_logic_vector(to_unsigned(96,8) ,
13089	 => std_logic_vector(to_unsigned(100,8) ,
13090	 => std_logic_vector(to_unsigned(90,8) ,
13091	 => std_logic_vector(to_unsigned(84,8) ,
13092	 => std_logic_vector(to_unsigned(90,8) ,
13093	 => std_logic_vector(to_unsigned(97,8) ,
13094	 => std_logic_vector(to_unsigned(108,8) ,
13095	 => std_logic_vector(to_unsigned(116,8) ,
13096	 => std_logic_vector(to_unsigned(124,8) ,
13097	 => std_logic_vector(to_unsigned(128,8) ,
13098	 => std_logic_vector(to_unsigned(128,8) ,
13099	 => std_logic_vector(to_unsigned(146,8) ,
13100	 => std_logic_vector(to_unsigned(159,8) ,
13101	 => std_logic_vector(to_unsigned(161,8) ,
13102	 => std_logic_vector(to_unsigned(161,8) ,
13103	 => std_logic_vector(to_unsigned(157,8) ,
13104	 => std_logic_vector(to_unsigned(161,8) ,
13105	 => std_logic_vector(to_unsigned(163,8) ,
13106	 => std_logic_vector(to_unsigned(161,8) ,
13107	 => std_logic_vector(to_unsigned(161,8) ,
13108	 => std_logic_vector(to_unsigned(156,8) ,
13109	 => std_logic_vector(to_unsigned(161,8) ,
13110	 => std_logic_vector(to_unsigned(161,8) ,
13111	 => std_logic_vector(to_unsigned(157,8) ,
13112	 => std_logic_vector(to_unsigned(159,8) ,
13113	 => std_logic_vector(to_unsigned(152,8) ,
13114	 => std_logic_vector(to_unsigned(144,8) ,
13115	 => std_logic_vector(to_unsigned(141,8) ,
13116	 => std_logic_vector(to_unsigned(139,8) ,
13117	 => std_logic_vector(to_unsigned(131,8) ,
13118	 => std_logic_vector(to_unsigned(134,8) ,
13119	 => std_logic_vector(to_unsigned(149,8) ,
13120	 => std_logic_vector(to_unsigned(156,8) ,
13121	 => std_logic_vector(to_unsigned(151,8) ,
13122	 => std_logic_vector(to_unsigned(151,8) ,
13123	 => std_logic_vector(to_unsigned(147,8) ,
13124	 => std_logic_vector(to_unsigned(152,8) ,
13125	 => std_logic_vector(to_unsigned(151,8) ,
13126	 => std_logic_vector(to_unsigned(147,8) ,
13127	 => std_logic_vector(to_unsigned(131,8) ,
13128	 => std_logic_vector(to_unsigned(130,8) ,
13129	 => std_logic_vector(to_unsigned(149,8) ,
13130	 => std_logic_vector(to_unsigned(149,8) ,
13131	 => std_logic_vector(to_unsigned(149,8) ,
13132	 => std_logic_vector(to_unsigned(154,8) ,
13133	 => std_logic_vector(to_unsigned(157,8) ,
13134	 => std_logic_vector(to_unsigned(157,8) ,
13135	 => std_logic_vector(to_unsigned(154,8) ,
13136	 => std_logic_vector(to_unsigned(154,8) ,
13137	 => std_logic_vector(to_unsigned(159,8) ,
13138	 => std_logic_vector(to_unsigned(157,8) ,
13139	 => std_logic_vector(to_unsigned(152,8) ,
13140	 => std_logic_vector(to_unsigned(159,8) ,
13141	 => std_logic_vector(to_unsigned(157,8) ,
13142	 => std_logic_vector(to_unsigned(156,8) ,
13143	 => std_logic_vector(to_unsigned(163,8) ,
13144	 => std_logic_vector(to_unsigned(159,8) ,
13145	 => std_logic_vector(to_unsigned(159,8) ,
13146	 => std_logic_vector(to_unsigned(159,8) ,
13147	 => std_logic_vector(to_unsigned(156,8) ,
13148	 => std_logic_vector(to_unsigned(152,8) ,
13149	 => std_logic_vector(to_unsigned(124,8) ,
13150	 => std_logic_vector(to_unsigned(112,8) ,
13151	 => std_logic_vector(to_unsigned(118,8) ,
13152	 => std_logic_vector(to_unsigned(116,8) ,
13153	 => std_logic_vector(to_unsigned(111,8) ,
13154	 => std_logic_vector(to_unsigned(119,8) ,
13155	 => std_logic_vector(to_unsigned(111,8) ,
13156	 => std_logic_vector(to_unsigned(107,8) ,
13157	 => std_logic_vector(to_unsigned(108,8) ,
13158	 => std_logic_vector(to_unsigned(108,8) ,
13159	 => std_logic_vector(to_unsigned(124,8) ,
13160	 => std_logic_vector(to_unsigned(141,8) ,
13161	 => std_logic_vector(to_unsigned(144,8) ,
13162	 => std_logic_vector(to_unsigned(144,8) ,
13163	 => std_logic_vector(to_unsigned(130,8) ,
13164	 => std_logic_vector(to_unsigned(127,8) ,
13165	 => std_logic_vector(to_unsigned(136,8) ,
13166	 => std_logic_vector(to_unsigned(128,8) ,
13167	 => std_logic_vector(to_unsigned(125,8) ,
13168	 => std_logic_vector(to_unsigned(133,8) ,
13169	 => std_logic_vector(to_unsigned(136,8) ,
13170	 => std_logic_vector(to_unsigned(136,8) ,
13171	 => std_logic_vector(to_unsigned(136,8) ,
13172	 => std_logic_vector(to_unsigned(122,8) ,
13173	 => std_logic_vector(to_unsigned(130,8) ,
13174	 => std_logic_vector(to_unsigned(138,8) ,
13175	 => std_logic_vector(to_unsigned(147,8) ,
13176	 => std_logic_vector(to_unsigned(151,8) ,
13177	 => std_logic_vector(to_unsigned(149,8) ,
13178	 => std_logic_vector(to_unsigned(151,8) ,
13179	 => std_logic_vector(to_unsigned(151,8) ,
13180	 => std_logic_vector(to_unsigned(149,8) ,
13181	 => std_logic_vector(to_unsigned(151,8) ,
13182	 => std_logic_vector(to_unsigned(154,8) ,
13183	 => std_logic_vector(to_unsigned(141,8) ,
13184	 => std_logic_vector(to_unsigned(128,8) ,
13185	 => std_logic_vector(to_unsigned(134,8) ,
13186	 => std_logic_vector(to_unsigned(134,8) ,
13187	 => std_logic_vector(to_unsigned(128,8) ,
13188	 => std_logic_vector(to_unsigned(127,8) ,
13189	 => std_logic_vector(to_unsigned(114,8) ,
13190	 => std_logic_vector(to_unsigned(116,8) ,
13191	 => std_logic_vector(to_unsigned(119,8) ,
13192	 => std_logic_vector(to_unsigned(125,8) ,
13193	 => std_logic_vector(to_unsigned(125,8) ,
13194	 => std_logic_vector(to_unsigned(124,8) ,
13195	 => std_logic_vector(to_unsigned(116,8) ,
13196	 => std_logic_vector(to_unsigned(108,8) ,
13197	 => std_logic_vector(to_unsigned(111,8) ,
13198	 => std_logic_vector(to_unsigned(112,8) ,
13199	 => std_logic_vector(to_unsigned(111,8) ,
13200	 => std_logic_vector(to_unsigned(121,8) ,
13201	 => std_logic_vector(to_unsigned(131,8) ,
13202	 => std_logic_vector(to_unsigned(144,8) ,
13203	 => std_logic_vector(to_unsigned(146,8) ,
13204	 => std_logic_vector(to_unsigned(144,8) ,
13205	 => std_logic_vector(to_unsigned(151,8) ,
13206	 => std_logic_vector(to_unsigned(151,8) ,
13207	 => std_logic_vector(to_unsigned(124,8) ,
13208	 => std_logic_vector(to_unsigned(146,8) ,
13209	 => std_logic_vector(to_unsigned(136,8) ,
13210	 => std_logic_vector(to_unsigned(149,8) ,
13211	 => std_logic_vector(to_unsigned(159,8) ,
13212	 => std_logic_vector(to_unsigned(149,8) ,
13213	 => std_logic_vector(to_unsigned(146,8) ,
13214	 => std_logic_vector(to_unsigned(133,8) ,
13215	 => std_logic_vector(to_unsigned(134,8) ,
13216	 => std_logic_vector(to_unsigned(147,8) ,
13217	 => std_logic_vector(to_unsigned(144,8) ,
13218	 => std_logic_vector(to_unsigned(134,8) ,
13219	 => std_logic_vector(to_unsigned(133,8) ,
13220	 => std_logic_vector(to_unsigned(138,8) ,
13221	 => std_logic_vector(to_unsigned(144,8) ,
13222	 => std_logic_vector(to_unsigned(142,8) ,
13223	 => std_logic_vector(to_unsigned(142,8) ,
13224	 => std_logic_vector(to_unsigned(127,8) ,
13225	 => std_logic_vector(to_unsigned(115,8) ,
13226	 => std_logic_vector(to_unsigned(121,8) ,
13227	 => std_logic_vector(to_unsigned(111,8) ,
13228	 => std_logic_vector(to_unsigned(122,8) ,
13229	 => std_logic_vector(to_unsigned(138,8) ,
13230	 => std_logic_vector(to_unsigned(121,8) ,
13231	 => std_logic_vector(to_unsigned(101,8) ,
13232	 => std_logic_vector(to_unsigned(93,8) ,
13233	 => std_logic_vector(to_unsigned(104,8) ,
13234	 => std_logic_vector(to_unsigned(114,8) ,
13235	 => std_logic_vector(to_unsigned(107,8) ,
13236	 => std_logic_vector(to_unsigned(107,8) ,
13237	 => std_logic_vector(to_unsigned(114,8) ,
13238	 => std_logic_vector(to_unsigned(131,8) ,
13239	 => std_logic_vector(to_unsigned(131,8) ,
13240	 => std_logic_vector(to_unsigned(122,8) ,
13241	 => std_logic_vector(to_unsigned(121,8) ,
13242	 => std_logic_vector(to_unsigned(119,8) ,
13243	 => std_logic_vector(to_unsigned(128,8) ,
13244	 => std_logic_vector(to_unsigned(142,8) ,
13245	 => std_logic_vector(to_unsigned(147,8) ,
13246	 => std_logic_vector(to_unsigned(124,8) ,
13247	 => std_logic_vector(to_unsigned(112,8) ,
13248	 => std_logic_vector(to_unsigned(127,8) ,
13249	 => std_logic_vector(to_unsigned(122,8) ,
13250	 => std_logic_vector(to_unsigned(125,8) ,
13251	 => std_logic_vector(to_unsigned(122,8) ,
13252	 => std_logic_vector(to_unsigned(105,8) ,
13253	 => std_logic_vector(to_unsigned(103,8) ,
13254	 => std_logic_vector(to_unsigned(95,8) ,
13255	 => std_logic_vector(to_unsigned(103,8) ,
13256	 => std_logic_vector(to_unsigned(100,8) ,
13257	 => std_logic_vector(to_unsigned(99,8) ,
13258	 => std_logic_vector(to_unsigned(115,8) ,
13259	 => std_logic_vector(to_unsigned(124,8) ,
13260	 => std_logic_vector(to_unsigned(125,8) ,
13261	 => std_logic_vector(to_unsigned(118,8) ,
13262	 => std_logic_vector(to_unsigned(96,8) ,
13263	 => std_logic_vector(to_unsigned(90,8) ,
13264	 => std_logic_vector(to_unsigned(116,8) ,
13265	 => std_logic_vector(to_unsigned(111,8) ,
13266	 => std_logic_vector(to_unsigned(107,8) ,
13267	 => std_logic_vector(to_unsigned(119,8) ,
13268	 => std_logic_vector(to_unsigned(115,8) ,
13269	 => std_logic_vector(to_unsigned(115,8) ,
13270	 => std_logic_vector(to_unsigned(116,8) ,
13271	 => std_logic_vector(to_unsigned(112,8) ,
13272	 => std_logic_vector(to_unsigned(90,8) ,
13273	 => std_logic_vector(to_unsigned(77,8) ,
13274	 => std_logic_vector(to_unsigned(79,8) ,
13275	 => std_logic_vector(to_unsigned(74,8) ,
13276	 => std_logic_vector(to_unsigned(103,8) ,
13277	 => std_logic_vector(to_unsigned(104,8) ,
13278	 => std_logic_vector(to_unsigned(103,8) ,
13279	 => std_logic_vector(to_unsigned(88,8) ,
13280	 => std_logic_vector(to_unsigned(80,8) ,
13281	 => std_logic_vector(to_unsigned(100,8) ,
13282	 => std_logic_vector(to_unsigned(97,8) ,
13283	 => std_logic_vector(to_unsigned(84,8) ,
13284	 => std_logic_vector(to_unsigned(99,8) ,
13285	 => std_logic_vector(to_unsigned(92,8) ,
13286	 => std_logic_vector(to_unsigned(86,8) ,
13287	 => std_logic_vector(to_unsigned(91,8) ,
13288	 => std_logic_vector(to_unsigned(80,8) ,
13289	 => std_logic_vector(to_unsigned(76,8) ,
13290	 => std_logic_vector(to_unsigned(70,8) ,
13291	 => std_logic_vector(to_unsigned(87,8) ,
13292	 => std_logic_vector(to_unsigned(125,8) ,
13293	 => std_logic_vector(to_unsigned(105,8) ,
13294	 => std_logic_vector(to_unsigned(86,8) ,
13295	 => std_logic_vector(to_unsigned(85,8) ,
13296	 => std_logic_vector(to_unsigned(87,8) ,
13297	 => std_logic_vector(to_unsigned(88,8) ,
13298	 => std_logic_vector(to_unsigned(86,8) ,
13299	 => std_logic_vector(to_unsigned(85,8) ,
13300	 => std_logic_vector(to_unsigned(73,8) ,
13301	 => std_logic_vector(to_unsigned(77,8) ,
13302	 => std_logic_vector(to_unsigned(97,8) ,
13303	 => std_logic_vector(to_unsigned(112,8) ,
13304	 => std_logic_vector(to_unsigned(108,8) ,
13305	 => std_logic_vector(to_unsigned(107,8) ,
13306	 => std_logic_vector(to_unsigned(104,8) ,
13307	 => std_logic_vector(to_unsigned(105,8) ,
13308	 => std_logic_vector(to_unsigned(108,8) ,
13309	 => std_logic_vector(to_unsigned(103,8) ,
13310	 => std_logic_vector(to_unsigned(97,8) ,
13311	 => std_logic_vector(to_unsigned(96,8) ,
13312	 => std_logic_vector(to_unsigned(104,8) ,
13313	 => std_logic_vector(to_unsigned(115,8) ,
13314	 => std_logic_vector(to_unsigned(100,8) ,
13315	 => std_logic_vector(to_unsigned(99,8) ,
13316	 => std_logic_vector(to_unsigned(99,8) ,
13317	 => std_logic_vector(to_unsigned(87,8) ,
13318	 => std_logic_vector(to_unsigned(92,8) ,
13319	 => std_logic_vector(to_unsigned(118,8) ,
13320	 => std_logic_vector(to_unsigned(124,8) ,
13321	 => std_logic_vector(to_unsigned(116,8) ,
13322	 => std_logic_vector(to_unsigned(103,8) ,
13323	 => std_logic_vector(to_unsigned(96,8) ,
13324	 => std_logic_vector(to_unsigned(114,8) ,
13325	 => std_logic_vector(to_unsigned(134,8) ,
13326	 => std_logic_vector(to_unsigned(99,8) ,
13327	 => std_logic_vector(to_unsigned(80,8) ,
13328	 => std_logic_vector(to_unsigned(87,8) ,
13329	 => std_logic_vector(to_unsigned(84,8) ,
13330	 => std_logic_vector(to_unsigned(86,8) ,
13331	 => std_logic_vector(to_unsigned(91,8) ,
13332	 => std_logic_vector(to_unsigned(87,8) ,
13333	 => std_logic_vector(to_unsigned(86,8) ,
13334	 => std_logic_vector(to_unsigned(86,8) ,
13335	 => std_logic_vector(to_unsigned(79,8) ,
13336	 => std_logic_vector(to_unsigned(88,8) ,
13337	 => std_logic_vector(to_unsigned(90,8) ,
13338	 => std_logic_vector(to_unsigned(93,8) ,
13339	 => std_logic_vector(to_unsigned(105,8) ,
13340	 => std_logic_vector(to_unsigned(107,8) ,
13341	 => std_logic_vector(to_unsigned(116,8) ,
13342	 => std_logic_vector(to_unsigned(124,8) ,
13343	 => std_logic_vector(to_unsigned(131,8) ,
13344	 => std_logic_vector(to_unsigned(115,8) ,
13345	 => std_logic_vector(to_unsigned(92,8) ,
13346	 => std_logic_vector(to_unsigned(86,8) ,
13347	 => std_logic_vector(to_unsigned(81,8) ,
13348	 => std_logic_vector(to_unsigned(82,8) ,
13349	 => std_logic_vector(to_unsigned(82,8) ,
13350	 => std_logic_vector(to_unsigned(86,8) ,
13351	 => std_logic_vector(to_unsigned(82,8) ,
13352	 => std_logic_vector(to_unsigned(88,8) ,
13353	 => std_logic_vector(to_unsigned(101,8) ,
13354	 => std_logic_vector(to_unsigned(103,8) ,
13355	 => std_logic_vector(to_unsigned(92,8) ,
13356	 => std_logic_vector(to_unsigned(87,8) ,
13357	 => std_logic_vector(to_unsigned(85,8) ,
13358	 => std_logic_vector(to_unsigned(84,8) ,
13359	 => std_logic_vector(to_unsigned(77,8) ,
13360	 => std_logic_vector(to_unsigned(71,8) ,
13361	 => std_logic_vector(to_unsigned(74,8) ,
13362	 => std_logic_vector(to_unsigned(63,8) ,
13363	 => std_logic_vector(to_unsigned(51,8) ,
13364	 => std_logic_vector(to_unsigned(48,8) ,
13365	 => std_logic_vector(to_unsigned(13,8) ,
13366	 => std_logic_vector(to_unsigned(0,8) ,
13367	 => std_logic_vector(to_unsigned(0,8) ,
13368	 => std_logic_vector(to_unsigned(3,8) ,
13369	 => std_logic_vector(to_unsigned(44,8) ,
13370	 => std_logic_vector(to_unsigned(50,8) ,
13371	 => std_logic_vector(to_unsigned(46,8) ,
13372	 => std_logic_vector(to_unsigned(45,8) ,
13373	 => std_logic_vector(to_unsigned(51,8) ,
13374	 => std_logic_vector(to_unsigned(48,8) ,
13375	 => std_logic_vector(to_unsigned(54,8) ,
13376	 => std_logic_vector(to_unsigned(52,8) ,
13377	 => std_logic_vector(to_unsigned(45,8) ,
13378	 => std_logic_vector(to_unsigned(38,8) ,
13379	 => std_logic_vector(to_unsigned(45,8) ,
13380	 => std_logic_vector(to_unsigned(53,8) ,
13381	 => std_logic_vector(to_unsigned(51,8) ,
13382	 => std_logic_vector(to_unsigned(51,8) ,
13383	 => std_logic_vector(to_unsigned(63,8) ,
13384	 => std_logic_vector(to_unsigned(86,8) ,
13385	 => std_logic_vector(to_unsigned(84,8) ,
13386	 => std_logic_vector(to_unsigned(61,8) ,
13387	 => std_logic_vector(to_unsigned(65,8) ,
13388	 => std_logic_vector(to_unsigned(66,8) ,
13389	 => std_logic_vector(to_unsigned(73,8) ,
13390	 => std_logic_vector(to_unsigned(67,8) ,
13391	 => std_logic_vector(to_unsigned(52,8) ,
13392	 => std_logic_vector(to_unsigned(53,8) ,
13393	 => std_logic_vector(to_unsigned(58,8) ,
13394	 => std_logic_vector(to_unsigned(57,8) ,
13395	 => std_logic_vector(to_unsigned(51,8) ,
13396	 => std_logic_vector(to_unsigned(55,8) ,
13397	 => std_logic_vector(to_unsigned(52,8) ,
13398	 => std_logic_vector(to_unsigned(54,8) ,
13399	 => std_logic_vector(to_unsigned(67,8) ,
13400	 => std_logic_vector(to_unsigned(70,8) ,
13401	 => std_logic_vector(to_unsigned(78,8) ,
13402	 => std_logic_vector(to_unsigned(88,8) ,
13403	 => std_logic_vector(to_unsigned(78,8) ,
13404	 => std_logic_vector(to_unsigned(82,8) ,
13405	 => std_logic_vector(to_unsigned(92,8) ,
13406	 => std_logic_vector(to_unsigned(91,8) ,
13407	 => std_logic_vector(to_unsigned(86,8) ,
13408	 => std_logic_vector(to_unsigned(88,8) ,
13409	 => std_logic_vector(to_unsigned(87,8) ,
13410	 => std_logic_vector(to_unsigned(88,8) ,
13411	 => std_logic_vector(to_unsigned(95,8) ,
13412	 => std_logic_vector(to_unsigned(104,8) ,
13413	 => std_logic_vector(to_unsigned(116,8) ,
13414	 => std_logic_vector(to_unsigned(115,8) ,
13415	 => std_logic_vector(to_unsigned(130,8) ,
13416	 => std_logic_vector(to_unsigned(146,8) ,
13417	 => std_logic_vector(to_unsigned(154,8) ,
13418	 => std_logic_vector(to_unsigned(159,8) ,
13419	 => std_logic_vector(to_unsigned(151,8) ,
13420	 => std_logic_vector(to_unsigned(161,8) ,
13421	 => std_logic_vector(to_unsigned(161,8) ,
13422	 => std_logic_vector(to_unsigned(154,8) ,
13423	 => std_logic_vector(to_unsigned(157,8) ,
13424	 => std_logic_vector(to_unsigned(161,8) ,
13425	 => std_logic_vector(to_unsigned(161,8) ,
13426	 => std_logic_vector(to_unsigned(163,8) ,
13427	 => std_logic_vector(to_unsigned(161,8) ,
13428	 => std_logic_vector(to_unsigned(164,8) ,
13429	 => std_logic_vector(to_unsigned(159,8) ,
13430	 => std_logic_vector(to_unsigned(163,8) ,
13431	 => std_logic_vector(to_unsigned(156,8) ,
13432	 => std_logic_vector(to_unsigned(136,8) ,
13433	 => std_logic_vector(to_unsigned(141,8) ,
13434	 => std_logic_vector(to_unsigned(142,8) ,
13435	 => std_logic_vector(to_unsigned(130,8) ,
13436	 => std_logic_vector(to_unsigned(125,8) ,
13437	 => std_logic_vector(to_unsigned(122,8) ,
13438	 => std_logic_vector(to_unsigned(127,8) ,
13439	 => std_logic_vector(to_unsigned(142,8) ,
13440	 => std_logic_vector(to_unsigned(151,8) ,
13441	 => std_logic_vector(to_unsigned(154,8) ,
13442	 => std_logic_vector(to_unsigned(151,8) ,
13443	 => std_logic_vector(to_unsigned(152,8) ,
13444	 => std_logic_vector(to_unsigned(151,8) ,
13445	 => std_logic_vector(to_unsigned(149,8) ,
13446	 => std_logic_vector(to_unsigned(147,8) ,
13447	 => std_logic_vector(to_unsigned(119,8) ,
13448	 => std_logic_vector(to_unsigned(127,8) ,
13449	 => std_logic_vector(to_unsigned(154,8) ,
13450	 => std_logic_vector(to_unsigned(152,8) ,
13451	 => std_logic_vector(to_unsigned(154,8) ,
13452	 => std_logic_vector(to_unsigned(152,8) ,
13453	 => std_logic_vector(to_unsigned(147,8) ,
13454	 => std_logic_vector(to_unsigned(149,8) ,
13455	 => std_logic_vector(to_unsigned(151,8) ,
13456	 => std_logic_vector(to_unsigned(157,8) ,
13457	 => std_logic_vector(to_unsigned(164,8) ,
13458	 => std_logic_vector(to_unsigned(156,8) ,
13459	 => std_logic_vector(to_unsigned(144,8) ,
13460	 => std_logic_vector(to_unsigned(156,8) ,
13461	 => std_logic_vector(to_unsigned(163,8) ,
13462	 => std_logic_vector(to_unsigned(159,8) ,
13463	 => std_logic_vector(to_unsigned(164,8) ,
13464	 => std_logic_vector(to_unsigned(161,8) ,
13465	 => std_logic_vector(to_unsigned(159,8) ,
13466	 => std_logic_vector(to_unsigned(157,8) ,
13467	 => std_logic_vector(to_unsigned(159,8) ,
13468	 => std_logic_vector(to_unsigned(152,8) ,
13469	 => std_logic_vector(to_unsigned(125,8) ,
13470	 => std_logic_vector(to_unsigned(116,8) ,
13471	 => std_logic_vector(to_unsigned(119,8) ,
13472	 => std_logic_vector(to_unsigned(122,8) ,
13473	 => std_logic_vector(to_unsigned(118,8) ,
13474	 => std_logic_vector(to_unsigned(121,8) ,
13475	 => std_logic_vector(to_unsigned(115,8) ,
13476	 => std_logic_vector(to_unsigned(119,8) ,
13477	 => std_logic_vector(to_unsigned(116,8) ,
13478	 => std_logic_vector(to_unsigned(130,8) ,
13479	 => std_logic_vector(to_unsigned(127,8) ,
13480	 => std_logic_vector(to_unsigned(134,8) ,
13481	 => std_logic_vector(to_unsigned(138,8) ,
13482	 => std_logic_vector(to_unsigned(134,8) ,
13483	 => std_logic_vector(to_unsigned(134,8) ,
13484	 => std_logic_vector(to_unsigned(128,8) ,
13485	 => std_logic_vector(to_unsigned(130,8) ,
13486	 => std_logic_vector(to_unsigned(122,8) ,
13487	 => std_logic_vector(to_unsigned(121,8) ,
13488	 => std_logic_vector(to_unsigned(130,8) ,
13489	 => std_logic_vector(to_unsigned(130,8) ,
13490	 => std_logic_vector(to_unsigned(144,8) ,
13491	 => std_logic_vector(to_unsigned(138,8) ,
13492	 => std_logic_vector(to_unsigned(139,8) ,
13493	 => std_logic_vector(to_unsigned(154,8) ,
13494	 => std_logic_vector(to_unsigned(156,8) ,
13495	 => std_logic_vector(to_unsigned(156,8) ,
13496	 => std_logic_vector(to_unsigned(152,8) ,
13497	 => std_logic_vector(to_unsigned(142,8) ,
13498	 => std_logic_vector(to_unsigned(149,8) ,
13499	 => std_logic_vector(to_unsigned(147,8) ,
13500	 => std_logic_vector(to_unsigned(144,8) ,
13501	 => std_logic_vector(to_unsigned(151,8) ,
13502	 => std_logic_vector(to_unsigned(151,8) ,
13503	 => std_logic_vector(to_unsigned(138,8) ,
13504	 => std_logic_vector(to_unsigned(128,8) ,
13505	 => std_logic_vector(to_unsigned(134,8) ,
13506	 => std_logic_vector(to_unsigned(134,8) ,
13507	 => std_logic_vector(to_unsigned(136,8) ,
13508	 => std_logic_vector(to_unsigned(128,8) ,
13509	 => std_logic_vector(to_unsigned(121,8) ,
13510	 => std_logic_vector(to_unsigned(125,8) ,
13511	 => std_logic_vector(to_unsigned(127,8) ,
13512	 => std_logic_vector(to_unsigned(130,8) ,
13513	 => std_logic_vector(to_unsigned(124,8) ,
13514	 => std_logic_vector(to_unsigned(138,8) ,
13515	 => std_logic_vector(to_unsigned(138,8) ,
13516	 => std_logic_vector(to_unsigned(95,8) ,
13517	 => std_logic_vector(to_unsigned(96,8) ,
13518	 => std_logic_vector(to_unsigned(105,8) ,
13519	 => std_logic_vector(to_unsigned(109,8) ,
13520	 => std_logic_vector(to_unsigned(119,8) ,
13521	 => std_logic_vector(to_unsigned(127,8) ,
13522	 => std_logic_vector(to_unsigned(131,8) ,
13523	 => std_logic_vector(to_unsigned(136,8) ,
13524	 => std_logic_vector(to_unsigned(131,8) ,
13525	 => std_logic_vector(to_unsigned(138,8) ,
13526	 => std_logic_vector(to_unsigned(139,8) ,
13527	 => std_logic_vector(to_unsigned(131,8) ,
13528	 => std_logic_vector(to_unsigned(138,8) ,
13529	 => std_logic_vector(to_unsigned(134,8) ,
13530	 => std_logic_vector(to_unsigned(141,8) ,
13531	 => std_logic_vector(to_unsigned(168,8) ,
13532	 => std_logic_vector(to_unsigned(168,8) ,
13533	 => std_logic_vector(to_unsigned(144,8) ,
13534	 => std_logic_vector(to_unsigned(131,8) ,
13535	 => std_logic_vector(to_unsigned(141,8) ,
13536	 => std_logic_vector(to_unsigned(151,8) ,
13537	 => std_logic_vector(to_unsigned(142,8) ,
13538	 => std_logic_vector(to_unsigned(134,8) ,
13539	 => std_logic_vector(to_unsigned(138,8) ,
13540	 => std_logic_vector(to_unsigned(144,8) ,
13541	 => std_logic_vector(to_unsigned(146,8) ,
13542	 => std_logic_vector(to_unsigned(136,8) ,
13543	 => std_logic_vector(to_unsigned(142,8) ,
13544	 => std_logic_vector(to_unsigned(134,8) ,
13545	 => std_logic_vector(to_unsigned(121,8) ,
13546	 => std_logic_vector(to_unsigned(125,8) ,
13547	 => std_logic_vector(to_unsigned(114,8) ,
13548	 => std_logic_vector(to_unsigned(118,8) ,
13549	 => std_logic_vector(to_unsigned(121,8) ,
13550	 => std_logic_vector(to_unsigned(114,8) ,
13551	 => std_logic_vector(to_unsigned(103,8) ,
13552	 => std_logic_vector(to_unsigned(97,8) ,
13553	 => std_logic_vector(to_unsigned(97,8) ,
13554	 => std_logic_vector(to_unsigned(96,8) ,
13555	 => std_logic_vector(to_unsigned(96,8) ,
13556	 => std_logic_vector(to_unsigned(95,8) ,
13557	 => std_logic_vector(to_unsigned(112,8) ,
13558	 => std_logic_vector(to_unsigned(134,8) ,
13559	 => std_logic_vector(to_unsigned(130,8) ,
13560	 => std_logic_vector(to_unsigned(116,8) ,
13561	 => std_logic_vector(to_unsigned(125,8) ,
13562	 => std_logic_vector(to_unsigned(130,8) ,
13563	 => std_logic_vector(to_unsigned(124,8) ,
13564	 => std_logic_vector(to_unsigned(134,8) ,
13565	 => std_logic_vector(to_unsigned(146,8) ,
13566	 => std_logic_vector(to_unsigned(130,8) ,
13567	 => std_logic_vector(to_unsigned(122,8) ,
13568	 => std_logic_vector(to_unsigned(152,8) ,
13569	 => std_logic_vector(to_unsigned(157,8) ,
13570	 => std_logic_vector(to_unsigned(146,8) ,
13571	 => std_logic_vector(to_unsigned(144,8) ,
13572	 => std_logic_vector(to_unsigned(147,8) ,
13573	 => std_logic_vector(to_unsigned(133,8) ,
13574	 => std_logic_vector(to_unsigned(125,8) ,
13575	 => std_logic_vector(to_unsigned(125,8) ,
13576	 => std_logic_vector(to_unsigned(118,8) ,
13577	 => std_logic_vector(to_unsigned(107,8) ,
13578	 => std_logic_vector(to_unsigned(109,8) ,
13579	 => std_logic_vector(to_unsigned(118,8) ,
13580	 => std_logic_vector(to_unsigned(118,8) ,
13581	 => std_logic_vector(to_unsigned(112,8) ,
13582	 => std_logic_vector(to_unsigned(108,8) ,
13583	 => std_logic_vector(to_unsigned(104,8) ,
13584	 => std_logic_vector(to_unsigned(109,8) ,
13585	 => std_logic_vector(to_unsigned(118,8) ,
13586	 => std_logic_vector(to_unsigned(121,8) ,
13587	 => std_logic_vector(to_unsigned(119,8) ,
13588	 => std_logic_vector(to_unsigned(118,8) ,
13589	 => std_logic_vector(to_unsigned(119,8) ,
13590	 => std_logic_vector(to_unsigned(114,8) ,
13591	 => std_logic_vector(to_unsigned(109,8) ,
13592	 => std_logic_vector(to_unsigned(100,8) ,
13593	 => std_logic_vector(to_unsigned(100,8) ,
13594	 => std_logic_vector(to_unsigned(88,8) ,
13595	 => std_logic_vector(to_unsigned(80,8) ,
13596	 => std_logic_vector(to_unsigned(105,8) ,
13597	 => std_logic_vector(to_unsigned(104,8) ,
13598	 => std_logic_vector(to_unsigned(95,8) ,
13599	 => std_logic_vector(to_unsigned(96,8) ,
13600	 => std_logic_vector(to_unsigned(86,8) ,
13601	 => std_logic_vector(to_unsigned(95,8) ,
13602	 => std_logic_vector(to_unsigned(104,8) ,
13603	 => std_logic_vector(to_unsigned(93,8) ,
13604	 => std_logic_vector(to_unsigned(95,8) ,
13605	 => std_logic_vector(to_unsigned(91,8) ,
13606	 => std_logic_vector(to_unsigned(91,8) ,
13607	 => std_logic_vector(to_unsigned(96,8) ,
13608	 => std_logic_vector(to_unsigned(70,8) ,
13609	 => std_logic_vector(to_unsigned(55,8) ,
13610	 => std_logic_vector(to_unsigned(55,8) ,
13611	 => std_logic_vector(to_unsigned(73,8) ,
13612	 => std_logic_vector(to_unsigned(118,8) ,
13613	 => std_logic_vector(to_unsigned(99,8) ,
13614	 => std_logic_vector(to_unsigned(84,8) ,
13615	 => std_logic_vector(to_unsigned(92,8) ,
13616	 => std_logic_vector(to_unsigned(95,8) ,
13617	 => std_logic_vector(to_unsigned(92,8) ,
13618	 => std_logic_vector(to_unsigned(95,8) ,
13619	 => std_logic_vector(to_unsigned(92,8) ,
13620	 => std_logic_vector(to_unsigned(74,8) ,
13621	 => std_logic_vector(to_unsigned(79,8) ,
13622	 => std_logic_vector(to_unsigned(99,8) ,
13623	 => std_logic_vector(to_unsigned(111,8) ,
13624	 => std_logic_vector(to_unsigned(105,8) ,
13625	 => std_logic_vector(to_unsigned(109,8) ,
13626	 => std_logic_vector(to_unsigned(93,8) ,
13627	 => std_logic_vector(to_unsigned(91,8) ,
13628	 => std_logic_vector(to_unsigned(108,8) ,
13629	 => std_logic_vector(to_unsigned(103,8) ,
13630	 => std_logic_vector(to_unsigned(92,8) ,
13631	 => std_logic_vector(to_unsigned(107,8) ,
13632	 => std_logic_vector(to_unsigned(112,8) ,
13633	 => std_logic_vector(to_unsigned(122,8) ,
13634	 => std_logic_vector(to_unsigned(118,8) ,
13635	 => std_logic_vector(to_unsigned(96,8) ,
13636	 => std_logic_vector(to_unsigned(104,8) ,
13637	 => std_logic_vector(to_unsigned(115,8) ,
13638	 => std_logic_vector(to_unsigned(107,8) ,
13639	 => std_logic_vector(to_unsigned(116,8) ,
13640	 => std_logic_vector(to_unsigned(118,8) ,
13641	 => std_logic_vector(to_unsigned(108,8) ,
13642	 => std_logic_vector(to_unsigned(103,8) ,
13643	 => std_logic_vector(to_unsigned(99,8) ,
13644	 => std_logic_vector(to_unsigned(101,8) ,
13645	 => std_logic_vector(to_unsigned(118,8) ,
13646	 => std_logic_vector(to_unsigned(104,8) ,
13647	 => std_logic_vector(to_unsigned(88,8) ,
13648	 => std_logic_vector(to_unsigned(82,8) ,
13649	 => std_logic_vector(to_unsigned(86,8) ,
13650	 => std_logic_vector(to_unsigned(84,8) ,
13651	 => std_logic_vector(to_unsigned(91,8) ,
13652	 => std_logic_vector(to_unsigned(78,8) ,
13653	 => std_logic_vector(to_unsigned(71,8) ,
13654	 => std_logic_vector(to_unsigned(66,8) ,
13655	 => std_logic_vector(to_unsigned(63,8) ,
13656	 => std_logic_vector(to_unsigned(79,8) ,
13657	 => std_logic_vector(to_unsigned(101,8) ,
13658	 => std_logic_vector(to_unsigned(100,8) ,
13659	 => std_logic_vector(to_unsigned(81,8) ,
13660	 => std_logic_vector(to_unsigned(78,8) ,
13661	 => std_logic_vector(to_unsigned(91,8) ,
13662	 => std_logic_vector(to_unsigned(124,8) ,
13663	 => std_logic_vector(to_unsigned(134,8) ,
13664	 => std_logic_vector(to_unsigned(121,8) ,
13665	 => std_logic_vector(to_unsigned(101,8) ,
13666	 => std_logic_vector(to_unsigned(84,8) ,
13667	 => std_logic_vector(to_unsigned(73,8) ,
13668	 => std_logic_vector(to_unsigned(71,8) ,
13669	 => std_logic_vector(to_unsigned(93,8) ,
13670	 => std_logic_vector(to_unsigned(87,8) ,
13671	 => std_logic_vector(to_unsigned(85,8) ,
13672	 => std_logic_vector(to_unsigned(101,8) ,
13673	 => std_logic_vector(to_unsigned(111,8) ,
13674	 => std_logic_vector(to_unsigned(107,8) ,
13675	 => std_logic_vector(to_unsigned(100,8) ,
13676	 => std_logic_vector(to_unsigned(103,8) ,
13677	 => std_logic_vector(to_unsigned(107,8) ,
13678	 => std_logic_vector(to_unsigned(87,8) ,
13679	 => std_logic_vector(to_unsigned(74,8) ,
13680	 => std_logic_vector(to_unsigned(70,8) ,
13681	 => std_logic_vector(to_unsigned(64,8) ,
13682	 => std_logic_vector(to_unsigned(55,8) ,
13683	 => std_logic_vector(to_unsigned(46,8) ,
13684	 => std_logic_vector(to_unsigned(58,8) ,
13685	 => std_logic_vector(to_unsigned(28,8) ,
13686	 => std_logic_vector(to_unsigned(1,8) ,
13687	 => std_logic_vector(to_unsigned(0,8) ,
13688	 => std_logic_vector(to_unsigned(1,8) ,
13689	 => std_logic_vector(to_unsigned(29,8) ,
13690	 => std_logic_vector(to_unsigned(56,8) ,
13691	 => std_logic_vector(to_unsigned(48,8) ,
13692	 => std_logic_vector(to_unsigned(51,8) ,
13693	 => std_logic_vector(to_unsigned(52,8) ,
13694	 => std_logic_vector(to_unsigned(52,8) ,
13695	 => std_logic_vector(to_unsigned(48,8) ,
13696	 => std_logic_vector(to_unsigned(49,8) ,
13697	 => std_logic_vector(to_unsigned(51,8) ,
13698	 => std_logic_vector(to_unsigned(46,8) ,
13699	 => std_logic_vector(to_unsigned(42,8) ,
13700	 => std_logic_vector(to_unsigned(51,8) ,
13701	 => std_logic_vector(to_unsigned(51,8) ,
13702	 => std_logic_vector(to_unsigned(51,8) ,
13703	 => std_logic_vector(to_unsigned(62,8) ,
13704	 => std_logic_vector(to_unsigned(77,8) ,
13705	 => std_logic_vector(to_unsigned(76,8) ,
13706	 => std_logic_vector(to_unsigned(56,8) ,
13707	 => std_logic_vector(to_unsigned(71,8) ,
13708	 => std_logic_vector(to_unsigned(82,8) ,
13709	 => std_logic_vector(to_unsigned(78,8) ,
13710	 => std_logic_vector(to_unsigned(62,8) ,
13711	 => std_logic_vector(to_unsigned(48,8) ,
13712	 => std_logic_vector(to_unsigned(51,8) ,
13713	 => std_logic_vector(to_unsigned(59,8) ,
13714	 => std_logic_vector(to_unsigned(56,8) ,
13715	 => std_logic_vector(to_unsigned(58,8) ,
13716	 => std_logic_vector(to_unsigned(62,8) ,
13717	 => std_logic_vector(to_unsigned(65,8) ,
13718	 => std_logic_vector(to_unsigned(65,8) ,
13719	 => std_logic_vector(to_unsigned(67,8) ,
13720	 => std_logic_vector(to_unsigned(66,8) ,
13721	 => std_logic_vector(to_unsigned(69,8) ,
13722	 => std_logic_vector(to_unsigned(91,8) ,
13723	 => std_logic_vector(to_unsigned(85,8) ,
13724	 => std_logic_vector(to_unsigned(81,8) ,
13725	 => std_logic_vector(to_unsigned(80,8) ,
13726	 => std_logic_vector(to_unsigned(84,8) ,
13727	 => std_logic_vector(to_unsigned(79,8) ,
13728	 => std_logic_vector(to_unsigned(77,8) ,
13729	 => std_logic_vector(to_unsigned(88,8) ,
13730	 => std_logic_vector(to_unsigned(104,8) ,
13731	 => std_logic_vector(to_unsigned(119,8) ,
13732	 => std_logic_vector(to_unsigned(119,8) ,
13733	 => std_logic_vector(to_unsigned(111,8) ,
13734	 => std_logic_vector(to_unsigned(114,8) ,
13735	 => std_logic_vector(to_unsigned(141,8) ,
13736	 => std_logic_vector(to_unsigned(156,8) ,
13737	 => std_logic_vector(to_unsigned(154,8) ,
13738	 => std_logic_vector(to_unsigned(161,8) ,
13739	 => std_logic_vector(to_unsigned(157,8) ,
13740	 => std_logic_vector(to_unsigned(161,8) ,
13741	 => std_logic_vector(to_unsigned(159,8) ,
13742	 => std_logic_vector(to_unsigned(161,8) ,
13743	 => std_logic_vector(to_unsigned(159,8) ,
13744	 => std_logic_vector(to_unsigned(163,8) ,
13745	 => std_logic_vector(to_unsigned(164,8) ,
13746	 => std_logic_vector(to_unsigned(159,8) ,
13747	 => std_logic_vector(to_unsigned(159,8) ,
13748	 => std_logic_vector(to_unsigned(161,8) ,
13749	 => std_logic_vector(to_unsigned(152,8) ,
13750	 => std_logic_vector(to_unsigned(147,8) ,
13751	 => std_logic_vector(to_unsigned(142,8) ,
13752	 => std_logic_vector(to_unsigned(128,8) ,
13753	 => std_logic_vector(to_unsigned(127,8) ,
13754	 => std_logic_vector(to_unsigned(128,8) ,
13755	 => std_logic_vector(to_unsigned(125,8) ,
13756	 => std_logic_vector(to_unsigned(134,8) ,
13757	 => std_logic_vector(to_unsigned(134,8) ,
13758	 => std_logic_vector(to_unsigned(142,8) ,
13759	 => std_logic_vector(to_unsigned(152,8) ,
13760	 => std_logic_vector(to_unsigned(152,8) ,
13761	 => std_logic_vector(to_unsigned(142,8) ,
13762	 => std_logic_vector(to_unsigned(142,8) ,
13763	 => std_logic_vector(to_unsigned(149,8) ,
13764	 => std_logic_vector(to_unsigned(144,8) ,
13765	 => std_logic_vector(to_unsigned(147,8) ,
13766	 => std_logic_vector(to_unsigned(152,8) ,
13767	 => std_logic_vector(to_unsigned(134,8) ,
13768	 => std_logic_vector(to_unsigned(133,8) ,
13769	 => std_logic_vector(to_unsigned(139,8) ,
13770	 => std_logic_vector(to_unsigned(144,8) ,
13771	 => std_logic_vector(to_unsigned(147,8) ,
13772	 => std_logic_vector(to_unsigned(151,8) ,
13773	 => std_logic_vector(to_unsigned(142,8) ,
13774	 => std_logic_vector(to_unsigned(139,8) ,
13775	 => std_logic_vector(to_unsigned(147,8) ,
13776	 => std_logic_vector(to_unsigned(149,8) ,
13777	 => std_logic_vector(to_unsigned(159,8) ,
13778	 => std_logic_vector(to_unsigned(152,8) ,
13779	 => std_logic_vector(to_unsigned(138,8) ,
13780	 => std_logic_vector(to_unsigned(146,8) ,
13781	 => std_logic_vector(to_unsigned(156,8) ,
13782	 => std_logic_vector(to_unsigned(157,8) ,
13783	 => std_logic_vector(to_unsigned(163,8) ,
13784	 => std_logic_vector(to_unsigned(161,8) ,
13785	 => std_logic_vector(to_unsigned(157,8) ,
13786	 => std_logic_vector(to_unsigned(161,8) ,
13787	 => std_logic_vector(to_unsigned(164,8) ,
13788	 => std_logic_vector(to_unsigned(152,8) ,
13789	 => std_logic_vector(to_unsigned(125,8) ,
13790	 => std_logic_vector(to_unsigned(115,8) ,
13791	 => std_logic_vector(to_unsigned(124,8) ,
13792	 => std_logic_vector(to_unsigned(128,8) ,
13793	 => std_logic_vector(to_unsigned(122,8) ,
13794	 => std_logic_vector(to_unsigned(122,8) ,
13795	 => std_logic_vector(to_unsigned(118,8) ,
13796	 => std_logic_vector(to_unsigned(116,8) ,
13797	 => std_logic_vector(to_unsigned(119,8) ,
13798	 => std_logic_vector(to_unsigned(127,8) ,
13799	 => std_logic_vector(to_unsigned(127,8) ,
13800	 => std_logic_vector(to_unsigned(138,8) ,
13801	 => std_logic_vector(to_unsigned(130,8) ,
13802	 => std_logic_vector(to_unsigned(121,8) ,
13803	 => std_logic_vector(to_unsigned(128,8) ,
13804	 => std_logic_vector(to_unsigned(136,8) ,
13805	 => std_logic_vector(to_unsigned(131,8) ,
13806	 => std_logic_vector(to_unsigned(128,8) ,
13807	 => std_logic_vector(to_unsigned(125,8) ,
13808	 => std_logic_vector(to_unsigned(130,8) ,
13809	 => std_logic_vector(to_unsigned(134,8) ,
13810	 => std_logic_vector(to_unsigned(142,8) ,
13811	 => std_logic_vector(to_unsigned(146,8) ,
13812	 => std_logic_vector(to_unsigned(151,8) ,
13813	 => std_logic_vector(to_unsigned(156,8) ,
13814	 => std_logic_vector(to_unsigned(156,8) ,
13815	 => std_logic_vector(to_unsigned(154,8) ,
13816	 => std_logic_vector(to_unsigned(151,8) ,
13817	 => std_logic_vector(to_unsigned(138,8) ,
13818	 => std_logic_vector(to_unsigned(142,8) ,
13819	 => std_logic_vector(to_unsigned(154,8) ,
13820	 => std_logic_vector(to_unsigned(151,8) ,
13821	 => std_logic_vector(to_unsigned(149,8) ,
13822	 => std_logic_vector(to_unsigned(152,8) ,
13823	 => std_logic_vector(to_unsigned(154,8) ,
13824	 => std_logic_vector(to_unsigned(147,8) ,
13825	 => std_logic_vector(to_unsigned(146,8) ,
13826	 => std_logic_vector(to_unsigned(151,8) ,
13827	 => std_logic_vector(to_unsigned(152,8) ,
13828	 => std_logic_vector(to_unsigned(146,8) ,
13829	 => std_logic_vector(to_unsigned(124,8) ,
13830	 => std_logic_vector(to_unsigned(124,8) ,
13831	 => std_logic_vector(to_unsigned(136,8) ,
13832	 => std_logic_vector(to_unsigned(134,8) ,
13833	 => std_logic_vector(to_unsigned(124,8) ,
13834	 => std_logic_vector(to_unsigned(133,8) ,
13835	 => std_logic_vector(to_unsigned(133,8) ,
13836	 => std_logic_vector(to_unsigned(97,8) ,
13837	 => std_logic_vector(to_unsigned(105,8) ,
13838	 => std_logic_vector(to_unsigned(133,8) ,
13839	 => std_logic_vector(to_unsigned(124,8) ,
13840	 => std_logic_vector(to_unsigned(121,8) ,
13841	 => std_logic_vector(to_unsigned(119,8) ,
13842	 => std_logic_vector(to_unsigned(107,8) ,
13843	 => std_logic_vector(to_unsigned(107,8) ,
13844	 => std_logic_vector(to_unsigned(116,8) ,
13845	 => std_logic_vector(to_unsigned(127,8) ,
13846	 => std_logic_vector(to_unsigned(125,8) ,
13847	 => std_logic_vector(to_unsigned(136,8) ,
13848	 => std_logic_vector(to_unsigned(138,8) ,
13849	 => std_logic_vector(to_unsigned(139,8) ,
13850	 => std_logic_vector(to_unsigned(146,8) ,
13851	 => std_logic_vector(to_unsigned(161,8) ,
13852	 => std_logic_vector(to_unsigned(164,8) ,
13853	 => std_logic_vector(to_unsigned(156,8) ,
13854	 => std_logic_vector(to_unsigned(151,8) ,
13855	 => std_logic_vector(to_unsigned(149,8) ,
13856	 => std_logic_vector(to_unsigned(147,8) ,
13857	 => std_logic_vector(to_unsigned(149,8) ,
13858	 => std_logic_vector(to_unsigned(151,8) ,
13859	 => std_logic_vector(to_unsigned(147,8) ,
13860	 => std_logic_vector(to_unsigned(146,8) ,
13861	 => std_logic_vector(to_unsigned(149,8) ,
13862	 => std_logic_vector(to_unsigned(146,8) ,
13863	 => std_logic_vector(to_unsigned(138,8) ,
13864	 => std_logic_vector(to_unsigned(133,8) ,
13865	 => std_logic_vector(to_unsigned(128,8) ,
13866	 => std_logic_vector(to_unsigned(124,8) ,
13867	 => std_logic_vector(to_unsigned(121,8) ,
13868	 => std_logic_vector(to_unsigned(128,8) ,
13869	 => std_logic_vector(to_unsigned(115,8) ,
13870	 => std_logic_vector(to_unsigned(104,8) ,
13871	 => std_logic_vector(to_unsigned(103,8) ,
13872	 => std_logic_vector(to_unsigned(108,8) ,
13873	 => std_logic_vector(to_unsigned(105,8) ,
13874	 => std_logic_vector(to_unsigned(93,8) ,
13875	 => std_logic_vector(to_unsigned(93,8) ,
13876	 => std_logic_vector(to_unsigned(100,8) ,
13877	 => std_logic_vector(to_unsigned(108,8) ,
13878	 => std_logic_vector(to_unsigned(105,8) ,
13879	 => std_logic_vector(to_unsigned(99,8) ,
13880	 => std_logic_vector(to_unsigned(105,8) ,
13881	 => std_logic_vector(to_unsigned(122,8) ,
13882	 => std_logic_vector(to_unsigned(130,8) ,
13883	 => std_logic_vector(to_unsigned(116,8) ,
13884	 => std_logic_vector(to_unsigned(121,8) ,
13885	 => std_logic_vector(to_unsigned(141,8) ,
13886	 => std_logic_vector(to_unsigned(136,8) ,
13887	 => std_logic_vector(to_unsigned(115,8) ,
13888	 => std_logic_vector(to_unsigned(133,8) ,
13889	 => std_logic_vector(to_unsigned(144,8) ,
13890	 => std_logic_vector(to_unsigned(133,8) ,
13891	 => std_logic_vector(to_unsigned(151,8) ,
13892	 => std_logic_vector(to_unsigned(152,8) ,
13893	 => std_logic_vector(to_unsigned(147,8) ,
13894	 => std_logic_vector(to_unsigned(147,8) ,
13895	 => std_logic_vector(to_unsigned(134,8) ,
13896	 => std_logic_vector(to_unsigned(134,8) ,
13897	 => std_logic_vector(to_unsigned(119,8) ,
13898	 => std_logic_vector(to_unsigned(100,8) ,
13899	 => std_logic_vector(to_unsigned(101,8) ,
13900	 => std_logic_vector(to_unsigned(97,8) ,
13901	 => std_logic_vector(to_unsigned(104,8) ,
13902	 => std_logic_vector(to_unsigned(104,8) ,
13903	 => std_logic_vector(to_unsigned(96,8) ,
13904	 => std_logic_vector(to_unsigned(101,8) ,
13905	 => std_logic_vector(to_unsigned(109,8) ,
13906	 => std_logic_vector(to_unsigned(116,8) ,
13907	 => std_logic_vector(to_unsigned(109,8) ,
13908	 => std_logic_vector(to_unsigned(105,8) ,
13909	 => std_logic_vector(to_unsigned(114,8) ,
13910	 => std_logic_vector(to_unsigned(105,8) ,
13911	 => std_logic_vector(to_unsigned(100,8) ,
13912	 => std_logic_vector(to_unsigned(93,8) ,
13913	 => std_logic_vector(to_unsigned(97,8) ,
13914	 => std_logic_vector(to_unsigned(92,8) ,
13915	 => std_logic_vector(to_unsigned(86,8) ,
13916	 => std_logic_vector(to_unsigned(93,8) ,
13917	 => std_logic_vector(to_unsigned(87,8) ,
13918	 => std_logic_vector(to_unsigned(97,8) ,
13919	 => std_logic_vector(to_unsigned(99,8) ,
13920	 => std_logic_vector(to_unsigned(97,8) ,
13921	 => std_logic_vector(to_unsigned(90,8) ,
13922	 => std_logic_vector(to_unsigned(78,8) ,
13923	 => std_logic_vector(to_unsigned(77,8) ,
13924	 => std_logic_vector(to_unsigned(95,8) ,
13925	 => std_logic_vector(to_unsigned(99,8) ,
13926	 => std_logic_vector(to_unsigned(91,8) ,
13927	 => std_logic_vector(to_unsigned(92,8) ,
13928	 => std_logic_vector(to_unsigned(85,8) ,
13929	 => std_logic_vector(to_unsigned(78,8) ,
13930	 => std_logic_vector(to_unsigned(85,8) ,
13931	 => std_logic_vector(to_unsigned(88,8) ,
13932	 => std_logic_vector(to_unsigned(105,8) ,
13933	 => std_logic_vector(to_unsigned(92,8) ,
13934	 => std_logic_vector(to_unsigned(85,8) ,
13935	 => std_logic_vector(to_unsigned(88,8) ,
13936	 => std_logic_vector(to_unsigned(96,8) ,
13937	 => std_logic_vector(to_unsigned(101,8) ,
13938	 => std_logic_vector(to_unsigned(103,8) ,
13939	 => std_logic_vector(to_unsigned(99,8) ,
13940	 => std_logic_vector(to_unsigned(80,8) ,
13941	 => std_logic_vector(to_unsigned(74,8) ,
13942	 => std_logic_vector(to_unsigned(86,8) ,
13943	 => std_logic_vector(to_unsigned(101,8) ,
13944	 => std_logic_vector(to_unsigned(103,8) ,
13945	 => std_logic_vector(to_unsigned(109,8) ,
13946	 => std_logic_vector(to_unsigned(86,8) ,
13947	 => std_logic_vector(to_unsigned(81,8) ,
13948	 => std_logic_vector(to_unsigned(114,8) ,
13949	 => std_logic_vector(to_unsigned(97,8) ,
13950	 => std_logic_vector(to_unsigned(95,8) ,
13951	 => std_logic_vector(to_unsigned(111,8) ,
13952	 => std_logic_vector(to_unsigned(101,8) ,
13953	 => std_logic_vector(to_unsigned(112,8) ,
13954	 => std_logic_vector(to_unsigned(108,8) ,
13955	 => std_logic_vector(to_unsigned(87,8) ,
13956	 => std_logic_vector(to_unsigned(96,8) ,
13957	 => std_logic_vector(to_unsigned(111,8) ,
13958	 => std_logic_vector(to_unsigned(97,8) ,
13959	 => std_logic_vector(to_unsigned(99,8) ,
13960	 => std_logic_vector(to_unsigned(96,8) ,
13961	 => std_logic_vector(to_unsigned(99,8) ,
13962	 => std_logic_vector(to_unsigned(111,8) ,
13963	 => std_logic_vector(to_unsigned(103,8) ,
13964	 => std_logic_vector(to_unsigned(86,8) ,
13965	 => std_logic_vector(to_unsigned(93,8) ,
13966	 => std_logic_vector(to_unsigned(109,8) ,
13967	 => std_logic_vector(to_unsigned(100,8) ,
13968	 => std_logic_vector(to_unsigned(80,8) ,
13969	 => std_logic_vector(to_unsigned(81,8) ,
13970	 => std_logic_vector(to_unsigned(77,8) ,
13971	 => std_logic_vector(to_unsigned(79,8) ,
13972	 => std_logic_vector(to_unsigned(74,8) ,
13973	 => std_logic_vector(to_unsigned(66,8) ,
13974	 => std_logic_vector(to_unsigned(49,8) ,
13975	 => std_logic_vector(to_unsigned(58,8) ,
13976	 => std_logic_vector(to_unsigned(84,8) ,
13977	 => std_logic_vector(to_unsigned(109,8) ,
13978	 => std_logic_vector(to_unsigned(108,8) ,
13979	 => std_logic_vector(to_unsigned(121,8) ,
13980	 => std_logic_vector(to_unsigned(134,8) ,
13981	 => std_logic_vector(to_unsigned(125,8) ,
13982	 => std_logic_vector(to_unsigned(108,8) ,
13983	 => std_logic_vector(to_unsigned(109,8) ,
13984	 => std_logic_vector(to_unsigned(115,8) ,
13985	 => std_logic_vector(to_unsigned(86,8) ,
13986	 => std_logic_vector(to_unsigned(81,8) ,
13987	 => std_logic_vector(to_unsigned(76,8) ,
13988	 => std_logic_vector(to_unsigned(56,8) ,
13989	 => std_logic_vector(to_unsigned(85,8) ,
13990	 => std_logic_vector(to_unsigned(72,8) ,
13991	 => std_logic_vector(to_unsigned(79,8) ,
13992	 => std_logic_vector(to_unsigned(99,8) ,
13993	 => std_logic_vector(to_unsigned(105,8) ,
13994	 => std_logic_vector(to_unsigned(107,8) ,
13995	 => std_logic_vector(to_unsigned(96,8) ,
13996	 => std_logic_vector(to_unsigned(85,8) ,
13997	 => std_logic_vector(to_unsigned(77,8) ,
13998	 => std_logic_vector(to_unsigned(63,8) ,
13999	 => std_logic_vector(to_unsigned(62,8) ,
14000	 => std_logic_vector(to_unsigned(63,8) ,
14001	 => std_logic_vector(to_unsigned(46,8) ,
14002	 => std_logic_vector(to_unsigned(45,8) ,
14003	 => std_logic_vector(to_unsigned(58,8) ,
14004	 => std_logic_vector(to_unsigned(67,8) ,
14005	 => std_logic_vector(to_unsigned(44,8) ,
14006	 => std_logic_vector(to_unsigned(3,8) ,
14007	 => std_logic_vector(to_unsigned(0,8) ,
14008	 => std_logic_vector(to_unsigned(0,8) ,
14009	 => std_logic_vector(to_unsigned(19,8) ,
14010	 => std_logic_vector(to_unsigned(66,8) ,
14011	 => std_logic_vector(to_unsigned(56,8) ,
14012	 => std_logic_vector(to_unsigned(54,8) ,
14013	 => std_logic_vector(to_unsigned(57,8) ,
14014	 => std_logic_vector(to_unsigned(63,8) ,
14015	 => std_logic_vector(to_unsigned(54,8) ,
14016	 => std_logic_vector(to_unsigned(47,8) ,
14017	 => std_logic_vector(to_unsigned(50,8) ,
14018	 => std_logic_vector(to_unsigned(51,8) ,
14019	 => std_logic_vector(to_unsigned(56,8) ,
14020	 => std_logic_vector(to_unsigned(56,8) ,
14021	 => std_logic_vector(to_unsigned(60,8) ,
14022	 => std_logic_vector(to_unsigned(67,8) ,
14023	 => std_logic_vector(to_unsigned(66,8) ,
14024	 => std_logic_vector(to_unsigned(56,8) ,
14025	 => std_logic_vector(to_unsigned(60,8) ,
14026	 => std_logic_vector(to_unsigned(56,8) ,
14027	 => std_logic_vector(to_unsigned(67,8) ,
14028	 => std_logic_vector(to_unsigned(67,8) ,
14029	 => std_logic_vector(to_unsigned(60,8) ,
14030	 => std_logic_vector(to_unsigned(61,8) ,
14031	 => std_logic_vector(to_unsigned(60,8) ,
14032	 => std_logic_vector(to_unsigned(63,8) ,
14033	 => std_logic_vector(to_unsigned(63,8) ,
14034	 => std_logic_vector(to_unsigned(60,8) ,
14035	 => std_logic_vector(to_unsigned(63,8) ,
14036	 => std_logic_vector(to_unsigned(67,8) ,
14037	 => std_logic_vector(to_unsigned(67,8) ,
14038	 => std_logic_vector(to_unsigned(66,8) ,
14039	 => std_logic_vector(to_unsigned(61,8) ,
14040	 => std_logic_vector(to_unsigned(64,8) ,
14041	 => std_logic_vector(to_unsigned(67,8) ,
14042	 => std_logic_vector(to_unsigned(76,8) ,
14043	 => std_logic_vector(to_unsigned(76,8) ,
14044	 => std_logic_vector(to_unsigned(77,8) ,
14045	 => std_logic_vector(to_unsigned(78,8) ,
14046	 => std_logic_vector(to_unsigned(91,8) ,
14047	 => std_logic_vector(to_unsigned(86,8) ,
14048	 => std_logic_vector(to_unsigned(100,8) ,
14049	 => std_logic_vector(to_unsigned(130,8) ,
14050	 => std_logic_vector(to_unsigned(139,8) ,
14051	 => std_logic_vector(to_unsigned(125,8) ,
14052	 => std_logic_vector(to_unsigned(127,8) ,
14053	 => std_logic_vector(to_unsigned(131,8) ,
14054	 => std_logic_vector(to_unsigned(128,8) ,
14055	 => std_logic_vector(to_unsigned(125,8) ,
14056	 => std_logic_vector(to_unsigned(139,8) ,
14057	 => std_logic_vector(to_unsigned(154,8) ,
14058	 => std_logic_vector(to_unsigned(147,8) ,
14059	 => std_logic_vector(to_unsigned(157,8) ,
14060	 => std_logic_vector(to_unsigned(156,8) ,
14061	 => std_logic_vector(to_unsigned(156,8) ,
14062	 => std_logic_vector(to_unsigned(161,8) ,
14063	 => std_logic_vector(to_unsigned(151,8) ,
14064	 => std_logic_vector(to_unsigned(157,8) ,
14065	 => std_logic_vector(to_unsigned(159,8) ,
14066	 => std_logic_vector(to_unsigned(163,8) ,
14067	 => std_logic_vector(to_unsigned(157,8) ,
14068	 => std_logic_vector(to_unsigned(156,8) ,
14069	 => std_logic_vector(to_unsigned(154,8) ,
14070	 => std_logic_vector(to_unsigned(147,8) ,
14071	 => std_logic_vector(to_unsigned(151,8) ,
14072	 => std_logic_vector(to_unsigned(149,8) ,
14073	 => std_logic_vector(to_unsigned(151,8) ,
14074	 => std_logic_vector(to_unsigned(147,8) ,
14075	 => std_logic_vector(to_unsigned(152,8) ,
14076	 => std_logic_vector(to_unsigned(156,8) ,
14077	 => std_logic_vector(to_unsigned(159,8) ,
14078	 => std_logic_vector(to_unsigned(161,8) ,
14079	 => std_logic_vector(to_unsigned(161,8) ,
14080	 => std_logic_vector(to_unsigned(164,8) ,
14081	 => std_logic_vector(to_unsigned(125,8) ,
14082	 => std_logic_vector(to_unsigned(125,8) ,
14083	 => std_logic_vector(to_unsigned(133,8) ,
14084	 => std_logic_vector(to_unsigned(136,8) ,
14085	 => std_logic_vector(to_unsigned(136,8) ,
14086	 => std_logic_vector(to_unsigned(144,8) ,
14087	 => std_logic_vector(to_unsigned(133,8) ,
14088	 => std_logic_vector(to_unsigned(124,8) ,
14089	 => std_logic_vector(to_unsigned(125,8) ,
14090	 => std_logic_vector(to_unsigned(128,8) ,
14091	 => std_logic_vector(to_unsigned(141,8) ,
14092	 => std_logic_vector(to_unsigned(146,8) ,
14093	 => std_logic_vector(to_unsigned(141,8) ,
14094	 => std_logic_vector(to_unsigned(141,8) ,
14095	 => std_logic_vector(to_unsigned(147,8) ,
14096	 => std_logic_vector(to_unsigned(146,8) ,
14097	 => std_logic_vector(to_unsigned(151,8) ,
14098	 => std_logic_vector(to_unsigned(147,8) ,
14099	 => std_logic_vector(to_unsigned(134,8) ,
14100	 => std_logic_vector(to_unsigned(133,8) ,
14101	 => std_logic_vector(to_unsigned(142,8) ,
14102	 => std_logic_vector(to_unsigned(147,8) ,
14103	 => std_logic_vector(to_unsigned(146,8) ,
14104	 => std_logic_vector(to_unsigned(152,8) ,
14105	 => std_logic_vector(to_unsigned(154,8) ,
14106	 => std_logic_vector(to_unsigned(159,8) ,
14107	 => std_logic_vector(to_unsigned(159,8) ,
14108	 => std_logic_vector(to_unsigned(149,8) ,
14109	 => std_logic_vector(to_unsigned(131,8) ,
14110	 => std_logic_vector(to_unsigned(127,8) ,
14111	 => std_logic_vector(to_unsigned(131,8) ,
14112	 => std_logic_vector(to_unsigned(125,8) ,
14113	 => std_logic_vector(to_unsigned(130,8) ,
14114	 => std_logic_vector(to_unsigned(130,8) ,
14115	 => std_logic_vector(to_unsigned(119,8) ,
14116	 => std_logic_vector(to_unsigned(109,8) ,
14117	 => std_logic_vector(to_unsigned(122,8) ,
14118	 => std_logic_vector(to_unsigned(127,8) ,
14119	 => std_logic_vector(to_unsigned(136,8) ,
14120	 => std_logic_vector(to_unsigned(147,8) ,
14121	 => std_logic_vector(to_unsigned(146,8) ,
14122	 => std_logic_vector(to_unsigned(144,8) ,
14123	 => std_logic_vector(to_unsigned(128,8) ,
14124	 => std_logic_vector(to_unsigned(130,8) ,
14125	 => std_logic_vector(to_unsigned(130,8) ,
14126	 => std_logic_vector(to_unsigned(128,8) ,
14127	 => std_logic_vector(to_unsigned(128,8) ,
14128	 => std_logic_vector(to_unsigned(136,8) ,
14129	 => std_logic_vector(to_unsigned(141,8) ,
14130	 => std_logic_vector(to_unsigned(139,8) ,
14131	 => std_logic_vector(to_unsigned(152,8) ,
14132	 => std_logic_vector(to_unsigned(154,8) ,
14133	 => std_logic_vector(to_unsigned(156,8) ,
14134	 => std_logic_vector(to_unsigned(154,8) ,
14135	 => std_logic_vector(to_unsigned(156,8) ,
14136	 => std_logic_vector(to_unsigned(152,8) ,
14137	 => std_logic_vector(to_unsigned(144,8) ,
14138	 => std_logic_vector(to_unsigned(144,8) ,
14139	 => std_logic_vector(to_unsigned(154,8) ,
14140	 => std_logic_vector(to_unsigned(154,8) ,
14141	 => std_logic_vector(to_unsigned(149,8) ,
14142	 => std_logic_vector(to_unsigned(152,8) ,
14143	 => std_logic_vector(to_unsigned(156,8) ,
14144	 => std_logic_vector(to_unsigned(156,8) ,
14145	 => std_logic_vector(to_unsigned(156,8) ,
14146	 => std_logic_vector(to_unsigned(161,8) ,
14147	 => std_logic_vector(to_unsigned(154,8) ,
14148	 => std_logic_vector(to_unsigned(163,8) ,
14149	 => std_logic_vector(to_unsigned(125,8) ,
14150	 => std_logic_vector(to_unsigned(104,8) ,
14151	 => std_logic_vector(to_unsigned(122,8) ,
14152	 => std_logic_vector(to_unsigned(119,8) ,
14153	 => std_logic_vector(to_unsigned(111,8) ,
14154	 => std_logic_vector(to_unsigned(107,8) ,
14155	 => std_logic_vector(to_unsigned(108,8) ,
14156	 => std_logic_vector(to_unsigned(114,8) ,
14157	 => std_logic_vector(to_unsigned(136,8) ,
14158	 => std_logic_vector(to_unsigned(134,8) ,
14159	 => std_logic_vector(to_unsigned(136,8) ,
14160	 => std_logic_vector(to_unsigned(134,8) ,
14161	 => std_logic_vector(to_unsigned(138,8) ,
14162	 => std_logic_vector(to_unsigned(127,8) ,
14163	 => std_logic_vector(to_unsigned(122,8) ,
14164	 => std_logic_vector(to_unsigned(139,8) ,
14165	 => std_logic_vector(to_unsigned(149,8) ,
14166	 => std_logic_vector(to_unsigned(147,8) ,
14167	 => std_logic_vector(to_unsigned(149,8) ,
14168	 => std_logic_vector(to_unsigned(149,8) ,
14169	 => std_logic_vector(to_unsigned(149,8) ,
14170	 => std_logic_vector(to_unsigned(152,8) ,
14171	 => std_logic_vector(to_unsigned(152,8) ,
14172	 => std_logic_vector(to_unsigned(151,8) ,
14173	 => std_logic_vector(to_unsigned(161,8) ,
14174	 => std_logic_vector(to_unsigned(163,8) ,
14175	 => std_logic_vector(to_unsigned(157,8) ,
14176	 => std_logic_vector(to_unsigned(156,8) ,
14177	 => std_logic_vector(to_unsigned(151,8) ,
14178	 => std_logic_vector(to_unsigned(157,8) ,
14179	 => std_logic_vector(to_unsigned(152,8) ,
14180	 => std_logic_vector(to_unsigned(147,8) ,
14181	 => std_logic_vector(to_unsigned(149,8) ,
14182	 => std_logic_vector(to_unsigned(147,8) ,
14183	 => std_logic_vector(to_unsigned(139,8) ,
14184	 => std_logic_vector(to_unsigned(147,8) ,
14185	 => std_logic_vector(to_unsigned(152,8) ,
14186	 => std_logic_vector(to_unsigned(128,8) ,
14187	 => std_logic_vector(to_unsigned(131,8) ,
14188	 => std_logic_vector(to_unsigned(142,8) ,
14189	 => std_logic_vector(to_unsigned(112,8) ,
14190	 => std_logic_vector(to_unsigned(93,8) ,
14191	 => std_logic_vector(to_unsigned(112,8) ,
14192	 => std_logic_vector(to_unsigned(116,8) ,
14193	 => std_logic_vector(to_unsigned(111,8) ,
14194	 => std_logic_vector(to_unsigned(109,8) ,
14195	 => std_logic_vector(to_unsigned(108,8) ,
14196	 => std_logic_vector(to_unsigned(112,8) ,
14197	 => std_logic_vector(to_unsigned(105,8) ,
14198	 => std_logic_vector(to_unsigned(108,8) ,
14199	 => std_logic_vector(to_unsigned(115,8) ,
14200	 => std_logic_vector(to_unsigned(104,8) ,
14201	 => std_logic_vector(to_unsigned(104,8) ,
14202	 => std_logic_vector(to_unsigned(119,8) ,
14203	 => std_logic_vector(to_unsigned(130,8) ,
14204	 => std_logic_vector(to_unsigned(128,8) ,
14205	 => std_logic_vector(to_unsigned(133,8) ,
14206	 => std_logic_vector(to_unsigned(119,8) ,
14207	 => std_logic_vector(to_unsigned(101,8) ,
14208	 => std_logic_vector(to_unsigned(116,8) ,
14209	 => std_logic_vector(to_unsigned(115,8) ,
14210	 => std_logic_vector(to_unsigned(114,8) ,
14211	 => std_logic_vector(to_unsigned(144,8) ,
14212	 => std_logic_vector(to_unsigned(154,8) ,
14213	 => std_logic_vector(to_unsigned(152,8) ,
14214	 => std_logic_vector(to_unsigned(152,8) ,
14215	 => std_logic_vector(to_unsigned(134,8) ,
14216	 => std_logic_vector(to_unsigned(127,8) ,
14217	 => std_logic_vector(to_unsigned(112,8) ,
14218	 => std_logic_vector(to_unsigned(99,8) ,
14219	 => std_logic_vector(to_unsigned(100,8) ,
14220	 => std_logic_vector(to_unsigned(105,8) ,
14221	 => std_logic_vector(to_unsigned(118,8) ,
14222	 => std_logic_vector(to_unsigned(112,8) ,
14223	 => std_logic_vector(to_unsigned(92,8) ,
14224	 => std_logic_vector(to_unsigned(97,8) ,
14225	 => std_logic_vector(to_unsigned(96,8) ,
14226	 => std_logic_vector(to_unsigned(105,8) ,
14227	 => std_logic_vector(to_unsigned(115,8) ,
14228	 => std_logic_vector(to_unsigned(101,8) ,
14229	 => std_logic_vector(to_unsigned(99,8) ,
14230	 => std_logic_vector(to_unsigned(91,8) ,
14231	 => std_logic_vector(to_unsigned(90,8) ,
14232	 => std_logic_vector(to_unsigned(87,8) ,
14233	 => std_logic_vector(to_unsigned(84,8) ,
14234	 => std_logic_vector(to_unsigned(88,8) ,
14235	 => std_logic_vector(to_unsigned(90,8) ,
14236	 => std_logic_vector(to_unsigned(80,8) ,
14237	 => std_logic_vector(to_unsigned(67,8) ,
14238	 => std_logic_vector(to_unsigned(65,8) ,
14239	 => std_logic_vector(to_unsigned(67,8) ,
14240	 => std_logic_vector(to_unsigned(107,8) ,
14241	 => std_logic_vector(to_unsigned(107,8) ,
14242	 => std_logic_vector(to_unsigned(88,8) ,
14243	 => std_logic_vector(to_unsigned(92,8) ,
14244	 => std_logic_vector(to_unsigned(90,8) ,
14245	 => std_logic_vector(to_unsigned(90,8) ,
14246	 => std_logic_vector(to_unsigned(85,8) ,
14247	 => std_logic_vector(to_unsigned(82,8) ,
14248	 => std_logic_vector(to_unsigned(92,8) ,
14249	 => std_logic_vector(to_unsigned(100,8) ,
14250	 => std_logic_vector(to_unsigned(86,8) ,
14251	 => std_logic_vector(to_unsigned(67,8) ,
14252	 => std_logic_vector(to_unsigned(69,8) ,
14253	 => std_logic_vector(to_unsigned(73,8) ,
14254	 => std_logic_vector(to_unsigned(86,8) ,
14255	 => std_logic_vector(to_unsigned(90,8) ,
14256	 => std_logic_vector(to_unsigned(91,8) ,
14257	 => std_logic_vector(to_unsigned(99,8) ,
14258	 => std_logic_vector(to_unsigned(104,8) ,
14259	 => std_logic_vector(to_unsigned(96,8) ,
14260	 => std_logic_vector(to_unsigned(82,8) ,
14261	 => std_logic_vector(to_unsigned(80,8) ,
14262	 => std_logic_vector(to_unsigned(91,8) ,
14263	 => std_logic_vector(to_unsigned(107,8) ,
14264	 => std_logic_vector(to_unsigned(101,8) ,
14265	 => std_logic_vector(to_unsigned(108,8) ,
14266	 => std_logic_vector(to_unsigned(88,8) ,
14267	 => std_logic_vector(to_unsigned(79,8) ,
14268	 => std_logic_vector(to_unsigned(118,8) ,
14269	 => std_logic_vector(to_unsigned(114,8) ,
14270	 => std_logic_vector(to_unsigned(107,8) ,
14271	 => std_logic_vector(to_unsigned(108,8) ,
14272	 => std_logic_vector(to_unsigned(97,8) ,
14273	 => std_logic_vector(to_unsigned(92,8) ,
14274	 => std_logic_vector(to_unsigned(91,8) ,
14275	 => std_logic_vector(to_unsigned(95,8) ,
14276	 => std_logic_vector(to_unsigned(97,8) ,
14277	 => std_logic_vector(to_unsigned(104,8) ,
14278	 => std_logic_vector(to_unsigned(99,8) ,
14279	 => std_logic_vector(to_unsigned(103,8) ,
14280	 => std_logic_vector(to_unsigned(90,8) ,
14281	 => std_logic_vector(to_unsigned(101,8) ,
14282	 => std_logic_vector(to_unsigned(109,8) ,
14283	 => std_logic_vector(to_unsigned(99,8) ,
14284	 => std_logic_vector(to_unsigned(93,8) ,
14285	 => std_logic_vector(to_unsigned(104,8) ,
14286	 => std_logic_vector(to_unsigned(116,8) ,
14287	 => std_logic_vector(to_unsigned(99,8) ,
14288	 => std_logic_vector(to_unsigned(92,8) ,
14289	 => std_logic_vector(to_unsigned(96,8) ,
14290	 => std_logic_vector(to_unsigned(65,8) ,
14291	 => std_logic_vector(to_unsigned(61,8) ,
14292	 => std_logic_vector(to_unsigned(62,8) ,
14293	 => std_logic_vector(to_unsigned(56,8) ,
14294	 => std_logic_vector(to_unsigned(48,8) ,
14295	 => std_logic_vector(to_unsigned(62,8) ,
14296	 => std_logic_vector(to_unsigned(84,8) ,
14297	 => std_logic_vector(to_unsigned(101,8) ,
14298	 => std_logic_vector(to_unsigned(108,8) ,
14299	 => std_logic_vector(to_unsigned(141,8) ,
14300	 => std_logic_vector(to_unsigned(164,8) ,
14301	 => std_logic_vector(to_unsigned(151,8) ,
14302	 => std_logic_vector(to_unsigned(109,8) ,
14303	 => std_logic_vector(to_unsigned(107,8) ,
14304	 => std_logic_vector(to_unsigned(108,8) ,
14305	 => std_logic_vector(to_unsigned(60,8) ,
14306	 => std_logic_vector(to_unsigned(60,8) ,
14307	 => std_logic_vector(to_unsigned(64,8) ,
14308	 => std_logic_vector(to_unsigned(51,8) ,
14309	 => std_logic_vector(to_unsigned(67,8) ,
14310	 => std_logic_vector(to_unsigned(70,8) ,
14311	 => std_logic_vector(to_unsigned(84,8) ,
14312	 => std_logic_vector(to_unsigned(93,8) ,
14313	 => std_logic_vector(to_unsigned(86,8) ,
14314	 => std_logic_vector(to_unsigned(79,8) ,
14315	 => std_logic_vector(to_unsigned(74,8) ,
14316	 => std_logic_vector(to_unsigned(64,8) ,
14317	 => std_logic_vector(to_unsigned(62,8) ,
14318	 => std_logic_vector(to_unsigned(60,8) ,
14319	 => std_logic_vector(to_unsigned(52,8) ,
14320	 => std_logic_vector(to_unsigned(51,8) ,
14321	 => std_logic_vector(to_unsigned(45,8) ,
14322	 => std_logic_vector(to_unsigned(47,8) ,
14323	 => std_logic_vector(to_unsigned(55,8) ,
14324	 => std_logic_vector(to_unsigned(53,8) ,
14325	 => std_logic_vector(to_unsigned(55,8) ,
14326	 => std_logic_vector(to_unsigned(12,8) ,
14327	 => std_logic_vector(to_unsigned(0,8) ,
14328	 => std_logic_vector(to_unsigned(0,8) ,
14329	 => std_logic_vector(to_unsigned(6,8) ,
14330	 => std_logic_vector(to_unsigned(55,8) ,
14331	 => std_logic_vector(to_unsigned(68,8) ,
14332	 => std_logic_vector(to_unsigned(62,8) ,
14333	 => std_logic_vector(to_unsigned(64,8) ,
14334	 => std_logic_vector(to_unsigned(62,8) ,
14335	 => std_logic_vector(to_unsigned(60,8) ,
14336	 => std_logic_vector(to_unsigned(52,8) ,
14337	 => std_logic_vector(to_unsigned(62,8) ,
14338	 => std_logic_vector(to_unsigned(64,8) ,
14339	 => std_logic_vector(to_unsigned(67,8) ,
14340	 => std_logic_vector(to_unsigned(76,8) ,
14341	 => std_logic_vector(to_unsigned(85,8) ,
14342	 => std_logic_vector(to_unsigned(87,8) ,
14343	 => std_logic_vector(to_unsigned(65,8) ,
14344	 => std_logic_vector(to_unsigned(52,8) ,
14345	 => std_logic_vector(to_unsigned(59,8) ,
14346	 => std_logic_vector(to_unsigned(54,8) ,
14347	 => std_logic_vector(to_unsigned(62,8) ,
14348	 => std_logic_vector(to_unsigned(64,8) ,
14349	 => std_logic_vector(to_unsigned(62,8) ,
14350	 => std_logic_vector(to_unsigned(82,8) ,
14351	 => std_logic_vector(to_unsigned(92,8) ,
14352	 => std_logic_vector(to_unsigned(80,8) ,
14353	 => std_logic_vector(to_unsigned(69,8) ,
14354	 => std_logic_vector(to_unsigned(56,8) ,
14355	 => std_logic_vector(to_unsigned(58,8) ,
14356	 => std_logic_vector(to_unsigned(67,8) ,
14357	 => std_logic_vector(to_unsigned(70,8) ,
14358	 => std_logic_vector(to_unsigned(64,8) ,
14359	 => std_logic_vector(to_unsigned(59,8) ,
14360	 => std_logic_vector(to_unsigned(70,8) ,
14361	 => std_logic_vector(to_unsigned(76,8) ,
14362	 => std_logic_vector(to_unsigned(80,8) ,
14363	 => std_logic_vector(to_unsigned(77,8) ,
14364	 => std_logic_vector(to_unsigned(74,8) ,
14365	 => std_logic_vector(to_unsigned(79,8) ,
14366	 => std_logic_vector(to_unsigned(93,8) ,
14367	 => std_logic_vector(to_unsigned(91,8) ,
14368	 => std_logic_vector(to_unsigned(99,8) ,
14369	 => std_logic_vector(to_unsigned(125,8) ,
14370	 => std_logic_vector(to_unsigned(131,8) ,
14371	 => std_logic_vector(to_unsigned(133,8) ,
14372	 => std_logic_vector(to_unsigned(128,8) ,
14373	 => std_logic_vector(to_unsigned(133,8) ,
14374	 => std_logic_vector(to_unsigned(136,8) ,
14375	 => std_logic_vector(to_unsigned(99,8) ,
14376	 => std_logic_vector(to_unsigned(124,8) ,
14377	 => std_logic_vector(to_unsigned(161,8) ,
14378	 => std_logic_vector(to_unsigned(141,8) ,
14379	 => std_logic_vector(to_unsigned(142,8) ,
14380	 => std_logic_vector(to_unsigned(152,8) ,
14381	 => std_logic_vector(to_unsigned(154,8) ,
14382	 => std_logic_vector(to_unsigned(147,8) ,
14383	 => std_logic_vector(to_unsigned(141,8) ,
14384	 => std_logic_vector(to_unsigned(146,8) ,
14385	 => std_logic_vector(to_unsigned(152,8) ,
14386	 => std_logic_vector(to_unsigned(154,8) ,
14387	 => std_logic_vector(to_unsigned(154,8) ,
14388	 => std_logic_vector(to_unsigned(154,8) ,
14389	 => std_logic_vector(to_unsigned(154,8) ,
14390	 => std_logic_vector(to_unsigned(156,8) ,
14391	 => std_logic_vector(to_unsigned(159,8) ,
14392	 => std_logic_vector(to_unsigned(161,8) ,
14393	 => std_logic_vector(to_unsigned(166,8) ,
14394	 => std_logic_vector(to_unsigned(168,8) ,
14395	 => std_logic_vector(to_unsigned(171,8) ,
14396	 => std_logic_vector(to_unsigned(164,8) ,
14397	 => std_logic_vector(to_unsigned(159,8) ,
14398	 => std_logic_vector(to_unsigned(163,8) ,
14399	 => std_logic_vector(to_unsigned(157,8) ,
14400	 => std_logic_vector(to_unsigned(159,8) ,
14401	 => std_logic_vector(to_unsigned(139,8) ,
14402	 => std_logic_vector(to_unsigned(136,8) ,
14403	 => std_logic_vector(to_unsigned(133,8) ,
14404	 => std_logic_vector(to_unsigned(134,8) ,
14405	 => std_logic_vector(to_unsigned(125,8) ,
14406	 => std_logic_vector(to_unsigned(142,8) ,
14407	 => std_logic_vector(to_unsigned(141,8) ,
14408	 => std_logic_vector(to_unsigned(133,8) ,
14409	 => std_logic_vector(to_unsigned(131,8) ,
14410	 => std_logic_vector(to_unsigned(128,8) ,
14411	 => std_logic_vector(to_unsigned(144,8) ,
14412	 => std_logic_vector(to_unsigned(138,8) ,
14413	 => std_logic_vector(to_unsigned(136,8) ,
14414	 => std_logic_vector(to_unsigned(141,8) ,
14415	 => std_logic_vector(to_unsigned(141,8) ,
14416	 => std_logic_vector(to_unsigned(151,8) ,
14417	 => std_logic_vector(to_unsigned(146,8) ,
14418	 => std_logic_vector(to_unsigned(133,8) ,
14419	 => std_logic_vector(to_unsigned(133,8) ,
14420	 => std_logic_vector(to_unsigned(142,8) ,
14421	 => std_logic_vector(to_unsigned(147,8) ,
14422	 => std_logic_vector(to_unsigned(144,8) ,
14423	 => std_logic_vector(to_unsigned(134,8) ,
14424	 => std_logic_vector(to_unsigned(151,8) ,
14425	 => std_logic_vector(to_unsigned(157,8) ,
14426	 => std_logic_vector(to_unsigned(151,8) ,
14427	 => std_logic_vector(to_unsigned(146,8) ,
14428	 => std_logic_vector(to_unsigned(141,8) ,
14429	 => std_logic_vector(to_unsigned(130,8) ,
14430	 => std_logic_vector(to_unsigned(138,8) ,
14431	 => std_logic_vector(to_unsigned(142,8) ,
14432	 => std_logic_vector(to_unsigned(134,8) ,
14433	 => std_logic_vector(to_unsigned(136,8) ,
14434	 => std_logic_vector(to_unsigned(133,8) ,
14435	 => std_logic_vector(to_unsigned(130,8) ,
14436	 => std_logic_vector(to_unsigned(133,8) ,
14437	 => std_logic_vector(to_unsigned(131,8) ,
14438	 => std_logic_vector(to_unsigned(134,8) ,
14439	 => std_logic_vector(to_unsigned(154,8) ,
14440	 => std_logic_vector(to_unsigned(146,8) ,
14441	 => std_logic_vector(to_unsigned(133,8) ,
14442	 => std_logic_vector(to_unsigned(134,8) ,
14443	 => std_logic_vector(to_unsigned(115,8) ,
14444	 => std_logic_vector(to_unsigned(114,8) ,
14445	 => std_logic_vector(to_unsigned(133,8) ,
14446	 => std_logic_vector(to_unsigned(136,8) ,
14447	 => std_logic_vector(to_unsigned(134,8) ,
14448	 => std_logic_vector(to_unsigned(141,8) ,
14449	 => std_logic_vector(to_unsigned(141,8) ,
14450	 => std_logic_vector(to_unsigned(144,8) ,
14451	 => std_logic_vector(to_unsigned(149,8) ,
14452	 => std_logic_vector(to_unsigned(152,8) ,
14453	 => std_logic_vector(to_unsigned(154,8) ,
14454	 => std_logic_vector(to_unsigned(154,8) ,
14455	 => std_logic_vector(to_unsigned(154,8) ,
14456	 => std_logic_vector(to_unsigned(149,8) ,
14457	 => std_logic_vector(to_unsigned(146,8) ,
14458	 => std_logic_vector(to_unsigned(151,8) ,
14459	 => std_logic_vector(to_unsigned(154,8) ,
14460	 => std_logic_vector(to_unsigned(152,8) ,
14461	 => std_logic_vector(to_unsigned(146,8) ,
14462	 => std_logic_vector(to_unsigned(151,8) ,
14463	 => std_logic_vector(to_unsigned(159,8) ,
14464	 => std_logic_vector(to_unsigned(157,8) ,
14465	 => std_logic_vector(to_unsigned(161,8) ,
14466	 => std_logic_vector(to_unsigned(157,8) ,
14467	 => std_logic_vector(to_unsigned(157,8) ,
14468	 => std_logic_vector(to_unsigned(159,8) ,
14469	 => std_logic_vector(to_unsigned(133,8) ,
14470	 => std_logic_vector(to_unsigned(114,8) ,
14471	 => std_logic_vector(to_unsigned(130,8) ,
14472	 => std_logic_vector(to_unsigned(134,8) ,
14473	 => std_logic_vector(to_unsigned(127,8) ,
14474	 => std_logic_vector(to_unsigned(114,8) ,
14475	 => std_logic_vector(to_unsigned(108,8) ,
14476	 => std_logic_vector(to_unsigned(115,8) ,
14477	 => std_logic_vector(to_unsigned(134,8) ,
14478	 => std_logic_vector(to_unsigned(115,8) ,
14479	 => std_logic_vector(to_unsigned(136,8) ,
14480	 => std_logic_vector(to_unsigned(144,8) ,
14481	 => std_logic_vector(to_unsigned(136,8) ,
14482	 => std_logic_vector(to_unsigned(133,8) ,
14483	 => std_logic_vector(to_unsigned(131,8) ,
14484	 => std_logic_vector(to_unsigned(131,8) ,
14485	 => std_logic_vector(to_unsigned(138,8) ,
14486	 => std_logic_vector(to_unsigned(149,8) ,
14487	 => std_logic_vector(to_unsigned(154,8) ,
14488	 => std_logic_vector(to_unsigned(157,8) ,
14489	 => std_logic_vector(to_unsigned(161,8) ,
14490	 => std_logic_vector(to_unsigned(157,8) ,
14491	 => std_logic_vector(to_unsigned(151,8) ,
14492	 => std_logic_vector(to_unsigned(152,8) ,
14493	 => std_logic_vector(to_unsigned(164,8) ,
14494	 => std_logic_vector(to_unsigned(173,8) ,
14495	 => std_logic_vector(to_unsigned(173,8) ,
14496	 => std_logic_vector(to_unsigned(175,8) ,
14497	 => std_logic_vector(to_unsigned(163,8) ,
14498	 => std_logic_vector(to_unsigned(157,8) ,
14499	 => std_logic_vector(to_unsigned(154,8) ,
14500	 => std_logic_vector(to_unsigned(152,8) ,
14501	 => std_logic_vector(to_unsigned(149,8) ,
14502	 => std_logic_vector(to_unsigned(149,8) ,
14503	 => std_logic_vector(to_unsigned(149,8) ,
14504	 => std_logic_vector(to_unsigned(161,8) ,
14505	 => std_logic_vector(to_unsigned(170,8) ,
14506	 => std_logic_vector(to_unsigned(134,8) ,
14507	 => std_logic_vector(to_unsigned(118,8) ,
14508	 => std_logic_vector(to_unsigned(125,8) ,
14509	 => std_logic_vector(to_unsigned(121,8) ,
14510	 => std_logic_vector(to_unsigned(114,8) ,
14511	 => std_logic_vector(to_unsigned(114,8) ,
14512	 => std_logic_vector(to_unsigned(107,8) ,
14513	 => std_logic_vector(to_unsigned(97,8) ,
14514	 => std_logic_vector(to_unsigned(93,8) ,
14515	 => std_logic_vector(to_unsigned(99,8) ,
14516	 => std_logic_vector(to_unsigned(104,8) ,
14517	 => std_logic_vector(to_unsigned(114,8) ,
14518	 => std_logic_vector(to_unsigned(125,8) ,
14519	 => std_logic_vector(to_unsigned(124,8) ,
14520	 => std_logic_vector(to_unsigned(114,8) ,
14521	 => std_logic_vector(to_unsigned(115,8) ,
14522	 => std_logic_vector(to_unsigned(125,8) ,
14523	 => std_logic_vector(to_unsigned(128,8) ,
14524	 => std_logic_vector(to_unsigned(119,8) ,
14525	 => std_logic_vector(to_unsigned(111,8) ,
14526	 => std_logic_vector(to_unsigned(99,8) ,
14527	 => std_logic_vector(to_unsigned(93,8) ,
14528	 => std_logic_vector(to_unsigned(108,8) ,
14529	 => std_logic_vector(to_unsigned(119,8) ,
14530	 => std_logic_vector(to_unsigned(115,8) ,
14531	 => std_logic_vector(to_unsigned(142,8) ,
14532	 => std_logic_vector(to_unsigned(152,8) ,
14533	 => std_logic_vector(to_unsigned(144,8) ,
14534	 => std_logic_vector(to_unsigned(133,8) ,
14535	 => std_logic_vector(to_unsigned(119,8) ,
14536	 => std_logic_vector(to_unsigned(108,8) ,
14537	 => std_logic_vector(to_unsigned(95,8) ,
14538	 => std_logic_vector(to_unsigned(104,8) ,
14539	 => std_logic_vector(to_unsigned(109,8) ,
14540	 => std_logic_vector(to_unsigned(112,8) ,
14541	 => std_logic_vector(to_unsigned(125,8) ,
14542	 => std_logic_vector(to_unsigned(128,8) ,
14543	 => std_logic_vector(to_unsigned(114,8) ,
14544	 => std_logic_vector(to_unsigned(112,8) ,
14545	 => std_logic_vector(to_unsigned(121,8) ,
14546	 => std_logic_vector(to_unsigned(134,8) ,
14547	 => std_logic_vector(to_unsigned(142,8) ,
14548	 => std_logic_vector(to_unsigned(104,8) ,
14549	 => std_logic_vector(to_unsigned(85,8) ,
14550	 => std_logic_vector(to_unsigned(87,8) ,
14551	 => std_logic_vector(to_unsigned(99,8) ,
14552	 => std_logic_vector(to_unsigned(105,8) ,
14553	 => std_logic_vector(to_unsigned(100,8) ,
14554	 => std_logic_vector(to_unsigned(92,8) ,
14555	 => std_logic_vector(to_unsigned(92,8) ,
14556	 => std_logic_vector(to_unsigned(88,8) ,
14557	 => std_logic_vector(to_unsigned(77,8) ,
14558	 => std_logic_vector(to_unsigned(68,8) ,
14559	 => std_logic_vector(to_unsigned(74,8) ,
14560	 => std_logic_vector(to_unsigned(84,8) ,
14561	 => std_logic_vector(to_unsigned(90,8) ,
14562	 => std_logic_vector(to_unsigned(104,8) ,
14563	 => std_logic_vector(to_unsigned(109,8) ,
14564	 => std_logic_vector(to_unsigned(96,8) ,
14565	 => std_logic_vector(to_unsigned(92,8) ,
14566	 => std_logic_vector(to_unsigned(93,8) ,
14567	 => std_logic_vector(to_unsigned(88,8) ,
14568	 => std_logic_vector(to_unsigned(99,8) ,
14569	 => std_logic_vector(to_unsigned(109,8) ,
14570	 => std_logic_vector(to_unsigned(61,8) ,
14571	 => std_logic_vector(to_unsigned(43,8) ,
14572	 => std_logic_vector(to_unsigned(56,8) ,
14573	 => std_logic_vector(to_unsigned(56,8) ,
14574	 => std_logic_vector(to_unsigned(70,8) ,
14575	 => std_logic_vector(to_unsigned(88,8) ,
14576	 => std_logic_vector(to_unsigned(90,8) ,
14577	 => std_logic_vector(to_unsigned(87,8) ,
14578	 => std_logic_vector(to_unsigned(93,8) ,
14579	 => std_logic_vector(to_unsigned(95,8) ,
14580	 => std_logic_vector(to_unsigned(86,8) ,
14581	 => std_logic_vector(to_unsigned(86,8) ,
14582	 => std_logic_vector(to_unsigned(96,8) ,
14583	 => std_logic_vector(to_unsigned(118,8) ,
14584	 => std_logic_vector(to_unsigned(107,8) ,
14585	 => std_logic_vector(to_unsigned(109,8) ,
14586	 => std_logic_vector(to_unsigned(95,8) ,
14587	 => std_logic_vector(to_unsigned(84,8) ,
14588	 => std_logic_vector(to_unsigned(109,8) ,
14589	 => std_logic_vector(to_unsigned(115,8) ,
14590	 => std_logic_vector(to_unsigned(115,8) ,
14591	 => std_logic_vector(to_unsigned(115,8) ,
14592	 => std_logic_vector(to_unsigned(108,8) ,
14593	 => std_logic_vector(to_unsigned(105,8) ,
14594	 => std_logic_vector(to_unsigned(99,8) ,
14595	 => std_logic_vector(to_unsigned(92,8) ,
14596	 => std_logic_vector(to_unsigned(93,8) ,
14597	 => std_logic_vector(to_unsigned(97,8) ,
14598	 => std_logic_vector(to_unsigned(95,8) ,
14599	 => std_logic_vector(to_unsigned(95,8) ,
14600	 => std_logic_vector(to_unsigned(96,8) ,
14601	 => std_logic_vector(to_unsigned(107,8) ,
14602	 => std_logic_vector(to_unsigned(109,8) ,
14603	 => std_logic_vector(to_unsigned(109,8) ,
14604	 => std_logic_vector(to_unsigned(93,8) ,
14605	 => std_logic_vector(to_unsigned(97,8) ,
14606	 => std_logic_vector(to_unsigned(100,8) ,
14607	 => std_logic_vector(to_unsigned(91,8) ,
14608	 => std_logic_vector(to_unsigned(104,8) ,
14609	 => std_logic_vector(to_unsigned(103,8) ,
14610	 => std_logic_vector(to_unsigned(73,8) ,
14611	 => std_logic_vector(to_unsigned(69,8) ,
14612	 => std_logic_vector(to_unsigned(85,8) ,
14613	 => std_logic_vector(to_unsigned(76,8) ,
14614	 => std_logic_vector(to_unsigned(54,8) ,
14615	 => std_logic_vector(to_unsigned(61,8) ,
14616	 => std_logic_vector(to_unsigned(81,8) ,
14617	 => std_logic_vector(to_unsigned(111,8) ,
14618	 => std_logic_vector(to_unsigned(111,8) ,
14619	 => std_logic_vector(to_unsigned(119,8) ,
14620	 => std_logic_vector(to_unsigned(114,8) ,
14621	 => std_logic_vector(to_unsigned(133,8) ,
14622	 => std_logic_vector(to_unsigned(115,8) ,
14623	 => std_logic_vector(to_unsigned(109,8) ,
14624	 => std_logic_vector(to_unsigned(100,8) ,
14625	 => std_logic_vector(to_unsigned(74,8) ,
14626	 => std_logic_vector(to_unsigned(70,8) ,
14627	 => std_logic_vector(to_unsigned(68,8) ,
14628	 => std_logic_vector(to_unsigned(71,8) ,
14629	 => std_logic_vector(to_unsigned(81,8) ,
14630	 => std_logic_vector(to_unsigned(91,8) ,
14631	 => std_logic_vector(to_unsigned(95,8) ,
14632	 => std_logic_vector(to_unsigned(81,8) ,
14633	 => std_logic_vector(to_unsigned(69,8) ,
14634	 => std_logic_vector(to_unsigned(67,8) ,
14635	 => std_logic_vector(to_unsigned(66,8) ,
14636	 => std_logic_vector(to_unsigned(61,8) ,
14637	 => std_logic_vector(to_unsigned(64,8) ,
14638	 => std_logic_vector(to_unsigned(66,8) ,
14639	 => std_logic_vector(to_unsigned(55,8) ,
14640	 => std_logic_vector(to_unsigned(54,8) ,
14641	 => std_logic_vector(to_unsigned(51,8) ,
14642	 => std_logic_vector(to_unsigned(51,8) ,
14643	 => std_logic_vector(to_unsigned(51,8) ,
14644	 => std_logic_vector(to_unsigned(46,8) ,
14645	 => std_logic_vector(to_unsigned(54,8) ,
14646	 => std_logic_vector(to_unsigned(22,8) ,
14647	 => std_logic_vector(to_unsigned(1,8) ,
14648	 => std_logic_vector(to_unsigned(0,8) ,
14649	 => std_logic_vector(to_unsigned(2,8) ,
14650	 => std_logic_vector(to_unsigned(46,8) ,
14651	 => std_logic_vector(to_unsigned(69,8) ,
14652	 => std_logic_vector(to_unsigned(54,8) ,
14653	 => std_logic_vector(to_unsigned(59,8) ,
14654	 => std_logic_vector(to_unsigned(57,8) ,
14655	 => std_logic_vector(to_unsigned(60,8) ,
14656	 => std_logic_vector(to_unsigned(68,8) ,
14657	 => std_logic_vector(to_unsigned(78,8) ,
14658	 => std_logic_vector(to_unsigned(82,8) ,
14659	 => std_logic_vector(to_unsigned(68,8) ,
14660	 => std_logic_vector(to_unsigned(71,8) ,
14661	 => std_logic_vector(to_unsigned(88,8) ,
14662	 => std_logic_vector(to_unsigned(86,8) ,
14663	 => std_logic_vector(to_unsigned(55,8) ,
14664	 => std_logic_vector(to_unsigned(64,8) ,
14665	 => std_logic_vector(to_unsigned(73,8) ,
14666	 => std_logic_vector(to_unsigned(69,8) ,
14667	 => std_logic_vector(to_unsigned(79,8) ,
14668	 => std_logic_vector(to_unsigned(74,8) ,
14669	 => std_logic_vector(to_unsigned(69,8) ,
14670	 => std_logic_vector(to_unsigned(85,8) ,
14671	 => std_logic_vector(to_unsigned(101,8) ,
14672	 => std_logic_vector(to_unsigned(90,8) ,
14673	 => std_logic_vector(to_unsigned(77,8) ,
14674	 => std_logic_vector(to_unsigned(56,8) ,
14675	 => std_logic_vector(to_unsigned(55,8) ,
14676	 => std_logic_vector(to_unsigned(66,8) ,
14677	 => std_logic_vector(to_unsigned(71,8) ,
14678	 => std_logic_vector(to_unsigned(68,8) ,
14679	 => std_logic_vector(to_unsigned(70,8) ,
14680	 => std_logic_vector(to_unsigned(70,8) ,
14681	 => std_logic_vector(to_unsigned(76,8) ,
14682	 => std_logic_vector(to_unsigned(80,8) ,
14683	 => std_logic_vector(to_unsigned(76,8) ,
14684	 => std_logic_vector(to_unsigned(70,8) ,
14685	 => std_logic_vector(to_unsigned(81,8) ,
14686	 => std_logic_vector(to_unsigned(91,8) ,
14687	 => std_logic_vector(to_unsigned(79,8) ,
14688	 => std_logic_vector(to_unsigned(84,8) ,
14689	 => std_logic_vector(to_unsigned(93,8) ,
14690	 => std_logic_vector(to_unsigned(99,8) ,
14691	 => std_logic_vector(to_unsigned(131,8) ,
14692	 => std_logic_vector(to_unsigned(103,8) ,
14693	 => std_logic_vector(to_unsigned(84,8) ,
14694	 => std_logic_vector(to_unsigned(95,8) ,
14695	 => std_logic_vector(to_unsigned(87,8) ,
14696	 => std_logic_vector(to_unsigned(114,8) ,
14697	 => std_logic_vector(to_unsigned(141,8) ,
14698	 => std_logic_vector(to_unsigned(154,8) ,
14699	 => std_logic_vector(to_unsigned(166,8) ,
14700	 => std_logic_vector(to_unsigned(164,8) ,
14701	 => std_logic_vector(to_unsigned(168,8) ,
14702	 => std_logic_vector(to_unsigned(163,8) ,
14703	 => std_logic_vector(to_unsigned(163,8) ,
14704	 => std_logic_vector(to_unsigned(159,8) ,
14705	 => std_logic_vector(to_unsigned(161,8) ,
14706	 => std_logic_vector(to_unsigned(161,8) ,
14707	 => std_logic_vector(to_unsigned(157,8) ,
14708	 => std_logic_vector(to_unsigned(163,8) ,
14709	 => std_logic_vector(to_unsigned(161,8) ,
14710	 => std_logic_vector(to_unsigned(164,8) ,
14711	 => std_logic_vector(to_unsigned(170,8) ,
14712	 => std_logic_vector(to_unsigned(159,8) ,
14713	 => std_logic_vector(to_unsigned(152,8) ,
14714	 => std_logic_vector(to_unsigned(168,8) ,
14715	 => std_logic_vector(to_unsigned(147,8) ,
14716	 => std_logic_vector(to_unsigned(154,8) ,
14717	 => std_logic_vector(to_unsigned(161,8) ,
14718	 => std_logic_vector(to_unsigned(163,8) ,
14719	 => std_logic_vector(to_unsigned(161,8) ,
14720	 => std_logic_vector(to_unsigned(154,8) ,
14721	 => std_logic_vector(to_unsigned(141,8) ,
14722	 => std_logic_vector(to_unsigned(142,8) ,
14723	 => std_logic_vector(to_unsigned(138,8) ,
14724	 => std_logic_vector(to_unsigned(127,8) ,
14725	 => std_logic_vector(to_unsigned(127,8) ,
14726	 => std_logic_vector(to_unsigned(151,8) ,
14727	 => std_logic_vector(to_unsigned(147,8) ,
14728	 => std_logic_vector(to_unsigned(142,8) ,
14729	 => std_logic_vector(to_unsigned(147,8) ,
14730	 => std_logic_vector(to_unsigned(146,8) ,
14731	 => std_logic_vector(to_unsigned(154,8) ,
14732	 => std_logic_vector(to_unsigned(144,8) ,
14733	 => std_logic_vector(to_unsigned(142,8) ,
14734	 => std_logic_vector(to_unsigned(142,8) ,
14735	 => std_logic_vector(to_unsigned(139,8) ,
14736	 => std_logic_vector(to_unsigned(149,8) ,
14737	 => std_logic_vector(to_unsigned(156,8) ,
14738	 => std_logic_vector(to_unsigned(146,8) ,
14739	 => std_logic_vector(to_unsigned(144,8) ,
14740	 => std_logic_vector(to_unsigned(159,8) ,
14741	 => std_logic_vector(to_unsigned(159,8) ,
14742	 => std_logic_vector(to_unsigned(152,8) ,
14743	 => std_logic_vector(to_unsigned(149,8) ,
14744	 => std_logic_vector(to_unsigned(157,8) ,
14745	 => std_logic_vector(to_unsigned(164,8) ,
14746	 => std_logic_vector(to_unsigned(149,8) ,
14747	 => std_logic_vector(to_unsigned(136,8) ,
14748	 => std_logic_vector(to_unsigned(133,8) ,
14749	 => std_logic_vector(to_unsigned(124,8) ,
14750	 => std_logic_vector(to_unsigned(131,8) ,
14751	 => std_logic_vector(to_unsigned(131,8) ,
14752	 => std_logic_vector(to_unsigned(134,8) ,
14753	 => std_logic_vector(to_unsigned(151,8) ,
14754	 => std_logic_vector(to_unsigned(142,8) ,
14755	 => std_logic_vector(to_unsigned(130,8) ,
14756	 => std_logic_vector(to_unsigned(141,8) ,
14757	 => std_logic_vector(to_unsigned(142,8) ,
14758	 => std_logic_vector(to_unsigned(144,8) ,
14759	 => std_logic_vector(to_unsigned(146,8) ,
14760	 => std_logic_vector(to_unsigned(139,8) ,
14761	 => std_logic_vector(to_unsigned(130,8) ,
14762	 => std_logic_vector(to_unsigned(134,8) ,
14763	 => std_logic_vector(to_unsigned(141,8) ,
14764	 => std_logic_vector(to_unsigned(131,8) ,
14765	 => std_logic_vector(to_unsigned(138,8) ,
14766	 => std_logic_vector(to_unsigned(138,8) ,
14767	 => std_logic_vector(to_unsigned(141,8) ,
14768	 => std_logic_vector(to_unsigned(142,8) ,
14769	 => std_logic_vector(to_unsigned(133,8) ,
14770	 => std_logic_vector(to_unsigned(136,8) ,
14771	 => std_logic_vector(to_unsigned(136,8) ,
14772	 => std_logic_vector(to_unsigned(147,8) ,
14773	 => std_logic_vector(to_unsigned(157,8) ,
14774	 => std_logic_vector(to_unsigned(156,8) ,
14775	 => std_logic_vector(to_unsigned(151,8) ,
14776	 => std_logic_vector(to_unsigned(147,8) ,
14777	 => std_logic_vector(to_unsigned(144,8) ,
14778	 => std_logic_vector(to_unsigned(149,8) ,
14779	 => std_logic_vector(to_unsigned(149,8) ,
14780	 => std_logic_vector(to_unsigned(152,8) ,
14781	 => std_logic_vector(to_unsigned(149,8) ,
14782	 => std_logic_vector(to_unsigned(149,8) ,
14783	 => std_logic_vector(to_unsigned(159,8) ,
14784	 => std_logic_vector(to_unsigned(157,8) ,
14785	 => std_logic_vector(to_unsigned(161,8) ,
14786	 => std_logic_vector(to_unsigned(156,8) ,
14787	 => std_logic_vector(to_unsigned(141,8) ,
14788	 => std_logic_vector(to_unsigned(138,8) ,
14789	 => std_logic_vector(to_unsigned(142,8) ,
14790	 => std_logic_vector(to_unsigned(133,8) ,
14791	 => std_logic_vector(to_unsigned(136,8) ,
14792	 => std_logic_vector(to_unsigned(138,8) ,
14793	 => std_logic_vector(to_unsigned(134,8) ,
14794	 => std_logic_vector(to_unsigned(121,8) ,
14795	 => std_logic_vector(to_unsigned(119,8) ,
14796	 => std_logic_vector(to_unsigned(119,8) ,
14797	 => std_logic_vector(to_unsigned(128,8) ,
14798	 => std_logic_vector(to_unsigned(121,8) ,
14799	 => std_logic_vector(to_unsigned(134,8) ,
14800	 => std_logic_vector(to_unsigned(146,8) ,
14801	 => std_logic_vector(to_unsigned(138,8) ,
14802	 => std_logic_vector(to_unsigned(133,8) ,
14803	 => std_logic_vector(to_unsigned(134,8) ,
14804	 => std_logic_vector(to_unsigned(122,8) ,
14805	 => std_logic_vector(to_unsigned(125,8) ,
14806	 => std_logic_vector(to_unsigned(144,8) ,
14807	 => std_logic_vector(to_unsigned(157,8) ,
14808	 => std_logic_vector(to_unsigned(161,8) ,
14809	 => std_logic_vector(to_unsigned(168,8) ,
14810	 => std_logic_vector(to_unsigned(168,8) ,
14811	 => std_logic_vector(to_unsigned(161,8) ,
14812	 => std_logic_vector(to_unsigned(156,8) ,
14813	 => std_logic_vector(to_unsigned(164,8) ,
14814	 => std_logic_vector(to_unsigned(171,8) ,
14815	 => std_logic_vector(to_unsigned(173,8) ,
14816	 => std_logic_vector(to_unsigned(173,8) ,
14817	 => std_logic_vector(to_unsigned(163,8) ,
14818	 => std_logic_vector(to_unsigned(154,8) ,
14819	 => std_logic_vector(to_unsigned(152,8) ,
14820	 => std_logic_vector(to_unsigned(151,8) ,
14821	 => std_logic_vector(to_unsigned(147,8) ,
14822	 => std_logic_vector(to_unsigned(156,8) ,
14823	 => std_logic_vector(to_unsigned(156,8) ,
14824	 => std_logic_vector(to_unsigned(156,8) ,
14825	 => std_logic_vector(to_unsigned(168,8) ,
14826	 => std_logic_vector(to_unsigned(141,8) ,
14827	 => std_logic_vector(to_unsigned(116,8) ,
14828	 => std_logic_vector(to_unsigned(118,8) ,
14829	 => std_logic_vector(to_unsigned(122,8) ,
14830	 => std_logic_vector(to_unsigned(130,8) ,
14831	 => std_logic_vector(to_unsigned(127,8) ,
14832	 => std_logic_vector(to_unsigned(111,8) ,
14833	 => std_logic_vector(to_unsigned(92,8) ,
14834	 => std_logic_vector(to_unsigned(93,8) ,
14835	 => std_logic_vector(to_unsigned(92,8) ,
14836	 => std_logic_vector(to_unsigned(93,8) ,
14837	 => std_logic_vector(to_unsigned(128,8) ,
14838	 => std_logic_vector(to_unsigned(121,8) ,
14839	 => std_logic_vector(to_unsigned(103,8) ,
14840	 => std_logic_vector(to_unsigned(121,8) ,
14841	 => std_logic_vector(to_unsigned(104,8) ,
14842	 => std_logic_vector(to_unsigned(112,8) ,
14843	 => std_logic_vector(to_unsigned(124,8) ,
14844	 => std_logic_vector(to_unsigned(103,8) ,
14845	 => std_logic_vector(to_unsigned(104,8) ,
14846	 => std_logic_vector(to_unsigned(107,8) ,
14847	 => std_logic_vector(to_unsigned(109,8) ,
14848	 => std_logic_vector(to_unsigned(111,8) ,
14849	 => std_logic_vector(to_unsigned(125,8) ,
14850	 => std_logic_vector(to_unsigned(139,8) ,
14851	 => std_logic_vector(to_unsigned(136,8) ,
14852	 => std_logic_vector(to_unsigned(141,8) ,
14853	 => std_logic_vector(to_unsigned(151,8) ,
14854	 => std_logic_vector(to_unsigned(124,8) ,
14855	 => std_logic_vector(to_unsigned(112,8) ,
14856	 => std_logic_vector(to_unsigned(115,8) ,
14857	 => std_logic_vector(to_unsigned(84,8) ,
14858	 => std_logic_vector(to_unsigned(103,8) ,
14859	 => std_logic_vector(to_unsigned(131,8) ,
14860	 => std_logic_vector(to_unsigned(122,8) ,
14861	 => std_logic_vector(to_unsigned(124,8) ,
14862	 => std_logic_vector(to_unsigned(125,8) ,
14863	 => std_logic_vector(to_unsigned(138,8) ,
14864	 => std_logic_vector(to_unsigned(136,8) ,
14865	 => std_logic_vector(to_unsigned(130,8) ,
14866	 => std_logic_vector(to_unsigned(114,8) ,
14867	 => std_logic_vector(to_unsigned(103,8) ,
14868	 => std_logic_vector(to_unsigned(81,8) ,
14869	 => std_logic_vector(to_unsigned(76,8) ,
14870	 => std_logic_vector(to_unsigned(77,8) ,
14871	 => std_logic_vector(to_unsigned(80,8) ,
14872	 => std_logic_vector(to_unsigned(95,8) ,
14873	 => std_logic_vector(to_unsigned(88,8) ,
14874	 => std_logic_vector(to_unsigned(82,8) ,
14875	 => std_logic_vector(to_unsigned(84,8) ,
14876	 => std_logic_vector(to_unsigned(84,8) ,
14877	 => std_logic_vector(to_unsigned(91,8) ,
14878	 => std_logic_vector(to_unsigned(112,8) ,
14879	 => std_logic_vector(to_unsigned(99,8) ,
14880	 => std_logic_vector(to_unsigned(57,8) ,
14881	 => std_logic_vector(to_unsigned(80,8) ,
14882	 => std_logic_vector(to_unsigned(104,8) ,
14883	 => std_logic_vector(to_unsigned(99,8) ,
14884	 => std_logic_vector(to_unsigned(96,8) ,
14885	 => std_logic_vector(to_unsigned(86,8) ,
14886	 => std_logic_vector(to_unsigned(90,8) ,
14887	 => std_logic_vector(to_unsigned(92,8) ,
14888	 => std_logic_vector(to_unsigned(96,8) ,
14889	 => std_logic_vector(to_unsigned(87,8) ,
14890	 => std_logic_vector(to_unsigned(54,8) ,
14891	 => std_logic_vector(to_unsigned(46,8) ,
14892	 => std_logic_vector(to_unsigned(61,8) ,
14893	 => std_logic_vector(to_unsigned(72,8) ,
14894	 => std_logic_vector(to_unsigned(74,8) ,
14895	 => std_logic_vector(to_unsigned(77,8) ,
14896	 => std_logic_vector(to_unsigned(86,8) ,
14897	 => std_logic_vector(to_unsigned(86,8) ,
14898	 => std_logic_vector(to_unsigned(88,8) ,
14899	 => std_logic_vector(to_unsigned(88,8) ,
14900	 => std_logic_vector(to_unsigned(86,8) ,
14901	 => std_logic_vector(to_unsigned(93,8) ,
14902	 => std_logic_vector(to_unsigned(99,8) ,
14903	 => std_logic_vector(to_unsigned(112,8) ,
14904	 => std_logic_vector(to_unsigned(105,8) ,
14905	 => std_logic_vector(to_unsigned(114,8) ,
14906	 => std_logic_vector(to_unsigned(111,8) ,
14907	 => std_logic_vector(to_unsigned(101,8) ,
14908	 => std_logic_vector(to_unsigned(107,8) ,
14909	 => std_logic_vector(to_unsigned(93,8) ,
14910	 => std_logic_vector(to_unsigned(101,8) ,
14911	 => std_logic_vector(to_unsigned(101,8) ,
14912	 => std_logic_vector(to_unsigned(99,8) ,
14913	 => std_logic_vector(to_unsigned(108,8) ,
14914	 => std_logic_vector(to_unsigned(91,8) ,
14915	 => std_logic_vector(to_unsigned(90,8) ,
14916	 => std_logic_vector(to_unsigned(100,8) ,
14917	 => std_logic_vector(to_unsigned(100,8) ,
14918	 => std_logic_vector(to_unsigned(108,8) ,
14919	 => std_logic_vector(to_unsigned(107,8) ,
14920	 => std_logic_vector(to_unsigned(107,8) ,
14921	 => std_logic_vector(to_unsigned(111,8) ,
14922	 => std_logic_vector(to_unsigned(112,8) ,
14923	 => std_logic_vector(to_unsigned(101,8) ,
14924	 => std_logic_vector(to_unsigned(91,8) ,
14925	 => std_logic_vector(to_unsigned(90,8) ,
14926	 => std_logic_vector(to_unsigned(92,8) ,
14927	 => std_logic_vector(to_unsigned(104,8) ,
14928	 => std_logic_vector(to_unsigned(111,8) ,
14929	 => std_logic_vector(to_unsigned(93,8) ,
14930	 => std_logic_vector(to_unsigned(91,8) ,
14931	 => std_logic_vector(to_unsigned(116,8) ,
14932	 => std_logic_vector(to_unsigned(131,8) ,
14933	 => std_logic_vector(to_unsigned(104,8) ,
14934	 => std_logic_vector(to_unsigned(51,8) ,
14935	 => std_logic_vector(to_unsigned(63,8) ,
14936	 => std_logic_vector(to_unsigned(86,8) ,
14937	 => std_logic_vector(to_unsigned(97,8) ,
14938	 => std_logic_vector(to_unsigned(103,8) ,
14939	 => std_logic_vector(to_unsigned(119,8) ,
14940	 => std_logic_vector(to_unsigned(86,8) ,
14941	 => std_logic_vector(to_unsigned(95,8) ,
14942	 => std_logic_vector(to_unsigned(112,8) ,
14943	 => std_logic_vector(to_unsigned(114,8) ,
14944	 => std_logic_vector(to_unsigned(107,8) ,
14945	 => std_logic_vector(to_unsigned(96,8) ,
14946	 => std_logic_vector(to_unsigned(92,8) ,
14947	 => std_logic_vector(to_unsigned(76,8) ,
14948	 => std_logic_vector(to_unsigned(71,8) ,
14949	 => std_logic_vector(to_unsigned(85,8) ,
14950	 => std_logic_vector(to_unsigned(85,8) ,
14951	 => std_logic_vector(to_unsigned(82,8) ,
14952	 => std_logic_vector(to_unsigned(76,8) ,
14953	 => std_logic_vector(to_unsigned(63,8) ,
14954	 => std_logic_vector(to_unsigned(66,8) ,
14955	 => std_logic_vector(to_unsigned(62,8) ,
14956	 => std_logic_vector(to_unsigned(63,8) ,
14957	 => std_logic_vector(to_unsigned(67,8) ,
14958	 => std_logic_vector(to_unsigned(66,8) ,
14959	 => std_logic_vector(to_unsigned(67,8) ,
14960	 => std_logic_vector(to_unsigned(60,8) ,
14961	 => std_logic_vector(to_unsigned(54,8) ,
14962	 => std_logic_vector(to_unsigned(56,8) ,
14963	 => std_logic_vector(to_unsigned(56,8) ,
14964	 => std_logic_vector(to_unsigned(56,8) ,
14965	 => std_logic_vector(to_unsigned(50,8) ,
14966	 => std_logic_vector(to_unsigned(39,8) ,
14967	 => std_logic_vector(to_unsigned(3,8) ,
14968	 => std_logic_vector(to_unsigned(0,8) ,
14969	 => std_logic_vector(to_unsigned(1,8) ,
14970	 => std_logic_vector(to_unsigned(27,8) ,
14971	 => std_logic_vector(to_unsigned(74,8) ,
14972	 => std_logic_vector(to_unsigned(60,8) ,
14973	 => std_logic_vector(to_unsigned(61,8) ,
14974	 => std_logic_vector(to_unsigned(62,8) ,
14975	 => std_logic_vector(to_unsigned(69,8) ,
14976	 => std_logic_vector(to_unsigned(70,8) ,
14977	 => std_logic_vector(to_unsigned(64,8) ,
14978	 => std_logic_vector(to_unsigned(65,8) ,
14979	 => std_logic_vector(to_unsigned(67,8) ,
14980	 => std_logic_vector(to_unsigned(63,8) ,
14981	 => std_logic_vector(to_unsigned(80,8) ,
14982	 => std_logic_vector(to_unsigned(81,8) ,
14983	 => std_logic_vector(to_unsigned(64,8) ,
14984	 => std_logic_vector(to_unsigned(63,8) ,
14985	 => std_logic_vector(to_unsigned(62,8) ,
14986	 => std_logic_vector(to_unsigned(70,8) ,
14987	 => std_logic_vector(to_unsigned(79,8) ,
14988	 => std_logic_vector(to_unsigned(65,8) ,
14989	 => std_logic_vector(to_unsigned(70,8) ,
14990	 => std_logic_vector(to_unsigned(81,8) ,
14991	 => std_logic_vector(to_unsigned(85,8) ,
14992	 => std_logic_vector(to_unsigned(74,8) ,
14993	 => std_logic_vector(to_unsigned(66,8) ,
14994	 => std_logic_vector(to_unsigned(62,8) ,
14995	 => std_logic_vector(to_unsigned(62,8) ,
14996	 => std_logic_vector(to_unsigned(62,8) ,
14997	 => std_logic_vector(to_unsigned(64,8) ,
14998	 => std_logic_vector(to_unsigned(68,8) ,
14999	 => std_logic_vector(to_unsigned(80,8) ,
15000	 => std_logic_vector(to_unsigned(72,8) ,
15001	 => std_logic_vector(to_unsigned(71,8) ,
15002	 => std_logic_vector(to_unsigned(68,8) ,
15003	 => std_logic_vector(to_unsigned(71,8) ,
15004	 => std_logic_vector(to_unsigned(76,8) ,
15005	 => std_logic_vector(to_unsigned(79,8) ,
15006	 => std_logic_vector(to_unsigned(76,8) ,
15007	 => std_logic_vector(to_unsigned(72,8) ,
15008	 => std_logic_vector(to_unsigned(80,8) ,
15009	 => std_logic_vector(to_unsigned(76,8) ,
15010	 => std_logic_vector(to_unsigned(81,8) ,
15011	 => std_logic_vector(to_unsigned(109,8) ,
15012	 => std_logic_vector(to_unsigned(93,8) ,
15013	 => std_logic_vector(to_unsigned(71,8) ,
15014	 => std_logic_vector(to_unsigned(74,8) ,
15015	 => std_logic_vector(to_unsigned(82,8) ,
15016	 => std_logic_vector(to_unsigned(80,8) ,
15017	 => std_logic_vector(to_unsigned(77,8) ,
15018	 => std_logic_vector(to_unsigned(112,8) ,
15019	 => std_logic_vector(to_unsigned(134,8) ,
15020	 => std_logic_vector(to_unsigned(133,8) ,
15021	 => std_logic_vector(to_unsigned(151,8) ,
15022	 => std_logic_vector(to_unsigned(157,8) ,
15023	 => std_logic_vector(to_unsigned(156,8) ,
15024	 => std_logic_vector(to_unsigned(159,8) ,
15025	 => std_logic_vector(to_unsigned(151,8) ,
15026	 => std_logic_vector(to_unsigned(163,8) ,
15027	 => std_logic_vector(to_unsigned(151,8) ,
15028	 => std_logic_vector(to_unsigned(131,8) ,
15029	 => std_logic_vector(to_unsigned(151,8) ,
15030	 => std_logic_vector(to_unsigned(147,8) ,
15031	 => std_logic_vector(to_unsigned(159,8) ,
15032	 => std_logic_vector(to_unsigned(139,8) ,
15033	 => std_logic_vector(to_unsigned(109,8) ,
15034	 => std_logic_vector(to_unsigned(124,8) ,
15035	 => std_logic_vector(to_unsigned(108,8) ,
15036	 => std_logic_vector(to_unsigned(131,8) ,
15037	 => std_logic_vector(to_unsigned(144,8) ,
15038	 => std_logic_vector(to_unsigned(144,8) ,
15039	 => std_logic_vector(to_unsigned(154,8) ,
15040	 => std_logic_vector(to_unsigned(139,8) ,
15041	 => std_logic_vector(to_unsigned(133,8) ,
15042	 => std_logic_vector(to_unsigned(141,8) ,
15043	 => std_logic_vector(to_unsigned(144,8) ,
15044	 => std_logic_vector(to_unsigned(130,8) ,
15045	 => std_logic_vector(to_unsigned(136,8) ,
15046	 => std_logic_vector(to_unsigned(149,8) ,
15047	 => std_logic_vector(to_unsigned(149,8) ,
15048	 => std_logic_vector(to_unsigned(146,8) ,
15049	 => std_logic_vector(to_unsigned(152,8) ,
15050	 => std_logic_vector(to_unsigned(156,8) ,
15051	 => std_logic_vector(to_unsigned(157,8) ,
15052	 => std_logic_vector(to_unsigned(156,8) ,
15053	 => std_logic_vector(to_unsigned(159,8) ,
15054	 => std_logic_vector(to_unsigned(154,8) ,
15055	 => std_logic_vector(to_unsigned(147,8) ,
15056	 => std_logic_vector(to_unsigned(151,8) ,
15057	 => std_logic_vector(to_unsigned(157,8) ,
15058	 => std_logic_vector(to_unsigned(157,8) ,
15059	 => std_logic_vector(to_unsigned(156,8) ,
15060	 => std_logic_vector(to_unsigned(161,8) ,
15061	 => std_logic_vector(to_unsigned(159,8) ,
15062	 => std_logic_vector(to_unsigned(156,8) ,
15063	 => std_logic_vector(to_unsigned(161,8) ,
15064	 => std_logic_vector(to_unsigned(161,8) ,
15065	 => std_logic_vector(to_unsigned(159,8) ,
15066	 => std_logic_vector(to_unsigned(154,8) ,
15067	 => std_logic_vector(to_unsigned(142,8) ,
15068	 => std_logic_vector(to_unsigned(138,8) ,
15069	 => std_logic_vector(to_unsigned(130,8) ,
15070	 => std_logic_vector(to_unsigned(134,8) ,
15071	 => std_logic_vector(to_unsigned(136,8) ,
15072	 => std_logic_vector(to_unsigned(136,8) ,
15073	 => std_logic_vector(to_unsigned(149,8) ,
15074	 => std_logic_vector(to_unsigned(142,8) ,
15075	 => std_logic_vector(to_unsigned(128,8) ,
15076	 => std_logic_vector(to_unsigned(139,8) ,
15077	 => std_logic_vector(to_unsigned(141,8) ,
15078	 => std_logic_vector(to_unsigned(142,8) ,
15079	 => std_logic_vector(to_unsigned(136,8) ,
15080	 => std_logic_vector(to_unsigned(134,8) ,
15081	 => std_logic_vector(to_unsigned(139,8) ,
15082	 => std_logic_vector(to_unsigned(139,8) ,
15083	 => std_logic_vector(to_unsigned(154,8) ,
15084	 => std_logic_vector(to_unsigned(146,8) ,
15085	 => std_logic_vector(to_unsigned(139,8) ,
15086	 => std_logic_vector(to_unsigned(131,8) ,
15087	 => std_logic_vector(to_unsigned(138,8) ,
15088	 => std_logic_vector(to_unsigned(141,8) ,
15089	 => std_logic_vector(to_unsigned(130,8) ,
15090	 => std_logic_vector(to_unsigned(133,8) ,
15091	 => std_logic_vector(to_unsigned(138,8) ,
15092	 => std_logic_vector(to_unsigned(146,8) ,
15093	 => std_logic_vector(to_unsigned(154,8) ,
15094	 => std_logic_vector(to_unsigned(157,8) ,
15095	 => std_logic_vector(to_unsigned(159,8) ,
15096	 => std_logic_vector(to_unsigned(159,8) ,
15097	 => std_logic_vector(to_unsigned(147,8) ,
15098	 => std_logic_vector(to_unsigned(139,8) ,
15099	 => std_logic_vector(to_unsigned(133,8) ,
15100	 => std_logic_vector(to_unsigned(141,8) ,
15101	 => std_logic_vector(to_unsigned(152,8) ,
15102	 => std_logic_vector(to_unsigned(152,8) ,
15103	 => std_logic_vector(to_unsigned(159,8) ,
15104	 => std_logic_vector(to_unsigned(152,8) ,
15105	 => std_logic_vector(to_unsigned(141,8) ,
15106	 => std_logic_vector(to_unsigned(138,8) ,
15107	 => std_logic_vector(to_unsigned(118,8) ,
15108	 => std_logic_vector(to_unsigned(125,8) ,
15109	 => std_logic_vector(to_unsigned(136,8) ,
15110	 => std_logic_vector(to_unsigned(125,8) ,
15111	 => std_logic_vector(to_unsigned(128,8) ,
15112	 => std_logic_vector(to_unsigned(131,8) ,
15113	 => std_logic_vector(to_unsigned(119,8) ,
15114	 => std_logic_vector(to_unsigned(108,8) ,
15115	 => std_logic_vector(to_unsigned(124,8) ,
15116	 => std_logic_vector(to_unsigned(128,8) ,
15117	 => std_logic_vector(to_unsigned(133,8) ,
15118	 => std_logic_vector(to_unsigned(121,8) ,
15119	 => std_logic_vector(to_unsigned(136,8) ,
15120	 => std_logic_vector(to_unsigned(152,8) ,
15121	 => std_logic_vector(to_unsigned(149,8) ,
15122	 => std_logic_vector(to_unsigned(138,8) ,
15123	 => std_logic_vector(to_unsigned(139,8) ,
15124	 => std_logic_vector(to_unsigned(138,8) ,
15125	 => std_logic_vector(to_unsigned(144,8) ,
15126	 => std_logic_vector(to_unsigned(159,8) ,
15127	 => std_logic_vector(to_unsigned(164,8) ,
15128	 => std_logic_vector(to_unsigned(166,8) ,
15129	 => std_logic_vector(to_unsigned(166,8) ,
15130	 => std_logic_vector(to_unsigned(168,8) ,
15131	 => std_logic_vector(to_unsigned(166,8) ,
15132	 => std_logic_vector(to_unsigned(159,8) ,
15133	 => std_logic_vector(to_unsigned(163,8) ,
15134	 => std_logic_vector(to_unsigned(171,8) ,
15135	 => std_logic_vector(to_unsigned(171,8) ,
15136	 => std_logic_vector(to_unsigned(170,8) ,
15137	 => std_logic_vector(to_unsigned(157,8) ,
15138	 => std_logic_vector(to_unsigned(156,8) ,
15139	 => std_logic_vector(to_unsigned(154,8) ,
15140	 => std_logic_vector(to_unsigned(154,8) ,
15141	 => std_logic_vector(to_unsigned(151,8) ,
15142	 => std_logic_vector(to_unsigned(157,8) ,
15143	 => std_logic_vector(to_unsigned(159,8) ,
15144	 => std_logic_vector(to_unsigned(152,8) ,
15145	 => std_logic_vector(to_unsigned(161,8) ,
15146	 => std_logic_vector(to_unsigned(144,8) ,
15147	 => std_logic_vector(to_unsigned(133,8) ,
15148	 => std_logic_vector(to_unsigned(138,8) ,
15149	 => std_logic_vector(to_unsigned(138,8) ,
15150	 => std_logic_vector(to_unsigned(128,8) ,
15151	 => std_logic_vector(to_unsigned(124,8) ,
15152	 => std_logic_vector(to_unsigned(124,8) ,
15153	 => std_logic_vector(to_unsigned(116,8) ,
15154	 => std_logic_vector(to_unsigned(119,8) ,
15155	 => std_logic_vector(to_unsigned(105,8) ,
15156	 => std_logic_vector(to_unsigned(92,8) ,
15157	 => std_logic_vector(to_unsigned(115,8) ,
15158	 => std_logic_vector(to_unsigned(131,8) ,
15159	 => std_logic_vector(to_unsigned(124,8) ,
15160	 => std_logic_vector(to_unsigned(116,8) ,
15161	 => std_logic_vector(to_unsigned(112,8) ,
15162	 => std_logic_vector(to_unsigned(128,8) ,
15163	 => std_logic_vector(to_unsigned(125,8) ,
15164	 => std_logic_vector(to_unsigned(112,8) ,
15165	 => std_logic_vector(to_unsigned(99,8) ,
15166	 => std_logic_vector(to_unsigned(108,8) ,
15167	 => std_logic_vector(to_unsigned(125,8) ,
15168	 => std_logic_vector(to_unsigned(121,8) ,
15169	 => std_logic_vector(to_unsigned(115,8) ,
15170	 => std_logic_vector(to_unsigned(125,8) ,
15171	 => std_logic_vector(to_unsigned(115,8) ,
15172	 => std_logic_vector(to_unsigned(112,8) ,
15173	 => std_logic_vector(to_unsigned(142,8) ,
15174	 => std_logic_vector(to_unsigned(122,8) ,
15175	 => std_logic_vector(to_unsigned(116,8) ,
15176	 => std_logic_vector(to_unsigned(131,8) ,
15177	 => std_logic_vector(to_unsigned(105,8) ,
15178	 => std_logic_vector(to_unsigned(101,8) ,
15179	 => std_logic_vector(to_unsigned(122,8) ,
15180	 => std_logic_vector(to_unsigned(109,8) ,
15181	 => std_logic_vector(to_unsigned(111,8) ,
15182	 => std_logic_vector(to_unsigned(114,8) ,
15183	 => std_logic_vector(to_unsigned(121,8) ,
15184	 => std_logic_vector(to_unsigned(107,8) ,
15185	 => std_logic_vector(to_unsigned(103,8) ,
15186	 => std_logic_vector(to_unsigned(68,8) ,
15187	 => std_logic_vector(to_unsigned(64,8) ,
15188	 => std_logic_vector(to_unsigned(71,8) ,
15189	 => std_logic_vector(to_unsigned(59,8) ,
15190	 => std_logic_vector(to_unsigned(66,8) ,
15191	 => std_logic_vector(to_unsigned(61,8) ,
15192	 => std_logic_vector(to_unsigned(82,8) ,
15193	 => std_logic_vector(to_unsigned(63,8) ,
15194	 => std_logic_vector(to_unsigned(73,8) ,
15195	 => std_logic_vector(to_unsigned(95,8) ,
15196	 => std_logic_vector(to_unsigned(99,8) ,
15197	 => std_logic_vector(to_unsigned(97,8) ,
15198	 => std_logic_vector(to_unsigned(101,8) ,
15199	 => std_logic_vector(to_unsigned(99,8) ,
15200	 => std_logic_vector(to_unsigned(62,8) ,
15201	 => std_logic_vector(to_unsigned(73,8) ,
15202	 => std_logic_vector(to_unsigned(99,8) ,
15203	 => std_logic_vector(to_unsigned(96,8) ,
15204	 => std_logic_vector(to_unsigned(88,8) ,
15205	 => std_logic_vector(to_unsigned(81,8) ,
15206	 => std_logic_vector(to_unsigned(86,8) ,
15207	 => std_logic_vector(to_unsigned(86,8) ,
15208	 => std_logic_vector(to_unsigned(87,8) ,
15209	 => std_logic_vector(to_unsigned(73,8) ,
15210	 => std_logic_vector(to_unsigned(67,8) ,
15211	 => std_logic_vector(to_unsigned(72,8) ,
15212	 => std_logic_vector(to_unsigned(80,8) ,
15213	 => std_logic_vector(to_unsigned(71,8) ,
15214	 => std_logic_vector(to_unsigned(66,8) ,
15215	 => std_logic_vector(to_unsigned(71,8) ,
15216	 => std_logic_vector(to_unsigned(84,8) ,
15217	 => std_logic_vector(to_unsigned(79,8) ,
15218	 => std_logic_vector(to_unsigned(85,8) ,
15219	 => std_logic_vector(to_unsigned(90,8) ,
15220	 => std_logic_vector(to_unsigned(90,8) ,
15221	 => std_logic_vector(to_unsigned(99,8) ,
15222	 => std_logic_vector(to_unsigned(103,8) ,
15223	 => std_logic_vector(to_unsigned(88,8) ,
15224	 => std_logic_vector(to_unsigned(82,8) ,
15225	 => std_logic_vector(to_unsigned(96,8) ,
15226	 => std_logic_vector(to_unsigned(100,8) ,
15227	 => std_logic_vector(to_unsigned(95,8) ,
15228	 => std_logic_vector(to_unsigned(107,8) ,
15229	 => std_logic_vector(to_unsigned(96,8) ,
15230	 => std_logic_vector(to_unsigned(86,8) ,
15231	 => std_logic_vector(to_unsigned(90,8) ,
15232	 => std_logic_vector(to_unsigned(95,8) ,
15233	 => std_logic_vector(to_unsigned(104,8) ,
15234	 => std_logic_vector(to_unsigned(109,8) ,
15235	 => std_logic_vector(to_unsigned(104,8) ,
15236	 => std_logic_vector(to_unsigned(107,8) ,
15237	 => std_logic_vector(to_unsigned(115,8) ,
15238	 => std_logic_vector(to_unsigned(119,8) ,
15239	 => std_logic_vector(to_unsigned(118,8) ,
15240	 => std_logic_vector(to_unsigned(118,8) ,
15241	 => std_logic_vector(to_unsigned(114,8) ,
15242	 => std_logic_vector(to_unsigned(112,8) ,
15243	 => std_logic_vector(to_unsigned(91,8) ,
15244	 => std_logic_vector(to_unsigned(88,8) ,
15245	 => std_logic_vector(to_unsigned(96,8) ,
15246	 => std_logic_vector(to_unsigned(107,8) ,
15247	 => std_logic_vector(to_unsigned(114,8) ,
15248	 => std_logic_vector(to_unsigned(115,8) ,
15249	 => std_logic_vector(to_unsigned(105,8) ,
15250	 => std_logic_vector(to_unsigned(73,8) ,
15251	 => std_logic_vector(to_unsigned(103,8) ,
15252	 => std_logic_vector(to_unsigned(108,8) ,
15253	 => std_logic_vector(to_unsigned(87,8) ,
15254	 => std_logic_vector(to_unsigned(59,8) ,
15255	 => std_logic_vector(to_unsigned(65,8) ,
15256	 => std_logic_vector(to_unsigned(72,8) ,
15257	 => std_logic_vector(to_unsigned(84,8) ,
15258	 => std_logic_vector(to_unsigned(108,8) ,
15259	 => std_logic_vector(to_unsigned(107,8) ,
15260	 => std_logic_vector(to_unsigned(100,8) ,
15261	 => std_logic_vector(to_unsigned(103,8) ,
15262	 => std_logic_vector(to_unsigned(109,8) ,
15263	 => std_logic_vector(to_unsigned(107,8) ,
15264	 => std_logic_vector(to_unsigned(97,8) ,
15265	 => std_logic_vector(to_unsigned(79,8) ,
15266	 => std_logic_vector(to_unsigned(65,8) ,
15267	 => std_logic_vector(to_unsigned(56,8) ,
15268	 => std_logic_vector(to_unsigned(55,8) ,
15269	 => std_logic_vector(to_unsigned(68,8) ,
15270	 => std_logic_vector(to_unsigned(81,8) ,
15271	 => std_logic_vector(to_unsigned(79,8) ,
15272	 => std_logic_vector(to_unsigned(68,8) ,
15273	 => std_logic_vector(to_unsigned(65,8) ,
15274	 => std_logic_vector(to_unsigned(68,8) ,
15275	 => std_logic_vector(to_unsigned(65,8) ,
15276	 => std_logic_vector(to_unsigned(51,8) ,
15277	 => std_logic_vector(to_unsigned(53,8) ,
15278	 => std_logic_vector(to_unsigned(60,8) ,
15279	 => std_logic_vector(to_unsigned(58,8) ,
15280	 => std_logic_vector(to_unsigned(54,8) ,
15281	 => std_logic_vector(to_unsigned(61,8) ,
15282	 => std_logic_vector(to_unsigned(59,8) ,
15283	 => std_logic_vector(to_unsigned(62,8) ,
15284	 => std_logic_vector(to_unsigned(62,8) ,
15285	 => std_logic_vector(to_unsigned(52,8) ,
15286	 => std_logic_vector(to_unsigned(54,8) ,
15287	 => std_logic_vector(to_unsigned(11,8) ,
15288	 => std_logic_vector(to_unsigned(0,8) ,
15289	 => std_logic_vector(to_unsigned(0,8) ,
15290	 => std_logic_vector(to_unsigned(12,8) ,
15291	 => std_logic_vector(to_unsigned(72,8) ,
15292	 => std_logic_vector(to_unsigned(72,8) ,
15293	 => std_logic_vector(to_unsigned(63,8) ,
15294	 => std_logic_vector(to_unsigned(69,8) ,
15295	 => std_logic_vector(to_unsigned(70,8) ,
15296	 => std_logic_vector(to_unsigned(63,8) ,
15297	 => std_logic_vector(to_unsigned(73,8) ,
15298	 => std_logic_vector(to_unsigned(64,8) ,
15299	 => std_logic_vector(to_unsigned(70,8) ,
15300	 => std_logic_vector(to_unsigned(77,8) ,
15301	 => std_logic_vector(to_unsigned(79,8) ,
15302	 => std_logic_vector(to_unsigned(78,8) ,
15303	 => std_logic_vector(to_unsigned(74,8) ,
15304	 => std_logic_vector(to_unsigned(64,8) ,
15305	 => std_logic_vector(to_unsigned(66,8) ,
15306	 => std_logic_vector(to_unsigned(70,8) ,
15307	 => std_logic_vector(to_unsigned(66,8) ,
15308	 => std_logic_vector(to_unsigned(68,8) ,
15309	 => std_logic_vector(to_unsigned(66,8) ,
15310	 => std_logic_vector(to_unsigned(71,8) ,
15311	 => std_logic_vector(to_unsigned(69,8) ,
15312	 => std_logic_vector(to_unsigned(62,8) ,
15313	 => std_logic_vector(to_unsigned(61,8) ,
15314	 => std_logic_vector(to_unsigned(69,8) ,
15315	 => std_logic_vector(to_unsigned(63,8) ,
15316	 => std_logic_vector(to_unsigned(66,8) ,
15317	 => std_logic_vector(to_unsigned(73,8) ,
15318	 => std_logic_vector(to_unsigned(64,8) ,
15319	 => std_logic_vector(to_unsigned(67,8) ,
15320	 => std_logic_vector(to_unsigned(69,8) ,
15321	 => std_logic_vector(to_unsigned(71,8) ,
15322	 => std_logic_vector(to_unsigned(69,8) ,
15323	 => std_logic_vector(to_unsigned(73,8) ,
15324	 => std_logic_vector(to_unsigned(72,8) ,
15325	 => std_logic_vector(to_unsigned(67,8) ,
15326	 => std_logic_vector(to_unsigned(67,8) ,
15327	 => std_logic_vector(to_unsigned(72,8) ,
15328	 => std_logic_vector(to_unsigned(73,8) ,
15329	 => std_logic_vector(to_unsigned(72,8) ,
15330	 => std_logic_vector(to_unsigned(80,8) ,
15331	 => std_logic_vector(to_unsigned(85,8) ,
15332	 => std_logic_vector(to_unsigned(86,8) ,
15333	 => std_logic_vector(to_unsigned(74,8) ,
15334	 => std_logic_vector(to_unsigned(69,8) ,
15335	 => std_logic_vector(to_unsigned(72,8) ,
15336	 => std_logic_vector(to_unsigned(72,8) ,
15337	 => std_logic_vector(to_unsigned(73,8) ,
15338	 => std_logic_vector(to_unsigned(79,8) ,
15339	 => std_logic_vector(to_unsigned(82,8) ,
15340	 => std_logic_vector(to_unsigned(86,8) ,
15341	 => std_logic_vector(to_unsigned(99,8) ,
15342	 => std_logic_vector(to_unsigned(100,8) ,
15343	 => std_logic_vector(to_unsigned(104,8) ,
15344	 => std_logic_vector(to_unsigned(121,8) ,
15345	 => std_logic_vector(to_unsigned(107,8) ,
15346	 => std_logic_vector(to_unsigned(118,8) ,
15347	 => std_logic_vector(to_unsigned(119,8) ,
15348	 => std_logic_vector(to_unsigned(93,8) ,
15349	 => std_logic_vector(to_unsigned(99,8) ,
15350	 => std_logic_vector(to_unsigned(104,8) ,
15351	 => std_logic_vector(to_unsigned(104,8) ,
15352	 => std_logic_vector(to_unsigned(109,8) ,
15353	 => std_logic_vector(to_unsigned(96,8) ,
15354	 => std_logic_vector(to_unsigned(88,8) ,
15355	 => std_logic_vector(to_unsigned(88,8) ,
15356	 => std_logic_vector(to_unsigned(105,8) ,
15357	 => std_logic_vector(to_unsigned(103,8) ,
15358	 => std_logic_vector(to_unsigned(109,8) ,
15359	 => std_logic_vector(to_unsigned(128,8) ,
15360	 => std_logic_vector(to_unsigned(111,8) ,
15361	 => std_logic_vector(to_unsigned(131,8) ,
15362	 => std_logic_vector(to_unsigned(139,8) ,
15363	 => std_logic_vector(to_unsigned(149,8) ,
15364	 => std_logic_vector(to_unsigned(146,8) ,
15365	 => std_logic_vector(to_unsigned(147,8) ,
15366	 => std_logic_vector(to_unsigned(151,8) ,
15367	 => std_logic_vector(to_unsigned(152,8) ,
15368	 => std_logic_vector(to_unsigned(146,8) ,
15369	 => std_logic_vector(to_unsigned(156,8) ,
15370	 => std_logic_vector(to_unsigned(159,8) ,
15371	 => std_logic_vector(to_unsigned(156,8) ,
15372	 => std_logic_vector(to_unsigned(154,8) ,
15373	 => std_logic_vector(to_unsigned(157,8) ,
15374	 => std_logic_vector(to_unsigned(151,8) ,
15375	 => std_logic_vector(to_unsigned(144,8) ,
15376	 => std_logic_vector(to_unsigned(146,8) ,
15377	 => std_logic_vector(to_unsigned(146,8) ,
15378	 => std_logic_vector(to_unsigned(144,8) ,
15379	 => std_logic_vector(to_unsigned(151,8) ,
15380	 => std_logic_vector(to_unsigned(159,8) ,
15381	 => std_logic_vector(to_unsigned(159,8) ,
15382	 => std_logic_vector(to_unsigned(157,8) ,
15383	 => std_logic_vector(to_unsigned(159,8) ,
15384	 => std_logic_vector(to_unsigned(159,8) ,
15385	 => std_logic_vector(to_unsigned(154,8) ,
15386	 => std_logic_vector(to_unsigned(147,8) ,
15387	 => std_logic_vector(to_unsigned(141,8) ,
15388	 => std_logic_vector(to_unsigned(136,8) ,
15389	 => std_logic_vector(to_unsigned(130,8) ,
15390	 => std_logic_vector(to_unsigned(130,8) ,
15391	 => std_logic_vector(to_unsigned(133,8) ,
15392	 => std_logic_vector(to_unsigned(139,8) ,
15393	 => std_logic_vector(to_unsigned(149,8) ,
15394	 => std_logic_vector(to_unsigned(142,8) ,
15395	 => std_logic_vector(to_unsigned(131,8) ,
15396	 => std_logic_vector(to_unsigned(138,8) ,
15397	 => std_logic_vector(to_unsigned(139,8) ,
15398	 => std_logic_vector(to_unsigned(138,8) ,
15399	 => std_logic_vector(to_unsigned(130,8) ,
15400	 => std_logic_vector(to_unsigned(131,8) ,
15401	 => std_logic_vector(to_unsigned(133,8) ,
15402	 => std_logic_vector(to_unsigned(125,8) ,
15403	 => std_logic_vector(to_unsigned(142,8) ,
15404	 => std_logic_vector(to_unsigned(144,8) ,
15405	 => std_logic_vector(to_unsigned(149,8) ,
15406	 => std_logic_vector(to_unsigned(146,8) ,
15407	 => std_logic_vector(to_unsigned(127,8) ,
15408	 => std_logic_vector(to_unsigned(122,8) ,
15409	 => std_logic_vector(to_unsigned(128,8) ,
15410	 => std_logic_vector(to_unsigned(133,8) ,
15411	 => std_logic_vector(to_unsigned(142,8) ,
15412	 => std_logic_vector(to_unsigned(149,8) ,
15413	 => std_logic_vector(to_unsigned(154,8) ,
15414	 => std_logic_vector(to_unsigned(157,8) ,
15415	 => std_logic_vector(to_unsigned(159,8) ,
15416	 => std_logic_vector(to_unsigned(159,8) ,
15417	 => std_logic_vector(to_unsigned(146,8) ,
15418	 => std_logic_vector(to_unsigned(131,8) ,
15419	 => std_logic_vector(to_unsigned(125,8) ,
15420	 => std_logic_vector(to_unsigned(125,8) ,
15421	 => std_logic_vector(to_unsigned(141,8) ,
15422	 => std_logic_vector(to_unsigned(154,8) ,
15423	 => std_logic_vector(to_unsigned(161,8) ,
15424	 => std_logic_vector(to_unsigned(146,8) ,
15425	 => std_logic_vector(to_unsigned(119,8) ,
15426	 => std_logic_vector(to_unsigned(122,8) ,
15427	 => std_logic_vector(to_unsigned(116,8) ,
15428	 => std_logic_vector(to_unsigned(118,8) ,
15429	 => std_logic_vector(to_unsigned(119,8) ,
15430	 => std_logic_vector(to_unsigned(115,8) ,
15431	 => std_logic_vector(to_unsigned(104,8) ,
15432	 => std_logic_vector(to_unsigned(114,8) ,
15433	 => std_logic_vector(to_unsigned(131,8) ,
15434	 => std_logic_vector(to_unsigned(127,8) ,
15435	 => std_logic_vector(to_unsigned(124,8) ,
15436	 => std_logic_vector(to_unsigned(127,8) ,
15437	 => std_logic_vector(to_unsigned(136,8) ,
15438	 => std_logic_vector(to_unsigned(125,8) ,
15439	 => std_logic_vector(to_unsigned(142,8) ,
15440	 => std_logic_vector(to_unsigned(157,8) ,
15441	 => std_logic_vector(to_unsigned(151,8) ,
15442	 => std_logic_vector(to_unsigned(139,8) ,
15443	 => std_logic_vector(to_unsigned(142,8) ,
15444	 => std_logic_vector(to_unsigned(146,8) ,
15445	 => std_logic_vector(to_unsigned(159,8) ,
15446	 => std_logic_vector(to_unsigned(161,8) ,
15447	 => std_logic_vector(to_unsigned(163,8) ,
15448	 => std_logic_vector(to_unsigned(164,8) ,
15449	 => std_logic_vector(to_unsigned(163,8) ,
15450	 => std_logic_vector(to_unsigned(163,8) ,
15451	 => std_logic_vector(to_unsigned(166,8) ,
15452	 => std_logic_vector(to_unsigned(166,8) ,
15453	 => std_logic_vector(to_unsigned(170,8) ,
15454	 => std_logic_vector(to_unsigned(173,8) ,
15455	 => std_logic_vector(to_unsigned(171,8) ,
15456	 => std_logic_vector(to_unsigned(168,8) ,
15457	 => std_logic_vector(to_unsigned(154,8) ,
15458	 => std_logic_vector(to_unsigned(156,8) ,
15459	 => std_logic_vector(to_unsigned(156,8) ,
15460	 => std_logic_vector(to_unsigned(157,8) ,
15461	 => std_logic_vector(to_unsigned(161,8) ,
15462	 => std_logic_vector(to_unsigned(159,8) ,
15463	 => std_logic_vector(to_unsigned(156,8) ,
15464	 => std_logic_vector(to_unsigned(151,8) ,
15465	 => std_logic_vector(to_unsigned(154,8) ,
15466	 => std_logic_vector(to_unsigned(149,8) ,
15467	 => std_logic_vector(to_unsigned(142,8) ,
15468	 => std_logic_vector(to_unsigned(142,8) ,
15469	 => std_logic_vector(to_unsigned(161,8) ,
15470	 => std_logic_vector(to_unsigned(159,8) ,
15471	 => std_logic_vector(to_unsigned(139,8) ,
15472	 => std_logic_vector(to_unsigned(136,8) ,
15473	 => std_logic_vector(to_unsigned(131,8) ,
15474	 => std_logic_vector(to_unsigned(130,8) ,
15475	 => std_logic_vector(to_unsigned(108,8) ,
15476	 => std_logic_vector(to_unsigned(92,8) ,
15477	 => std_logic_vector(to_unsigned(95,8) ,
15478	 => std_logic_vector(to_unsigned(122,8) ,
15479	 => std_logic_vector(to_unsigned(128,8) ,
15480	 => std_logic_vector(to_unsigned(114,8) ,
15481	 => std_logic_vector(to_unsigned(124,8) ,
15482	 => std_logic_vector(to_unsigned(139,8) ,
15483	 => std_logic_vector(to_unsigned(139,8) ,
15484	 => std_logic_vector(to_unsigned(128,8) ,
15485	 => std_logic_vector(to_unsigned(86,8) ,
15486	 => std_logic_vector(to_unsigned(87,8) ,
15487	 => std_logic_vector(to_unsigned(115,8) ,
15488	 => std_logic_vector(to_unsigned(121,8) ,
15489	 => std_logic_vector(to_unsigned(108,8) ,
15490	 => std_logic_vector(to_unsigned(99,8) ,
15491	 => std_logic_vector(to_unsigned(100,8) ,
15492	 => std_logic_vector(to_unsigned(99,8) ,
15493	 => std_logic_vector(to_unsigned(119,8) ,
15494	 => std_logic_vector(to_unsigned(112,8) ,
15495	 => std_logic_vector(to_unsigned(109,8) ,
15496	 => std_logic_vector(to_unsigned(115,8) ,
15497	 => std_logic_vector(to_unsigned(118,8) ,
15498	 => std_logic_vector(to_unsigned(104,8) ,
15499	 => std_logic_vector(to_unsigned(111,8) ,
15500	 => std_logic_vector(to_unsigned(103,8) ,
15501	 => std_logic_vector(to_unsigned(103,8) ,
15502	 => std_logic_vector(to_unsigned(109,8) ,
15503	 => std_logic_vector(to_unsigned(116,8) ,
15504	 => std_logic_vector(to_unsigned(101,8) ,
15505	 => std_logic_vector(to_unsigned(93,8) ,
15506	 => std_logic_vector(to_unsigned(76,8) ,
15507	 => std_logic_vector(to_unsigned(67,8) ,
15508	 => std_logic_vector(to_unsigned(66,8) ,
15509	 => std_logic_vector(to_unsigned(62,8) ,
15510	 => std_logic_vector(to_unsigned(59,8) ,
15511	 => std_logic_vector(to_unsigned(58,8) ,
15512	 => std_logic_vector(to_unsigned(91,8) ,
15513	 => std_logic_vector(to_unsigned(67,8) ,
15514	 => std_logic_vector(to_unsigned(72,8) ,
15515	 => std_logic_vector(to_unsigned(104,8) ,
15516	 => std_logic_vector(to_unsigned(103,8) ,
15517	 => std_logic_vector(to_unsigned(86,8) ,
15518	 => std_logic_vector(to_unsigned(87,8) ,
15519	 => std_logic_vector(to_unsigned(87,8) ,
15520	 => std_logic_vector(to_unsigned(74,8) ,
15521	 => std_logic_vector(to_unsigned(70,8) ,
15522	 => std_logic_vector(to_unsigned(93,8) ,
15523	 => std_logic_vector(to_unsigned(97,8) ,
15524	 => std_logic_vector(to_unsigned(92,8) ,
15525	 => std_logic_vector(to_unsigned(92,8) ,
15526	 => std_logic_vector(to_unsigned(91,8) ,
15527	 => std_logic_vector(to_unsigned(86,8) ,
15528	 => std_logic_vector(to_unsigned(87,8) ,
15529	 => std_logic_vector(to_unsigned(85,8) ,
15530	 => std_logic_vector(to_unsigned(88,8) ,
15531	 => std_logic_vector(to_unsigned(85,8) ,
15532	 => std_logic_vector(to_unsigned(76,8) ,
15533	 => std_logic_vector(to_unsigned(73,8) ,
15534	 => std_logic_vector(to_unsigned(69,8) ,
15535	 => std_logic_vector(to_unsigned(78,8) ,
15536	 => std_logic_vector(to_unsigned(85,8) ,
15537	 => std_logic_vector(to_unsigned(71,8) ,
15538	 => std_logic_vector(to_unsigned(80,8) ,
15539	 => std_logic_vector(to_unsigned(100,8) ,
15540	 => std_logic_vector(to_unsigned(107,8) ,
15541	 => std_logic_vector(to_unsigned(109,8) ,
15542	 => std_logic_vector(to_unsigned(107,8) ,
15543	 => std_logic_vector(to_unsigned(88,8) ,
15544	 => std_logic_vector(to_unsigned(88,8) ,
15545	 => std_logic_vector(to_unsigned(92,8) ,
15546	 => std_logic_vector(to_unsigned(84,8) ,
15547	 => std_logic_vector(to_unsigned(80,8) ,
15548	 => std_logic_vector(to_unsigned(97,8) ,
15549	 => std_logic_vector(to_unsigned(104,8) ,
15550	 => std_logic_vector(to_unsigned(87,8) ,
15551	 => std_logic_vector(to_unsigned(97,8) ,
15552	 => std_logic_vector(to_unsigned(109,8) ,
15553	 => std_logic_vector(to_unsigned(108,8) ,
15554	 => std_logic_vector(to_unsigned(130,8) ,
15555	 => std_logic_vector(to_unsigned(109,8) ,
15556	 => std_logic_vector(to_unsigned(105,8) ,
15557	 => std_logic_vector(to_unsigned(131,8) ,
15558	 => std_logic_vector(to_unsigned(119,8) ,
15559	 => std_logic_vector(to_unsigned(114,8) ,
15560	 => std_logic_vector(to_unsigned(125,8) ,
15561	 => std_logic_vector(to_unsigned(124,8) ,
15562	 => std_logic_vector(to_unsigned(108,8) ,
15563	 => std_logic_vector(to_unsigned(100,8) ,
15564	 => std_logic_vector(to_unsigned(92,8) ,
15565	 => std_logic_vector(to_unsigned(93,8) ,
15566	 => std_logic_vector(to_unsigned(100,8) ,
15567	 => std_logic_vector(to_unsigned(108,8) ,
15568	 => std_logic_vector(to_unsigned(119,8) ,
15569	 => std_logic_vector(to_unsigned(114,8) ,
15570	 => std_logic_vector(to_unsigned(68,8) ,
15571	 => std_logic_vector(to_unsigned(81,8) ,
15572	 => std_logic_vector(to_unsigned(104,8) ,
15573	 => std_logic_vector(to_unsigned(97,8) ,
15574	 => std_logic_vector(to_unsigned(69,8) ,
15575	 => std_logic_vector(to_unsigned(69,8) ,
15576	 => std_logic_vector(to_unsigned(66,8) ,
15577	 => std_logic_vector(to_unsigned(71,8) ,
15578	 => std_logic_vector(to_unsigned(92,8) ,
15579	 => std_logic_vector(to_unsigned(85,8) ,
15580	 => std_logic_vector(to_unsigned(93,8) ,
15581	 => std_logic_vector(to_unsigned(116,8) ,
15582	 => std_logic_vector(to_unsigned(90,8) ,
15583	 => std_logic_vector(to_unsigned(76,8) ,
15584	 => std_logic_vector(to_unsigned(64,8) ,
15585	 => std_logic_vector(to_unsigned(73,8) ,
15586	 => std_logic_vector(to_unsigned(65,8) ,
15587	 => std_logic_vector(to_unsigned(56,8) ,
15588	 => std_logic_vector(to_unsigned(67,8) ,
15589	 => std_logic_vector(to_unsigned(65,8) ,
15590	 => std_logic_vector(to_unsigned(67,8) ,
15591	 => std_logic_vector(to_unsigned(74,8) ,
15592	 => std_logic_vector(to_unsigned(73,8) ,
15593	 => std_logic_vector(to_unsigned(66,8) ,
15594	 => std_logic_vector(to_unsigned(67,8) ,
15595	 => std_logic_vector(to_unsigned(67,8) ,
15596	 => std_logic_vector(to_unsigned(56,8) ,
15597	 => std_logic_vector(to_unsigned(57,8) ,
15598	 => std_logic_vector(to_unsigned(63,8) ,
15599	 => std_logic_vector(to_unsigned(63,8) ,
15600	 => std_logic_vector(to_unsigned(64,8) ,
15601	 => std_logic_vector(to_unsigned(61,8) ,
15602	 => std_logic_vector(to_unsigned(55,8) ,
15603	 => std_logic_vector(to_unsigned(61,8) ,
15604	 => std_logic_vector(to_unsigned(60,8) ,
15605	 => std_logic_vector(to_unsigned(57,8) ,
15606	 => std_logic_vector(to_unsigned(60,8) ,
15607	 => std_logic_vector(to_unsigned(18,8) ,
15608	 => std_logic_vector(to_unsigned(0,8) ,
15609	 => std_logic_vector(to_unsigned(0,8) ,
15610	 => std_logic_vector(to_unsigned(5,8) ,
15611	 => std_logic_vector(to_unsigned(62,8) ,
15612	 => std_logic_vector(to_unsigned(69,8) ,
15613	 => std_logic_vector(to_unsigned(60,8) ,
15614	 => std_logic_vector(to_unsigned(73,8) ,
15615	 => std_logic_vector(to_unsigned(87,8) ,
15616	 => std_logic_vector(to_unsigned(74,8) ,
15617	 => std_logic_vector(to_unsigned(86,8) ,
15618	 => std_logic_vector(to_unsigned(80,8) ,
15619	 => std_logic_vector(to_unsigned(74,8) ,
15620	 => std_logic_vector(to_unsigned(79,8) ,
15621	 => std_logic_vector(to_unsigned(77,8) ,
15622	 => std_logic_vector(to_unsigned(74,8) ,
15623	 => std_logic_vector(to_unsigned(66,8) ,
15624	 => std_logic_vector(to_unsigned(70,8) ,
15625	 => std_logic_vector(to_unsigned(81,8) ,
15626	 => std_logic_vector(to_unsigned(73,8) ,
15627	 => std_logic_vector(to_unsigned(69,8) ,
15628	 => std_logic_vector(to_unsigned(77,8) ,
15629	 => std_logic_vector(to_unsigned(72,8) ,
15630	 => std_logic_vector(to_unsigned(68,8) ,
15631	 => std_logic_vector(to_unsigned(67,8) ,
15632	 => std_logic_vector(to_unsigned(62,8) ,
15633	 => std_logic_vector(to_unsigned(62,8) ,
15634	 => std_logic_vector(to_unsigned(64,8) ,
15635	 => std_logic_vector(to_unsigned(51,8) ,
15636	 => std_logic_vector(to_unsigned(59,8) ,
15637	 => std_logic_vector(to_unsigned(71,8) ,
15638	 => std_logic_vector(to_unsigned(57,8) ,
15639	 => std_logic_vector(to_unsigned(57,8) ,
15640	 => std_logic_vector(to_unsigned(68,8) ,
15641	 => std_logic_vector(to_unsigned(73,8) ,
15642	 => std_logic_vector(to_unsigned(68,8) ,
15643	 => std_logic_vector(to_unsigned(70,8) ,
15644	 => std_logic_vector(to_unsigned(76,8) ,
15645	 => std_logic_vector(to_unsigned(70,8) ,
15646	 => std_logic_vector(to_unsigned(73,8) ,
15647	 => std_logic_vector(to_unsigned(74,8) ,
15648	 => std_logic_vector(to_unsigned(66,8) ,
15649	 => std_logic_vector(to_unsigned(77,8) ,
15650	 => std_logic_vector(to_unsigned(77,8) ,
15651	 => std_logic_vector(to_unsigned(77,8) ,
15652	 => std_logic_vector(to_unsigned(79,8) ,
15653	 => std_logic_vector(to_unsigned(72,8) ,
15654	 => std_logic_vector(to_unsigned(71,8) ,
15655	 => std_logic_vector(to_unsigned(74,8) ,
15656	 => std_logic_vector(to_unsigned(76,8) ,
15657	 => std_logic_vector(to_unsigned(90,8) ,
15658	 => std_logic_vector(to_unsigned(81,8) ,
15659	 => std_logic_vector(to_unsigned(80,8) ,
15660	 => std_logic_vector(to_unsigned(80,8) ,
15661	 => std_logic_vector(to_unsigned(86,8) ,
15662	 => std_logic_vector(to_unsigned(81,8) ,
15663	 => std_logic_vector(to_unsigned(85,8) ,
15664	 => std_logic_vector(to_unsigned(99,8) ,
15665	 => std_logic_vector(to_unsigned(91,8) ,
15666	 => std_logic_vector(to_unsigned(87,8) ,
15667	 => std_logic_vector(to_unsigned(93,8) ,
15668	 => std_logic_vector(to_unsigned(87,8) ,
15669	 => std_logic_vector(to_unsigned(79,8) ,
15670	 => std_logic_vector(to_unsigned(95,8) ,
15671	 => std_logic_vector(to_unsigned(95,8) ,
15672	 => std_logic_vector(to_unsigned(96,8) ,
15673	 => std_logic_vector(to_unsigned(91,8) ,
15674	 => std_logic_vector(to_unsigned(86,8) ,
15675	 => std_logic_vector(to_unsigned(80,8) ,
15676	 => std_logic_vector(to_unsigned(86,8) ,
15677	 => std_logic_vector(to_unsigned(96,8) ,
15678	 => std_logic_vector(to_unsigned(100,8) ,
15679	 => std_logic_vector(to_unsigned(101,8) ,
15680	 => std_logic_vector(to_unsigned(97,8) ,
15681	 => std_logic_vector(to_unsigned(139,8) ,
15682	 => std_logic_vector(to_unsigned(142,8) ,
15683	 => std_logic_vector(to_unsigned(146,8) ,
15684	 => std_logic_vector(to_unsigned(157,8) ,
15685	 => std_logic_vector(to_unsigned(152,8) ,
15686	 => std_logic_vector(to_unsigned(149,8) ,
15687	 => std_logic_vector(to_unsigned(152,8) ,
15688	 => std_logic_vector(to_unsigned(149,8) ,
15689	 => std_logic_vector(to_unsigned(157,8) ,
15690	 => std_logic_vector(to_unsigned(163,8) ,
15691	 => std_logic_vector(to_unsigned(157,8) ,
15692	 => std_logic_vector(to_unsigned(156,8) ,
15693	 => std_logic_vector(to_unsigned(154,8) ,
15694	 => std_logic_vector(to_unsigned(151,8) ,
15695	 => std_logic_vector(to_unsigned(147,8) ,
15696	 => std_logic_vector(to_unsigned(151,8) ,
15697	 => std_logic_vector(to_unsigned(149,8) ,
15698	 => std_logic_vector(to_unsigned(151,8) ,
15699	 => std_logic_vector(to_unsigned(156,8) ,
15700	 => std_logic_vector(to_unsigned(157,8) ,
15701	 => std_logic_vector(to_unsigned(156,8) ,
15702	 => std_logic_vector(to_unsigned(157,8) ,
15703	 => std_logic_vector(to_unsigned(156,8) ,
15704	 => std_logic_vector(to_unsigned(159,8) ,
15705	 => std_logic_vector(to_unsigned(156,8) ,
15706	 => std_logic_vector(to_unsigned(147,8) ,
15707	 => std_logic_vector(to_unsigned(146,8) ,
15708	 => std_logic_vector(to_unsigned(142,8) ,
15709	 => std_logic_vector(to_unsigned(138,8) ,
15710	 => std_logic_vector(to_unsigned(138,8) ,
15711	 => std_logic_vector(to_unsigned(146,8) ,
15712	 => std_logic_vector(to_unsigned(149,8) ,
15713	 => std_logic_vector(to_unsigned(151,8) ,
15714	 => std_logic_vector(to_unsigned(149,8) ,
15715	 => std_logic_vector(to_unsigned(134,8) ,
15716	 => std_logic_vector(to_unsigned(134,8) ,
15717	 => std_logic_vector(to_unsigned(142,8) ,
15718	 => std_logic_vector(to_unsigned(139,8) ,
15719	 => std_logic_vector(to_unsigned(131,8) ,
15720	 => std_logic_vector(to_unsigned(134,8) ,
15721	 => std_logic_vector(to_unsigned(131,8) ,
15722	 => std_logic_vector(to_unsigned(127,8) ,
15723	 => std_logic_vector(to_unsigned(131,8) ,
15724	 => std_logic_vector(to_unsigned(141,8) ,
15725	 => std_logic_vector(to_unsigned(157,8) ,
15726	 => std_logic_vector(to_unsigned(159,8) ,
15727	 => std_logic_vector(to_unsigned(141,8) ,
15728	 => std_logic_vector(to_unsigned(127,8) ,
15729	 => std_logic_vector(to_unsigned(133,8) ,
15730	 => std_logic_vector(to_unsigned(149,8) ,
15731	 => std_logic_vector(to_unsigned(156,8) ,
15732	 => std_logic_vector(to_unsigned(157,8) ,
15733	 => std_logic_vector(to_unsigned(152,8) ,
15734	 => std_logic_vector(to_unsigned(147,8) ,
15735	 => std_logic_vector(to_unsigned(138,8) ,
15736	 => std_logic_vector(to_unsigned(131,8) ,
15737	 => std_logic_vector(to_unsigned(133,8) ,
15738	 => std_logic_vector(to_unsigned(138,8) ,
15739	 => std_logic_vector(to_unsigned(133,8) ,
15740	 => std_logic_vector(to_unsigned(119,8) ,
15741	 => std_logic_vector(to_unsigned(127,8) ,
15742	 => std_logic_vector(to_unsigned(144,8) ,
15743	 => std_logic_vector(to_unsigned(157,8) ,
15744	 => std_logic_vector(to_unsigned(149,8) ,
15745	 => std_logic_vector(to_unsigned(133,8) ,
15746	 => std_logic_vector(to_unsigned(131,8) ,
15747	 => std_logic_vector(to_unsigned(133,8) ,
15748	 => std_logic_vector(to_unsigned(128,8) ,
15749	 => std_logic_vector(to_unsigned(118,8) ,
15750	 => std_logic_vector(to_unsigned(128,8) ,
15751	 => std_logic_vector(to_unsigned(128,8) ,
15752	 => std_logic_vector(to_unsigned(124,8) ,
15753	 => std_logic_vector(to_unsigned(142,8) ,
15754	 => std_logic_vector(to_unsigned(159,8) ,
15755	 => std_logic_vector(to_unsigned(152,8) ,
15756	 => std_logic_vector(to_unsigned(144,8) ,
15757	 => std_logic_vector(to_unsigned(144,8) ,
15758	 => std_logic_vector(to_unsigned(136,8) ,
15759	 => std_logic_vector(to_unsigned(139,8) ,
15760	 => std_logic_vector(to_unsigned(144,8) ,
15761	 => std_logic_vector(to_unsigned(147,8) ,
15762	 => std_logic_vector(to_unsigned(154,8) ,
15763	 => std_logic_vector(to_unsigned(154,8) ,
15764	 => std_logic_vector(to_unsigned(152,8) ,
15765	 => std_logic_vector(to_unsigned(157,8) ,
15766	 => std_logic_vector(to_unsigned(159,8) ,
15767	 => std_logic_vector(to_unsigned(161,8) ,
15768	 => std_logic_vector(to_unsigned(163,8) ,
15769	 => std_logic_vector(to_unsigned(161,8) ,
15770	 => std_logic_vector(to_unsigned(164,8) ,
15771	 => std_logic_vector(to_unsigned(161,8) ,
15772	 => std_logic_vector(to_unsigned(163,8) ,
15773	 => std_logic_vector(to_unsigned(166,8) ,
15774	 => std_logic_vector(to_unsigned(170,8) ,
15775	 => std_logic_vector(to_unsigned(173,8) ,
15776	 => std_logic_vector(to_unsigned(171,8) ,
15777	 => std_logic_vector(to_unsigned(152,8) ,
15778	 => std_logic_vector(to_unsigned(151,8) ,
15779	 => std_logic_vector(to_unsigned(159,8) ,
15780	 => std_logic_vector(to_unsigned(156,8) ,
15781	 => std_logic_vector(to_unsigned(157,8) ,
15782	 => std_logic_vector(to_unsigned(159,8) ,
15783	 => std_logic_vector(to_unsigned(154,8) ,
15784	 => std_logic_vector(to_unsigned(151,8) ,
15785	 => std_logic_vector(to_unsigned(151,8) ,
15786	 => std_logic_vector(to_unsigned(151,8) ,
15787	 => std_logic_vector(to_unsigned(151,8) ,
15788	 => std_logic_vector(to_unsigned(151,8) ,
15789	 => std_logic_vector(to_unsigned(156,8) ,
15790	 => std_logic_vector(to_unsigned(164,8) ,
15791	 => std_logic_vector(to_unsigned(151,8) ,
15792	 => std_logic_vector(to_unsigned(139,8) ,
15793	 => std_logic_vector(to_unsigned(125,8) ,
15794	 => std_logic_vector(to_unsigned(131,8) ,
15795	 => std_logic_vector(to_unsigned(109,8) ,
15796	 => std_logic_vector(to_unsigned(114,8) ,
15797	 => std_logic_vector(to_unsigned(104,8) ,
15798	 => std_logic_vector(to_unsigned(121,8) ,
15799	 => std_logic_vector(to_unsigned(127,8) ,
15800	 => std_logic_vector(to_unsigned(107,8) ,
15801	 => std_logic_vector(to_unsigned(133,8) ,
15802	 => std_logic_vector(to_unsigned(146,8) ,
15803	 => std_logic_vector(to_unsigned(146,8) ,
15804	 => std_logic_vector(to_unsigned(136,8) ,
15805	 => std_logic_vector(to_unsigned(97,8) ,
15806	 => std_logic_vector(to_unsigned(97,8) ,
15807	 => std_logic_vector(to_unsigned(119,8) ,
15808	 => std_logic_vector(to_unsigned(130,8) ,
15809	 => std_logic_vector(to_unsigned(109,8) ,
15810	 => std_logic_vector(to_unsigned(112,8) ,
15811	 => std_logic_vector(to_unsigned(122,8) ,
15812	 => std_logic_vector(to_unsigned(124,8) ,
15813	 => std_logic_vector(to_unsigned(125,8) ,
15814	 => std_logic_vector(to_unsigned(122,8) ,
15815	 => std_logic_vector(to_unsigned(119,8) ,
15816	 => std_logic_vector(to_unsigned(119,8) ,
15817	 => std_logic_vector(to_unsigned(116,8) ,
15818	 => std_logic_vector(to_unsigned(118,8) ,
15819	 => std_logic_vector(to_unsigned(118,8) ,
15820	 => std_logic_vector(to_unsigned(112,8) ,
15821	 => std_logic_vector(to_unsigned(109,8) ,
15822	 => std_logic_vector(to_unsigned(114,8) ,
15823	 => std_logic_vector(to_unsigned(115,8) ,
15824	 => std_logic_vector(to_unsigned(114,8) ,
15825	 => std_logic_vector(to_unsigned(108,8) ,
15826	 => std_logic_vector(to_unsigned(112,8) ,
15827	 => std_logic_vector(to_unsigned(95,8) ,
15828	 => std_logic_vector(to_unsigned(88,8) ,
15829	 => std_logic_vector(to_unsigned(90,8) ,
15830	 => std_logic_vector(to_unsigned(90,8) ,
15831	 => std_logic_vector(to_unsigned(84,8) ,
15832	 => std_logic_vector(to_unsigned(100,8) ,
15833	 => std_logic_vector(to_unsigned(100,8) ,
15834	 => std_logic_vector(to_unsigned(82,8) ,
15835	 => std_logic_vector(to_unsigned(91,8) ,
15836	 => std_logic_vector(to_unsigned(96,8) ,
15837	 => std_logic_vector(to_unsigned(81,8) ,
15838	 => std_logic_vector(to_unsigned(82,8) ,
15839	 => std_logic_vector(to_unsigned(87,8) ,
15840	 => std_logic_vector(to_unsigned(79,8) ,
15841	 => std_logic_vector(to_unsigned(81,8) ,
15842	 => std_logic_vector(to_unsigned(108,8) ,
15843	 => std_logic_vector(to_unsigned(107,8) ,
15844	 => std_logic_vector(to_unsigned(91,8) ,
15845	 => std_logic_vector(to_unsigned(90,8) ,
15846	 => std_logic_vector(to_unsigned(93,8) ,
15847	 => std_logic_vector(to_unsigned(95,8) ,
15848	 => std_logic_vector(to_unsigned(93,8) ,
15849	 => std_logic_vector(to_unsigned(86,8) ,
15850	 => std_logic_vector(to_unsigned(91,8) ,
15851	 => std_logic_vector(to_unsigned(97,8) ,
15852	 => std_logic_vector(to_unsigned(78,8) ,
15853	 => std_logic_vector(to_unsigned(82,8) ,
15854	 => std_logic_vector(to_unsigned(91,8) ,
15855	 => std_logic_vector(to_unsigned(81,8) ,
15856	 => std_logic_vector(to_unsigned(87,8) ,
15857	 => std_logic_vector(to_unsigned(90,8) ,
15858	 => std_logic_vector(to_unsigned(96,8) ,
15859	 => std_logic_vector(to_unsigned(109,8) ,
15860	 => std_logic_vector(to_unsigned(105,8) ,
15861	 => std_logic_vector(to_unsigned(103,8) ,
15862	 => std_logic_vector(to_unsigned(105,8) ,
15863	 => std_logic_vector(to_unsigned(96,8) ,
15864	 => std_logic_vector(to_unsigned(100,8) ,
15865	 => std_logic_vector(to_unsigned(96,8) ,
15866	 => std_logic_vector(to_unsigned(79,8) ,
15867	 => std_logic_vector(to_unsigned(78,8) ,
15868	 => std_logic_vector(to_unsigned(103,8) ,
15869	 => std_logic_vector(to_unsigned(104,8) ,
15870	 => std_logic_vector(to_unsigned(95,8) ,
15871	 => std_logic_vector(to_unsigned(90,8) ,
15872	 => std_logic_vector(to_unsigned(112,8) ,
15873	 => std_logic_vector(to_unsigned(124,8) ,
15874	 => std_logic_vector(to_unsigned(133,8) ,
15875	 => std_logic_vector(to_unsigned(119,8) ,
15876	 => std_logic_vector(to_unsigned(122,8) ,
15877	 => std_logic_vector(to_unsigned(131,8) ,
15878	 => std_logic_vector(to_unsigned(121,8) ,
15879	 => std_logic_vector(to_unsigned(125,8) ,
15880	 => std_logic_vector(to_unsigned(131,8) ,
15881	 => std_logic_vector(to_unsigned(122,8) ,
15882	 => std_logic_vector(to_unsigned(108,8) ,
15883	 => std_logic_vector(to_unsigned(108,8) ,
15884	 => std_logic_vector(to_unsigned(96,8) ,
15885	 => std_logic_vector(to_unsigned(100,8) ,
15886	 => std_logic_vector(to_unsigned(99,8) ,
15887	 => std_logic_vector(to_unsigned(101,8) ,
15888	 => std_logic_vector(to_unsigned(127,8) ,
15889	 => std_logic_vector(to_unsigned(114,8) ,
15890	 => std_logic_vector(to_unsigned(71,8) ,
15891	 => std_logic_vector(to_unsigned(86,8) ,
15892	 => std_logic_vector(to_unsigned(99,8) ,
15893	 => std_logic_vector(to_unsigned(91,8) ,
15894	 => std_logic_vector(to_unsigned(71,8) ,
15895	 => std_logic_vector(to_unsigned(73,8) ,
15896	 => std_logic_vector(to_unsigned(73,8) ,
15897	 => std_logic_vector(to_unsigned(79,8) ,
15898	 => std_logic_vector(to_unsigned(87,8) ,
15899	 => std_logic_vector(to_unsigned(80,8) ,
15900	 => std_logic_vector(to_unsigned(86,8) ,
15901	 => std_logic_vector(to_unsigned(101,8) ,
15902	 => std_logic_vector(to_unsigned(90,8) ,
15903	 => std_logic_vector(to_unsigned(85,8) ,
15904	 => std_logic_vector(to_unsigned(73,8) ,
15905	 => std_logic_vector(to_unsigned(76,8) ,
15906	 => std_logic_vector(to_unsigned(80,8) ,
15907	 => std_logic_vector(to_unsigned(69,8) ,
15908	 => std_logic_vector(to_unsigned(70,8) ,
15909	 => std_logic_vector(to_unsigned(66,8) ,
15910	 => std_logic_vector(to_unsigned(71,8) ,
15911	 => std_logic_vector(to_unsigned(78,8) ,
15912	 => std_logic_vector(to_unsigned(63,8) ,
15913	 => std_logic_vector(to_unsigned(63,8) ,
15914	 => std_logic_vector(to_unsigned(64,8) ,
15915	 => std_logic_vector(to_unsigned(58,8) ,
15916	 => std_logic_vector(to_unsigned(62,8) ,
15917	 => std_logic_vector(to_unsigned(63,8) ,
15918	 => std_logic_vector(to_unsigned(62,8) ,
15919	 => std_logic_vector(to_unsigned(61,8) ,
15920	 => std_logic_vector(to_unsigned(68,8) ,
15921	 => std_logic_vector(to_unsigned(61,8) ,
15922	 => std_logic_vector(to_unsigned(63,8) ,
15923	 => std_logic_vector(to_unsigned(68,8) ,
15924	 => std_logic_vector(to_unsigned(69,8) ,
15925	 => std_logic_vector(to_unsigned(64,8) ,
15926	 => std_logic_vector(to_unsigned(59,8) ,
15927	 => std_logic_vector(to_unsigned(32,8) ,
15928	 => std_logic_vector(to_unsigned(1,8) ,
15929	 => std_logic_vector(to_unsigned(0,8) ,
15930	 => std_logic_vector(to_unsigned(2,8) ,
15931	 => std_logic_vector(to_unsigned(46,8) ,
15932	 => std_logic_vector(to_unsigned(70,8) ,
15933	 => std_logic_vector(to_unsigned(67,8) ,
15934	 => std_logic_vector(to_unsigned(66,8) ,
15935	 => std_logic_vector(to_unsigned(77,8) ,
15936	 => std_logic_vector(to_unsigned(77,8) ,
15937	 => std_logic_vector(to_unsigned(78,8) ,
15938	 => std_logic_vector(to_unsigned(79,8) ,
15939	 => std_logic_vector(to_unsigned(85,8) ,
15940	 => std_logic_vector(to_unsigned(80,8) ,
15941	 => std_logic_vector(to_unsigned(76,8) ,
15942	 => std_logic_vector(to_unsigned(79,8) ,
15943	 => std_logic_vector(to_unsigned(68,8) ,
15944	 => std_logic_vector(to_unsigned(65,8) ,
15945	 => std_logic_vector(to_unsigned(73,8) ,
15946	 => std_logic_vector(to_unsigned(73,8) ,
15947	 => std_logic_vector(to_unsigned(81,8) ,
15948	 => std_logic_vector(to_unsigned(87,8) ,
15949	 => std_logic_vector(to_unsigned(86,8) ,
15950	 => std_logic_vector(to_unsigned(80,8) ,
15951	 => std_logic_vector(to_unsigned(74,8) ,
15952	 => std_logic_vector(to_unsigned(70,8) ,
15953	 => std_logic_vector(to_unsigned(64,8) ,
15954	 => std_logic_vector(to_unsigned(69,8) ,
15955	 => std_logic_vector(to_unsigned(57,8) ,
15956	 => std_logic_vector(to_unsigned(58,8) ,
15957	 => std_logic_vector(to_unsigned(69,8) ,
15958	 => std_logic_vector(to_unsigned(69,8) ,
15959	 => std_logic_vector(to_unsigned(68,8) ,
15960	 => std_logic_vector(to_unsigned(68,8) ,
15961	 => std_logic_vector(to_unsigned(65,8) ,
15962	 => std_logic_vector(to_unsigned(71,8) ,
15963	 => std_logic_vector(to_unsigned(80,8) ,
15964	 => std_logic_vector(to_unsigned(81,8) ,
15965	 => std_logic_vector(to_unsigned(76,8) ,
15966	 => std_logic_vector(to_unsigned(74,8) ,
15967	 => std_logic_vector(to_unsigned(70,8) ,
15968	 => std_logic_vector(to_unsigned(70,8) ,
15969	 => std_logic_vector(to_unsigned(88,8) ,
15970	 => std_logic_vector(to_unsigned(73,8) ,
15971	 => std_logic_vector(to_unsigned(65,8) ,
15972	 => std_logic_vector(to_unsigned(77,8) ,
15973	 => std_logic_vector(to_unsigned(81,8) ,
15974	 => std_logic_vector(to_unsigned(79,8) ,
15975	 => std_logic_vector(to_unsigned(78,8) ,
15976	 => std_logic_vector(to_unsigned(85,8) ,
15977	 => std_logic_vector(to_unsigned(95,8) ,
15978	 => std_logic_vector(to_unsigned(79,8) ,
15979	 => std_logic_vector(to_unsigned(77,8) ,
15980	 => std_logic_vector(to_unsigned(76,8) ,
15981	 => std_logic_vector(to_unsigned(80,8) ,
15982	 => std_logic_vector(to_unsigned(80,8) ,
15983	 => std_logic_vector(to_unsigned(85,8) ,
15984	 => std_logic_vector(to_unsigned(86,8) ,
15985	 => std_logic_vector(to_unsigned(88,8) ,
15986	 => std_logic_vector(to_unsigned(93,8) ,
15987	 => std_logic_vector(to_unsigned(91,8) ,
15988	 => std_logic_vector(to_unsigned(87,8) ,
15989	 => std_logic_vector(to_unsigned(82,8) ,
15990	 => std_logic_vector(to_unsigned(87,8) ,
15991	 => std_logic_vector(to_unsigned(90,8) ,
15992	 => std_logic_vector(to_unsigned(95,8) ,
15993	 => std_logic_vector(to_unsigned(88,8) ,
15994	 => std_logic_vector(to_unsigned(88,8) ,
15995	 => std_logic_vector(to_unsigned(81,8) ,
15996	 => std_logic_vector(to_unsigned(79,8) ,
15997	 => std_logic_vector(to_unsigned(90,8) ,
15998	 => std_logic_vector(to_unsigned(95,8) ,
15999	 => std_logic_vector(to_unsigned(92,8) ,
16000	 => std_logic_vector(to_unsigned(96,8) ,
16001	 => std_logic_vector(to_unsigned(144,8) ,
16002	 => std_logic_vector(to_unsigned(146,8) ,
16003	 => std_logic_vector(to_unsigned(154,8) ,
16004	 => std_logic_vector(to_unsigned(161,8) ,
16005	 => std_logic_vector(to_unsigned(161,8) ,
16006	 => std_logic_vector(to_unsigned(159,8) ,
16007	 => std_logic_vector(to_unsigned(156,8) ,
16008	 => std_logic_vector(to_unsigned(154,8) ,
16009	 => std_logic_vector(to_unsigned(159,8) ,
16010	 => std_logic_vector(to_unsigned(163,8) ,
16011	 => std_logic_vector(to_unsigned(161,8) ,
16012	 => std_logic_vector(to_unsigned(159,8) ,
16013	 => std_logic_vector(to_unsigned(157,8) ,
16014	 => std_logic_vector(to_unsigned(156,8) ,
16015	 => std_logic_vector(to_unsigned(154,8) ,
16016	 => std_logic_vector(to_unsigned(154,8) ,
16017	 => std_logic_vector(to_unsigned(154,8) ,
16018	 => std_logic_vector(to_unsigned(156,8) ,
16019	 => std_logic_vector(to_unsigned(154,8) ,
16020	 => std_logic_vector(to_unsigned(161,8) ,
16021	 => std_logic_vector(to_unsigned(157,8) ,
16022	 => std_logic_vector(to_unsigned(154,8) ,
16023	 => std_logic_vector(to_unsigned(159,8) ,
16024	 => std_logic_vector(to_unsigned(161,8) ,
16025	 => std_logic_vector(to_unsigned(157,8) ,
16026	 => std_logic_vector(to_unsigned(156,8) ,
16027	 => std_logic_vector(to_unsigned(152,8) ,
16028	 => std_logic_vector(to_unsigned(142,8) ,
16029	 => std_logic_vector(to_unsigned(141,8) ,
16030	 => std_logic_vector(to_unsigned(146,8) ,
16031	 => std_logic_vector(to_unsigned(149,8) ,
16032	 => std_logic_vector(to_unsigned(141,8) ,
16033	 => std_logic_vector(to_unsigned(139,8) ,
16034	 => std_logic_vector(to_unsigned(142,8) ,
16035	 => std_logic_vector(to_unsigned(136,8) ,
16036	 => std_logic_vector(to_unsigned(136,8) ,
16037	 => std_logic_vector(to_unsigned(139,8) ,
16038	 => std_logic_vector(to_unsigned(142,8) ,
16039	 => std_logic_vector(to_unsigned(141,8) ,
16040	 => std_logic_vector(to_unsigned(138,8) ,
16041	 => std_logic_vector(to_unsigned(141,8) ,
16042	 => std_logic_vector(to_unsigned(146,8) ,
16043	 => std_logic_vector(to_unsigned(141,8) ,
16044	 => std_logic_vector(to_unsigned(147,8) ,
16045	 => std_logic_vector(to_unsigned(154,8) ,
16046	 => std_logic_vector(to_unsigned(154,8) ,
16047	 => std_logic_vector(to_unsigned(154,8) ,
16048	 => std_logic_vector(to_unsigned(151,8) ,
16049	 => std_logic_vector(to_unsigned(149,8) ,
16050	 => std_logic_vector(to_unsigned(157,8) ,
16051	 => std_logic_vector(to_unsigned(157,8) ,
16052	 => std_logic_vector(to_unsigned(156,8) ,
16053	 => std_logic_vector(to_unsigned(152,8) ,
16054	 => std_logic_vector(to_unsigned(147,8) ,
16055	 => std_logic_vector(to_unsigned(133,8) ,
16056	 => std_logic_vector(to_unsigned(127,8) ,
16057	 => std_logic_vector(to_unsigned(134,8) ,
16058	 => std_logic_vector(to_unsigned(138,8) ,
16059	 => std_logic_vector(to_unsigned(121,8) ,
16060	 => std_logic_vector(to_unsigned(122,8) ,
16061	 => std_logic_vector(to_unsigned(127,8) ,
16062	 => std_logic_vector(to_unsigned(139,8) ,
16063	 => std_logic_vector(to_unsigned(152,8) ,
16064	 => std_logic_vector(to_unsigned(141,8) ,
16065	 => std_logic_vector(to_unsigned(130,8) ,
16066	 => std_logic_vector(to_unsigned(131,8) ,
16067	 => std_logic_vector(to_unsigned(144,8) ,
16068	 => std_logic_vector(to_unsigned(149,8) ,
16069	 => std_logic_vector(to_unsigned(136,8) ,
16070	 => std_logic_vector(to_unsigned(130,8) ,
16071	 => std_logic_vector(to_unsigned(151,8) ,
16072	 => std_logic_vector(to_unsigned(152,8) ,
16073	 => std_logic_vector(to_unsigned(147,8) ,
16074	 => std_logic_vector(to_unsigned(156,8) ,
16075	 => std_logic_vector(to_unsigned(163,8) ,
16076	 => std_logic_vector(to_unsigned(166,8) ,
16077	 => std_logic_vector(to_unsigned(163,8) ,
16078	 => std_logic_vector(to_unsigned(156,8) ,
16079	 => std_logic_vector(to_unsigned(149,8) ,
16080	 => std_logic_vector(to_unsigned(121,8) ,
16081	 => std_logic_vector(to_unsigned(112,8) ,
16082	 => std_logic_vector(to_unsigned(141,8) ,
16083	 => std_logic_vector(to_unsigned(151,8) ,
16084	 => std_logic_vector(to_unsigned(147,8) ,
16085	 => std_logic_vector(to_unsigned(156,8) ,
16086	 => std_logic_vector(to_unsigned(161,8) ,
16087	 => std_logic_vector(to_unsigned(163,8) ,
16088	 => std_logic_vector(to_unsigned(163,8) ,
16089	 => std_logic_vector(to_unsigned(163,8) ,
16090	 => std_logic_vector(to_unsigned(159,8) ,
16091	 => std_logic_vector(to_unsigned(163,8) ,
16092	 => std_logic_vector(to_unsigned(177,8) ,
16093	 => std_logic_vector(to_unsigned(190,8) ,
16094	 => std_logic_vector(to_unsigned(194,8) ,
16095	 => std_logic_vector(to_unsigned(186,8) ,
16096	 => std_logic_vector(to_unsigned(186,8) ,
16097	 => std_logic_vector(to_unsigned(179,8) ,
16098	 => std_logic_vector(to_unsigned(177,8) ,
16099	 => std_logic_vector(to_unsigned(163,8) ,
16100	 => std_logic_vector(to_unsigned(152,8) ,
16101	 => std_logic_vector(to_unsigned(156,8) ,
16102	 => std_logic_vector(to_unsigned(159,8) ,
16103	 => std_logic_vector(to_unsigned(157,8) ,
16104	 => std_logic_vector(to_unsigned(154,8) ,
16105	 => std_logic_vector(to_unsigned(154,8) ,
16106	 => std_logic_vector(to_unsigned(142,8) ,
16107	 => std_logic_vector(to_unsigned(139,8) ,
16108	 => std_logic_vector(to_unsigned(147,8) ,
16109	 => std_logic_vector(to_unsigned(154,8) ,
16110	 => std_logic_vector(to_unsigned(166,8) ,
16111	 => std_logic_vector(to_unsigned(141,8) ,
16112	 => std_logic_vector(to_unsigned(131,8) ,
16113	 => std_logic_vector(to_unsigned(125,8) ,
16114	 => std_logic_vector(to_unsigned(127,8) ,
16115	 => std_logic_vector(to_unsigned(121,8) ,
16116	 => std_logic_vector(to_unsigned(121,8) ,
16117	 => std_logic_vector(to_unsigned(114,8) ,
16118	 => std_logic_vector(to_unsigned(124,8) ,
16119	 => std_logic_vector(to_unsigned(124,8) ,
16120	 => std_logic_vector(to_unsigned(101,8) ,
16121	 => std_logic_vector(to_unsigned(131,8) ,
16122	 => std_logic_vector(to_unsigned(146,8) ,
16123	 => std_logic_vector(to_unsigned(134,8) ,
16124	 => std_logic_vector(to_unsigned(119,8) ,
16125	 => std_logic_vector(to_unsigned(101,8) ,
16126	 => std_logic_vector(to_unsigned(107,8) ,
16127	 => std_logic_vector(to_unsigned(125,8) ,
16128	 => std_logic_vector(to_unsigned(131,8) ,
16129	 => std_logic_vector(to_unsigned(114,8) ,
16130	 => std_logic_vector(to_unsigned(114,8) ,
16131	 => std_logic_vector(to_unsigned(116,8) ,
16132	 => std_logic_vector(to_unsigned(116,8) ,
16133	 => std_logic_vector(to_unsigned(121,8) ,
16134	 => std_logic_vector(to_unsigned(119,8) ,
16135	 => std_logic_vector(to_unsigned(122,8) ,
16136	 => std_logic_vector(to_unsigned(128,8) ,
16137	 => std_logic_vector(to_unsigned(124,8) ,
16138	 => std_logic_vector(to_unsigned(124,8) ,
16139	 => std_logic_vector(to_unsigned(118,8) ,
16140	 => std_logic_vector(to_unsigned(109,8) ,
16141	 => std_logic_vector(to_unsigned(111,8) ,
16142	 => std_logic_vector(to_unsigned(116,8) ,
16143	 => std_logic_vector(to_unsigned(116,8) ,
16144	 => std_logic_vector(to_unsigned(122,8) ,
16145	 => std_logic_vector(to_unsigned(125,8) ,
16146	 => std_logic_vector(to_unsigned(101,8) ,
16147	 => std_logic_vector(to_unsigned(80,8) ,
16148	 => std_logic_vector(to_unsigned(86,8) ,
16149	 => std_logic_vector(to_unsigned(81,8) ,
16150	 => std_logic_vector(to_unsigned(82,8) ,
16151	 => std_logic_vector(to_unsigned(71,8) ,
16152	 => std_logic_vector(to_unsigned(85,8) ,
16153	 => std_logic_vector(to_unsigned(84,8) ,
16154	 => std_logic_vector(to_unsigned(114,8) ,
16155	 => std_logic_vector(to_unsigned(107,8) ,
16156	 => std_logic_vector(to_unsigned(91,8) ,
16157	 => std_logic_vector(to_unsigned(86,8) ,
16158	 => std_logic_vector(to_unsigned(82,8) ,
16159	 => std_logic_vector(to_unsigned(80,8) ,
16160	 => std_logic_vector(to_unsigned(80,8) ,
16161	 => std_logic_vector(to_unsigned(85,8) ,
16162	 => std_logic_vector(to_unsigned(96,8) ,
16163	 => std_logic_vector(to_unsigned(107,8) ,
16164	 => std_logic_vector(to_unsigned(96,8) ,
16165	 => std_logic_vector(to_unsigned(88,8) ,
16166	 => std_logic_vector(to_unsigned(88,8) ,
16167	 => std_logic_vector(to_unsigned(87,8) ,
16168	 => std_logic_vector(to_unsigned(95,8) ,
16169	 => std_logic_vector(to_unsigned(93,8) ,
16170	 => std_logic_vector(to_unsigned(92,8) ,
16171	 => std_logic_vector(to_unsigned(104,8) ,
16172	 => std_logic_vector(to_unsigned(80,8) ,
16173	 => std_logic_vector(to_unsigned(65,8) ,
16174	 => std_logic_vector(to_unsigned(78,8) ,
16175	 => std_logic_vector(to_unsigned(86,8) ,
16176	 => std_logic_vector(to_unsigned(92,8) ,
16177	 => std_logic_vector(to_unsigned(84,8) ,
16178	 => std_logic_vector(to_unsigned(87,8) ,
16179	 => std_logic_vector(to_unsigned(104,8) ,
16180	 => std_logic_vector(to_unsigned(100,8) ,
16181	 => std_logic_vector(to_unsigned(95,8) ,
16182	 => std_logic_vector(to_unsigned(99,8) ,
16183	 => std_logic_vector(to_unsigned(99,8) ,
16184	 => std_logic_vector(to_unsigned(73,8) ,
16185	 => std_logic_vector(to_unsigned(73,8) ,
16186	 => std_logic_vector(to_unsigned(78,8) ,
16187	 => std_logic_vector(to_unsigned(86,8) ,
16188	 => std_logic_vector(to_unsigned(99,8) ,
16189	 => std_logic_vector(to_unsigned(86,8) ,
16190	 => std_logic_vector(to_unsigned(76,8) ,
16191	 => std_logic_vector(to_unsigned(81,8) ,
16192	 => std_logic_vector(to_unsigned(111,8) ,
16193	 => std_logic_vector(to_unsigned(128,8) ,
16194	 => std_logic_vector(to_unsigned(133,8) ,
16195	 => std_logic_vector(to_unsigned(119,8) ,
16196	 => std_logic_vector(to_unsigned(121,8) ,
16197	 => std_logic_vector(to_unsigned(130,8) ,
16198	 => std_logic_vector(to_unsigned(121,8) ,
16199	 => std_logic_vector(to_unsigned(122,8) ,
16200	 => std_logic_vector(to_unsigned(128,8) ,
16201	 => std_logic_vector(to_unsigned(109,8) ,
16202	 => std_logic_vector(to_unsigned(104,8) ,
16203	 => std_logic_vector(to_unsigned(111,8) ,
16204	 => std_logic_vector(to_unsigned(92,8) ,
16205	 => std_logic_vector(to_unsigned(96,8) ,
16206	 => std_logic_vector(to_unsigned(99,8) ,
16207	 => std_logic_vector(to_unsigned(105,8) ,
16208	 => std_logic_vector(to_unsigned(116,8) ,
16209	 => std_logic_vector(to_unsigned(97,8) ,
16210	 => std_logic_vector(to_unsigned(70,8) ,
16211	 => std_logic_vector(to_unsigned(90,8) ,
16212	 => std_logic_vector(to_unsigned(92,8) ,
16213	 => std_logic_vector(to_unsigned(80,8) ,
16214	 => std_logic_vector(to_unsigned(77,8) ,
16215	 => std_logic_vector(to_unsigned(65,8) ,
16216	 => std_logic_vector(to_unsigned(68,8) ,
16217	 => std_logic_vector(to_unsigned(72,8) ,
16218	 => std_logic_vector(to_unsigned(73,8) ,
16219	 => std_logic_vector(to_unsigned(68,8) ,
16220	 => std_logic_vector(to_unsigned(67,8) ,
16221	 => std_logic_vector(to_unsigned(79,8) ,
16222	 => std_logic_vector(to_unsigned(90,8) ,
16223	 => std_logic_vector(to_unsigned(91,8) ,
16224	 => std_logic_vector(to_unsigned(79,8) ,
16225	 => std_logic_vector(to_unsigned(74,8) ,
16226	 => std_logic_vector(to_unsigned(85,8) ,
16227	 => std_logic_vector(to_unsigned(72,8) ,
16228	 => std_logic_vector(to_unsigned(72,8) ,
16229	 => std_logic_vector(to_unsigned(73,8) ,
16230	 => std_logic_vector(to_unsigned(68,8) ,
16231	 => std_logic_vector(to_unsigned(64,8) ,
16232	 => std_logic_vector(to_unsigned(53,8) ,
16233	 => std_logic_vector(to_unsigned(57,8) ,
16234	 => std_logic_vector(to_unsigned(59,8) ,
16235	 => std_logic_vector(to_unsigned(56,8) ,
16236	 => std_logic_vector(to_unsigned(58,8) ,
16237	 => std_logic_vector(to_unsigned(56,8) ,
16238	 => std_logic_vector(to_unsigned(67,8) ,
16239	 => std_logic_vector(to_unsigned(64,8) ,
16240	 => std_logic_vector(to_unsigned(65,8) ,
16241	 => std_logic_vector(to_unsigned(66,8) ,
16242	 => std_logic_vector(to_unsigned(72,8) ,
16243	 => std_logic_vector(to_unsigned(80,8) ,
16244	 => std_logic_vector(to_unsigned(78,8) ,
16245	 => std_logic_vector(to_unsigned(70,8) ,
16246	 => std_logic_vector(to_unsigned(60,8) ,
16247	 => std_logic_vector(to_unsigned(52,8) ,
16248	 => std_logic_vector(to_unsigned(5,8) ,
16249	 => std_logic_vector(to_unsigned(0,8) ,
16250	 => std_logic_vector(to_unsigned(0,8) ,
16251	 => std_logic_vector(to_unsigned(25,8) ,
16252	 => std_logic_vector(to_unsigned(74,8) ,
16253	 => std_logic_vector(to_unsigned(73,8) ,
16254	 => std_logic_vector(to_unsigned(74,8) ,
16255	 => std_logic_vector(to_unsigned(68,8) ,
16256	 => std_logic_vector(to_unsigned(64,8) ,
16257	 => std_logic_vector(to_unsigned(69,8) ,
16258	 => std_logic_vector(to_unsigned(84,8) ,
16259	 => std_logic_vector(to_unsigned(86,8) ,
16260	 => std_logic_vector(to_unsigned(80,8) ,
16261	 => std_logic_vector(to_unsigned(72,8) ,
16262	 => std_logic_vector(to_unsigned(72,8) ,
16263	 => std_logic_vector(to_unsigned(76,8) ,
16264	 => std_logic_vector(to_unsigned(78,8) ,
16265	 => std_logic_vector(to_unsigned(77,8) ,
16266	 => std_logic_vector(to_unsigned(80,8) ,
16267	 => std_logic_vector(to_unsigned(86,8) ,
16268	 => std_logic_vector(to_unsigned(81,8) ,
16269	 => std_logic_vector(to_unsigned(86,8) ,
16270	 => std_logic_vector(to_unsigned(87,8) ,
16271	 => std_logic_vector(to_unsigned(76,8) ,
16272	 => std_logic_vector(to_unsigned(62,8) ,
16273	 => std_logic_vector(to_unsigned(68,8) ,
16274	 => std_logic_vector(to_unsigned(73,8) ,
16275	 => std_logic_vector(to_unsigned(69,8) ,
16276	 => std_logic_vector(to_unsigned(76,8) ,
16277	 => std_logic_vector(to_unsigned(70,8) ,
16278	 => std_logic_vector(to_unsigned(74,8) ,
16279	 => std_logic_vector(to_unsigned(77,8) ,
16280	 => std_logic_vector(to_unsigned(69,8) ,
16281	 => std_logic_vector(to_unsigned(71,8) ,
16282	 => std_logic_vector(to_unsigned(78,8) ,
16283	 => std_logic_vector(to_unsigned(82,8) ,
16284	 => std_logic_vector(to_unsigned(77,8) ,
16285	 => std_logic_vector(to_unsigned(72,8) ,
16286	 => std_logic_vector(to_unsigned(76,8) ,
16287	 => std_logic_vector(to_unsigned(76,8) ,
16288	 => std_logic_vector(to_unsigned(76,8) ,
16289	 => std_logic_vector(to_unsigned(72,8) ,
16290	 => std_logic_vector(to_unsigned(77,8) ,
16291	 => std_logic_vector(to_unsigned(76,8) ,
16292	 => std_logic_vector(to_unsigned(81,8) ,
16293	 => std_logic_vector(to_unsigned(81,8) ,
16294	 => std_logic_vector(to_unsigned(65,8) ,
16295	 => std_logic_vector(to_unsigned(74,8) ,
16296	 => std_logic_vector(to_unsigned(92,8) ,
16297	 => std_logic_vector(to_unsigned(96,8) ,
16298	 => std_logic_vector(to_unsigned(86,8) ,
16299	 => std_logic_vector(to_unsigned(79,8) ,
16300	 => std_logic_vector(to_unsigned(72,8) ,
16301	 => std_logic_vector(to_unsigned(77,8) ,
16302	 => std_logic_vector(to_unsigned(81,8) ,
16303	 => std_logic_vector(to_unsigned(86,8) ,
16304	 => std_logic_vector(to_unsigned(87,8) ,
16305	 => std_logic_vector(to_unsigned(86,8) ,
16306	 => std_logic_vector(to_unsigned(88,8) ,
16307	 => std_logic_vector(to_unsigned(87,8) ,
16308	 => std_logic_vector(to_unsigned(84,8) ,
16309	 => std_logic_vector(to_unsigned(82,8) ,
16310	 => std_logic_vector(to_unsigned(86,8) ,
16311	 => std_logic_vector(to_unsigned(90,8) ,
16312	 => std_logic_vector(to_unsigned(96,8) ,
16313	 => std_logic_vector(to_unsigned(93,8) ,
16314	 => std_logic_vector(to_unsigned(87,8) ,
16315	 => std_logic_vector(to_unsigned(93,8) ,
16316	 => std_logic_vector(to_unsigned(95,8) ,
16317	 => std_logic_vector(to_unsigned(90,8) ,
16318	 => std_logic_vector(to_unsigned(88,8) ,
16319	 => std_logic_vector(to_unsigned(90,8) ,
16320	 => std_logic_vector(to_unsigned(93,8) ,
16321	 => std_logic_vector(to_unsigned(149,8) ,
16322	 => std_logic_vector(to_unsigned(146,8) ,
16323	 => std_logic_vector(to_unsigned(147,8) ,
16324	 => std_logic_vector(to_unsigned(154,8) ,
16325	 => std_logic_vector(to_unsigned(157,8) ,
16326	 => std_logic_vector(to_unsigned(156,8) ,
16327	 => std_logic_vector(to_unsigned(152,8) ,
16328	 => std_logic_vector(to_unsigned(154,8) ,
16329	 => std_logic_vector(to_unsigned(154,8) ,
16330	 => std_logic_vector(to_unsigned(157,8) ,
16331	 => std_logic_vector(to_unsigned(161,8) ,
16332	 => std_logic_vector(to_unsigned(159,8) ,
16333	 => std_logic_vector(to_unsigned(157,8) ,
16334	 => std_logic_vector(to_unsigned(156,8) ,
16335	 => std_logic_vector(to_unsigned(152,8) ,
16336	 => std_logic_vector(to_unsigned(152,8) ,
16337	 => std_logic_vector(to_unsigned(152,8) ,
16338	 => std_logic_vector(to_unsigned(147,8) ,
16339	 => std_logic_vector(to_unsigned(149,8) ,
16340	 => std_logic_vector(to_unsigned(159,8) ,
16341	 => std_logic_vector(to_unsigned(154,8) ,
16342	 => std_logic_vector(to_unsigned(151,8) ,
16343	 => std_logic_vector(to_unsigned(161,8) ,
16344	 => std_logic_vector(to_unsigned(161,8) ,
16345	 => std_logic_vector(to_unsigned(156,8) ,
16346	 => std_logic_vector(to_unsigned(157,8) ,
16347	 => std_logic_vector(to_unsigned(154,8) ,
16348	 => std_logic_vector(to_unsigned(144,8) ,
16349	 => std_logic_vector(to_unsigned(149,8) ,
16350	 => std_logic_vector(to_unsigned(146,8) ,
16351	 => std_logic_vector(to_unsigned(144,8) ,
16352	 => std_logic_vector(to_unsigned(131,8) ,
16353	 => std_logic_vector(to_unsigned(119,8) ,
16354	 => std_logic_vector(to_unsigned(125,8) ,
16355	 => std_logic_vector(to_unsigned(141,8) ,
16356	 => std_logic_vector(to_unsigned(144,8) ,
16357	 => std_logic_vector(to_unsigned(136,8) ,
16358	 => std_logic_vector(to_unsigned(138,8) ,
16359	 => std_logic_vector(to_unsigned(139,8) ,
16360	 => std_logic_vector(to_unsigned(133,8) ,
16361	 => std_logic_vector(to_unsigned(136,8) ,
16362	 => std_logic_vector(to_unsigned(144,8) ,
16363	 => std_logic_vector(to_unsigned(138,8) ,
16364	 => std_logic_vector(to_unsigned(142,8) ,
16365	 => std_logic_vector(to_unsigned(157,8) ,
16366	 => std_logic_vector(to_unsigned(157,8) ,
16367	 => std_logic_vector(to_unsigned(149,8) ,
16368	 => std_logic_vector(to_unsigned(151,8) ,
16369	 => std_logic_vector(to_unsigned(156,8) ,
16370	 => std_logic_vector(to_unsigned(156,8) ,
16371	 => std_logic_vector(to_unsigned(156,8) ,
16372	 => std_logic_vector(to_unsigned(154,8) ,
16373	 => std_logic_vector(to_unsigned(156,8) ,
16374	 => std_logic_vector(to_unsigned(152,8) ,
16375	 => std_logic_vector(to_unsigned(138,8) ,
16376	 => std_logic_vector(to_unsigned(142,8) ,
16377	 => std_logic_vector(to_unsigned(152,8) ,
16378	 => std_logic_vector(to_unsigned(142,8) ,
16379	 => std_logic_vector(to_unsigned(131,8) ,
16380	 => std_logic_vector(to_unsigned(138,8) ,
16381	 => std_logic_vector(to_unsigned(128,8) ,
16382	 => std_logic_vector(to_unsigned(125,8) ,
16383	 => std_logic_vector(to_unsigned(133,8) ,
16384	 => std_logic_vector(to_unsigned(146,8) ,
16385	 => std_logic_vector(to_unsigned(133,8) ,
16386	 => std_logic_vector(to_unsigned(134,8) ,
16387	 => std_logic_vector(to_unsigned(141,8) ,
16388	 => std_logic_vector(to_unsigned(154,8) ,
16389	 => std_logic_vector(to_unsigned(157,8) ,
16390	 => std_logic_vector(to_unsigned(131,8) ,
16391	 => std_logic_vector(to_unsigned(142,8) ,
16392	 => std_logic_vector(to_unsigned(156,8) ,
16393	 => std_logic_vector(to_unsigned(157,8) ,
16394	 => std_logic_vector(to_unsigned(151,8) ,
16395	 => std_logic_vector(to_unsigned(154,8) ,
16396	 => std_logic_vector(to_unsigned(154,8) ,
16397	 => std_logic_vector(to_unsigned(157,8) ,
16398	 => std_logic_vector(to_unsigned(157,8) ,
16399	 => std_logic_vector(to_unsigned(141,8) ,
16400	 => std_logic_vector(to_unsigned(118,8) ,
16401	 => std_logic_vector(to_unsigned(115,8) ,
16402	 => std_logic_vector(to_unsigned(122,8) ,
16403	 => std_logic_vector(to_unsigned(138,8) ,
16404	 => std_logic_vector(to_unsigned(151,8) ,
16405	 => std_logic_vector(to_unsigned(159,8) ,
16406	 => std_logic_vector(to_unsigned(161,8) ,
16407	 => std_logic_vector(to_unsigned(164,8) ,
16408	 => std_logic_vector(to_unsigned(168,8) ,
16409	 => std_logic_vector(to_unsigned(156,8) ,
16410	 => std_logic_vector(to_unsigned(164,8) ,
16411	 => std_logic_vector(to_unsigned(190,8) ,
16412	 => std_logic_vector(to_unsigned(152,8) ,
16413	 => std_logic_vector(to_unsigned(76,8) ,
16414	 => std_logic_vector(to_unsigned(46,8) ,
16415	 => std_logic_vector(to_unsigned(30,8) ,
16416	 => std_logic_vector(to_unsigned(32,8) ,
16417	 => std_logic_vector(to_unsigned(58,8) ,
16418	 => std_logic_vector(to_unsigned(109,8) ,
16419	 => std_logic_vector(to_unsigned(170,8) ,
16420	 => std_logic_vector(to_unsigned(175,8) ,
16421	 => std_logic_vector(to_unsigned(157,8) ,
16422	 => std_logic_vector(to_unsigned(164,8) ,
16423	 => std_logic_vector(to_unsigned(164,8) ,
16424	 => std_logic_vector(to_unsigned(154,8) ,
16425	 => std_logic_vector(to_unsigned(161,8) ,
16426	 => std_logic_vector(to_unsigned(154,8) ,
16427	 => std_logic_vector(to_unsigned(144,8) ,
16428	 => std_logic_vector(to_unsigned(146,8) ,
16429	 => std_logic_vector(to_unsigned(154,8) ,
16430	 => std_logic_vector(to_unsigned(149,8) ,
16431	 => std_logic_vector(to_unsigned(131,8) ,
16432	 => std_logic_vector(to_unsigned(141,8) ,
16433	 => std_logic_vector(to_unsigned(149,8) ,
16434	 => std_logic_vector(to_unsigned(125,8) ,
16435	 => std_logic_vector(to_unsigned(99,8) ,
16436	 => std_logic_vector(to_unsigned(95,8) ,
16437	 => std_logic_vector(to_unsigned(103,8) ,
16438	 => std_logic_vector(to_unsigned(116,8) ,
16439	 => std_logic_vector(to_unsigned(121,8) ,
16440	 => std_logic_vector(to_unsigned(111,8) ,
16441	 => std_logic_vector(to_unsigned(122,8) ,
16442	 => std_logic_vector(to_unsigned(116,8) ,
16443	 => std_logic_vector(to_unsigned(114,8) ,
16444	 => std_logic_vector(to_unsigned(100,8) ,
16445	 => std_logic_vector(to_unsigned(99,8) ,
16446	 => std_logic_vector(to_unsigned(99,8) ,
16447	 => std_logic_vector(to_unsigned(114,8) ,
16448	 => std_logic_vector(to_unsigned(128,8) ,
16449	 => std_logic_vector(to_unsigned(121,8) ,
16450	 => std_logic_vector(to_unsigned(116,8) ,
16451	 => std_logic_vector(to_unsigned(107,8) ,
16452	 => std_logic_vector(to_unsigned(109,8) ,
16453	 => std_logic_vector(to_unsigned(107,8) ,
16454	 => std_logic_vector(to_unsigned(119,8) ,
16455	 => std_logic_vector(to_unsigned(130,8) ,
16456	 => std_logic_vector(to_unsigned(133,8) ,
16457	 => std_logic_vector(to_unsigned(139,8) ,
16458	 => std_logic_vector(to_unsigned(136,8) ,
16459	 => std_logic_vector(to_unsigned(124,8) ,
16460	 => std_logic_vector(to_unsigned(111,8) ,
16461	 => std_logic_vector(to_unsigned(105,8) ,
16462	 => std_logic_vector(to_unsigned(111,8) ,
16463	 => std_logic_vector(to_unsigned(116,8) ,
16464	 => std_logic_vector(to_unsigned(119,8) ,
16465	 => std_logic_vector(to_unsigned(127,8) ,
16466	 => std_logic_vector(to_unsigned(97,8) ,
16467	 => std_logic_vector(to_unsigned(68,8) ,
16468	 => std_logic_vector(to_unsigned(63,8) ,
16469	 => std_logic_vector(to_unsigned(69,8) ,
16470	 => std_logic_vector(to_unsigned(60,8) ,
16471	 => std_logic_vector(to_unsigned(60,8) ,
16472	 => std_logic_vector(to_unsigned(65,8) ,
16473	 => std_logic_vector(to_unsigned(60,8) ,
16474	 => std_logic_vector(to_unsigned(108,8) ,
16475	 => std_logic_vector(to_unsigned(112,8) ,
16476	 => std_logic_vector(to_unsigned(104,8) ,
16477	 => std_logic_vector(to_unsigned(99,8) ,
16478	 => std_logic_vector(to_unsigned(100,8) ,
16479	 => std_logic_vector(to_unsigned(91,8) ,
16480	 => std_logic_vector(to_unsigned(86,8) ,
16481	 => std_logic_vector(to_unsigned(92,8) ,
16482	 => std_logic_vector(to_unsigned(95,8) ,
16483	 => std_logic_vector(to_unsigned(107,8) ,
16484	 => std_logic_vector(to_unsigned(104,8) ,
16485	 => std_logic_vector(to_unsigned(100,8) ,
16486	 => std_logic_vector(to_unsigned(92,8) ,
16487	 => std_logic_vector(to_unsigned(87,8) ,
16488	 => std_logic_vector(to_unsigned(88,8) ,
16489	 => std_logic_vector(to_unsigned(97,8) ,
16490	 => std_logic_vector(to_unsigned(92,8) ,
16491	 => std_logic_vector(to_unsigned(104,8) ,
16492	 => std_logic_vector(to_unsigned(79,8) ,
16493	 => std_logic_vector(to_unsigned(78,8) ,
16494	 => std_logic_vector(to_unsigned(92,8) ,
16495	 => std_logic_vector(to_unsigned(88,8) ,
16496	 => std_logic_vector(to_unsigned(97,8) ,
16497	 => std_logic_vector(to_unsigned(90,8) ,
16498	 => std_logic_vector(to_unsigned(92,8) ,
16499	 => std_logic_vector(to_unsigned(101,8) ,
16500	 => std_logic_vector(to_unsigned(104,8) ,
16501	 => std_logic_vector(to_unsigned(109,8) ,
16502	 => std_logic_vector(to_unsigned(104,8) ,
16503	 => std_logic_vector(to_unsigned(101,8) ,
16504	 => std_logic_vector(to_unsigned(67,8) ,
16505	 => std_logic_vector(to_unsigned(66,8) ,
16506	 => std_logic_vector(to_unsigned(82,8) ,
16507	 => std_logic_vector(to_unsigned(87,8) ,
16508	 => std_logic_vector(to_unsigned(79,8) ,
16509	 => std_logic_vector(to_unsigned(77,8) ,
16510	 => std_logic_vector(to_unsigned(77,8) ,
16511	 => std_logic_vector(to_unsigned(99,8) ,
16512	 => std_logic_vector(to_unsigned(112,8) ,
16513	 => std_logic_vector(to_unsigned(119,8) ,
16514	 => std_logic_vector(to_unsigned(131,8) ,
16515	 => std_logic_vector(to_unsigned(121,8) ,
16516	 => std_logic_vector(to_unsigned(116,8) ,
16517	 => std_logic_vector(to_unsigned(127,8) ,
16518	 => std_logic_vector(to_unsigned(111,8) ,
16519	 => std_logic_vector(to_unsigned(121,8) ,
16520	 => std_logic_vector(to_unsigned(127,8) ,
16521	 => std_logic_vector(to_unsigned(108,8) ,
16522	 => std_logic_vector(to_unsigned(107,8) ,
16523	 => std_logic_vector(to_unsigned(111,8) ,
16524	 => std_logic_vector(to_unsigned(107,8) ,
16525	 => std_logic_vector(to_unsigned(99,8) ,
16526	 => std_logic_vector(to_unsigned(97,8) ,
16527	 => std_logic_vector(to_unsigned(105,8) ,
16528	 => std_logic_vector(to_unsigned(82,8) ,
16529	 => std_logic_vector(to_unsigned(79,8) ,
16530	 => std_logic_vector(to_unsigned(77,8) ,
16531	 => std_logic_vector(to_unsigned(68,8) ,
16532	 => std_logic_vector(to_unsigned(60,8) ,
16533	 => std_logic_vector(to_unsigned(59,8) ,
16534	 => std_logic_vector(to_unsigned(55,8) ,
16535	 => std_logic_vector(to_unsigned(42,8) ,
16536	 => std_logic_vector(to_unsigned(41,8) ,
16537	 => std_logic_vector(to_unsigned(45,8) ,
16538	 => std_logic_vector(to_unsigned(51,8) ,
16539	 => std_logic_vector(to_unsigned(60,8) ,
16540	 => std_logic_vector(to_unsigned(60,8) ,
16541	 => std_logic_vector(to_unsigned(59,8) ,
16542	 => std_logic_vector(to_unsigned(70,8) ,
16543	 => std_logic_vector(to_unsigned(67,8) ,
16544	 => std_logic_vector(to_unsigned(59,8) ,
16545	 => std_logic_vector(to_unsigned(63,8) ,
16546	 => std_logic_vector(to_unsigned(70,8) ,
16547	 => std_logic_vector(to_unsigned(70,8) ,
16548	 => std_logic_vector(to_unsigned(71,8) ,
16549	 => std_logic_vector(to_unsigned(76,8) ,
16550	 => std_logic_vector(to_unsigned(61,8) ,
16551	 => std_logic_vector(to_unsigned(54,8) ,
16552	 => std_logic_vector(to_unsigned(59,8) ,
16553	 => std_logic_vector(to_unsigned(56,8) ,
16554	 => std_logic_vector(to_unsigned(65,8) ,
16555	 => std_logic_vector(to_unsigned(68,8) ,
16556	 => std_logic_vector(to_unsigned(62,8) ,
16557	 => std_logic_vector(to_unsigned(55,8) ,
16558	 => std_logic_vector(to_unsigned(67,8) ,
16559	 => std_logic_vector(to_unsigned(72,8) ,
16560	 => std_logic_vector(to_unsigned(67,8) ,
16561	 => std_logic_vector(to_unsigned(67,8) ,
16562	 => std_logic_vector(to_unsigned(71,8) ,
16563	 => std_logic_vector(to_unsigned(80,8) ,
16564	 => std_logic_vector(to_unsigned(73,8) ,
16565	 => std_logic_vector(to_unsigned(69,8) ,
16566	 => std_logic_vector(to_unsigned(66,8) ,
16567	 => std_logic_vector(to_unsigned(64,8) ,
16568	 => std_logic_vector(to_unsigned(8,8) ,
16569	 => std_logic_vector(to_unsigned(0,8) ,
16570	 => std_logic_vector(to_unsigned(0,8) ,
16571	 => std_logic_vector(to_unsigned(11,8) ,
16572	 => std_logic_vector(to_unsigned(71,8) ,
16573	 => std_logic_vector(to_unsigned(70,8) ,
16574	 => std_logic_vector(to_unsigned(81,8) ,
16575	 => std_logic_vector(to_unsigned(74,8) ,
16576	 => std_logic_vector(to_unsigned(71,8) ,
16577	 => std_logic_vector(to_unsigned(77,8) ,
16578	 => std_logic_vector(to_unsigned(81,8) ,
16579	 => std_logic_vector(to_unsigned(81,8) ,
16580	 => std_logic_vector(to_unsigned(79,8) ,
16581	 => std_logic_vector(to_unsigned(73,8) ,
16582	 => std_logic_vector(to_unsigned(71,8) ,
16583	 => std_logic_vector(to_unsigned(81,8) ,
16584	 => std_logic_vector(to_unsigned(88,8) ,
16585	 => std_logic_vector(to_unsigned(86,8) ,
16586	 => std_logic_vector(to_unsigned(86,8) ,
16587	 => std_logic_vector(to_unsigned(81,8) ,
16588	 => std_logic_vector(to_unsigned(79,8) ,
16589	 => std_logic_vector(to_unsigned(93,8) ,
16590	 => std_logic_vector(to_unsigned(88,8) ,
16591	 => std_logic_vector(to_unsigned(71,8) ,
16592	 => std_logic_vector(to_unsigned(64,8) ,
16593	 => std_logic_vector(to_unsigned(70,8) ,
16594	 => std_logic_vector(to_unsigned(65,8) ,
16595	 => std_logic_vector(to_unsigned(64,8) ,
16596	 => std_logic_vector(to_unsigned(72,8) ,
16597	 => std_logic_vector(to_unsigned(74,8) ,
16598	 => std_logic_vector(to_unsigned(69,8) ,
16599	 => std_logic_vector(to_unsigned(65,8) ,
16600	 => std_logic_vector(to_unsigned(73,8) ,
16601	 => std_logic_vector(to_unsigned(74,8) ,
16602	 => std_logic_vector(to_unsigned(73,8) ,
16603	 => std_logic_vector(to_unsigned(76,8) ,
16604	 => std_logic_vector(to_unsigned(73,8) ,
16605	 => std_logic_vector(to_unsigned(76,8) ,
16606	 => std_logic_vector(to_unsigned(79,8) ,
16607	 => std_logic_vector(to_unsigned(74,8) ,
16608	 => std_logic_vector(to_unsigned(76,8) ,
16609	 => std_logic_vector(to_unsigned(77,8) ,
16610	 => std_logic_vector(to_unsigned(73,8) ,
16611	 => std_logic_vector(to_unsigned(79,8) ,
16612	 => std_logic_vector(to_unsigned(73,8) ,
16613	 => std_logic_vector(to_unsigned(73,8) ,
16614	 => std_logic_vector(to_unsigned(77,8) ,
16615	 => std_logic_vector(to_unsigned(80,8) ,
16616	 => std_logic_vector(to_unsigned(79,8) ,
16617	 => std_logic_vector(to_unsigned(86,8) ,
16618	 => std_logic_vector(to_unsigned(90,8) ,
16619	 => std_logic_vector(to_unsigned(84,8) ,
16620	 => std_logic_vector(to_unsigned(73,8) ,
16621	 => std_logic_vector(to_unsigned(79,8) ,
16622	 => std_logic_vector(to_unsigned(80,8) ,
16623	 => std_logic_vector(to_unsigned(82,8) ,
16624	 => std_logic_vector(to_unsigned(86,8) ,
16625	 => std_logic_vector(to_unsigned(87,8) ,
16626	 => std_logic_vector(to_unsigned(91,8) ,
16627	 => std_logic_vector(to_unsigned(88,8) ,
16628	 => std_logic_vector(to_unsigned(82,8) ,
16629	 => std_logic_vector(to_unsigned(82,8) ,
16630	 => std_logic_vector(to_unsigned(85,8) ,
16631	 => std_logic_vector(to_unsigned(90,8) ,
16632	 => std_logic_vector(to_unsigned(88,8) ,
16633	 => std_logic_vector(to_unsigned(81,8) ,
16634	 => std_logic_vector(to_unsigned(77,8) ,
16635	 => std_logic_vector(to_unsigned(84,8) ,
16636	 => std_logic_vector(to_unsigned(85,8) ,
16637	 => std_logic_vector(to_unsigned(80,8) ,
16638	 => std_logic_vector(to_unsigned(86,8) ,
16639	 => std_logic_vector(to_unsigned(88,8) ,
16640	 => std_logic_vector(to_unsigned(84,8) ,
16641	 => std_logic_vector(to_unsigned(156,8) ,
16642	 => std_logic_vector(to_unsigned(152,8) ,
16643	 => std_logic_vector(to_unsigned(147,8) ,
16644	 => std_logic_vector(to_unsigned(151,8) ,
16645	 => std_logic_vector(to_unsigned(156,8) ,
16646	 => std_logic_vector(to_unsigned(151,8) ,
16647	 => std_logic_vector(to_unsigned(152,8) ,
16648	 => std_logic_vector(to_unsigned(157,8) ,
16649	 => std_logic_vector(to_unsigned(156,8) ,
16650	 => std_logic_vector(to_unsigned(157,8) ,
16651	 => std_logic_vector(to_unsigned(161,8) ,
16652	 => std_logic_vector(to_unsigned(163,8) ,
16653	 => std_logic_vector(to_unsigned(161,8) ,
16654	 => std_logic_vector(to_unsigned(157,8) ,
16655	 => std_logic_vector(to_unsigned(156,8) ,
16656	 => std_logic_vector(to_unsigned(154,8) ,
16657	 => std_logic_vector(to_unsigned(154,8) ,
16658	 => std_logic_vector(to_unsigned(149,8) ,
16659	 => std_logic_vector(to_unsigned(151,8) ,
16660	 => std_logic_vector(to_unsigned(156,8) ,
16661	 => std_logic_vector(to_unsigned(151,8) ,
16662	 => std_logic_vector(to_unsigned(152,8) ,
16663	 => std_logic_vector(to_unsigned(159,8) ,
16664	 => std_logic_vector(to_unsigned(161,8) ,
16665	 => std_logic_vector(to_unsigned(157,8) ,
16666	 => std_logic_vector(to_unsigned(154,8) ,
16667	 => std_logic_vector(to_unsigned(154,8) ,
16668	 => std_logic_vector(to_unsigned(152,8) ,
16669	 => std_logic_vector(to_unsigned(156,8) ,
16670	 => std_logic_vector(to_unsigned(139,8) ,
16671	 => std_logic_vector(to_unsigned(131,8) ,
16672	 => std_logic_vector(to_unsigned(146,8) ,
16673	 => std_logic_vector(to_unsigned(142,8) ,
16674	 => std_logic_vector(to_unsigned(138,8) ,
16675	 => std_logic_vector(to_unsigned(136,8) ,
16676	 => std_logic_vector(to_unsigned(133,8) ,
16677	 => std_logic_vector(to_unsigned(139,8) ,
16678	 => std_logic_vector(to_unsigned(141,8) ,
16679	 => std_logic_vector(to_unsigned(139,8) ,
16680	 => std_logic_vector(to_unsigned(138,8) ,
16681	 => std_logic_vector(to_unsigned(138,8) ,
16682	 => std_logic_vector(to_unsigned(142,8) ,
16683	 => std_logic_vector(to_unsigned(138,8) ,
16684	 => std_logic_vector(to_unsigned(141,8) ,
16685	 => std_logic_vector(to_unsigned(159,8) ,
16686	 => std_logic_vector(to_unsigned(157,8) ,
16687	 => std_logic_vector(to_unsigned(149,8) ,
16688	 => std_logic_vector(to_unsigned(146,8) ,
16689	 => std_logic_vector(to_unsigned(147,8) ,
16690	 => std_logic_vector(to_unsigned(152,8) ,
16691	 => std_logic_vector(to_unsigned(159,8) ,
16692	 => std_logic_vector(to_unsigned(156,8) ,
16693	 => std_logic_vector(to_unsigned(152,8) ,
16694	 => std_logic_vector(to_unsigned(154,8) ,
16695	 => std_logic_vector(to_unsigned(163,8) ,
16696	 => std_logic_vector(to_unsigned(164,8) ,
16697	 => std_logic_vector(to_unsigned(164,8) ,
16698	 => std_logic_vector(to_unsigned(179,8) ,
16699	 => std_logic_vector(to_unsigned(181,8) ,
16700	 => std_logic_vector(to_unsigned(175,8) ,
16701	 => std_logic_vector(to_unsigned(136,8) ,
16702	 => std_logic_vector(to_unsigned(118,8) ,
16703	 => std_logic_vector(to_unsigned(131,8) ,
16704	 => std_logic_vector(to_unsigned(149,8) ,
16705	 => std_logic_vector(to_unsigned(146,8) ,
16706	 => std_logic_vector(to_unsigned(136,8) ,
16707	 => std_logic_vector(to_unsigned(144,8) ,
16708	 => std_logic_vector(to_unsigned(141,8) ,
16709	 => std_logic_vector(to_unsigned(134,8) ,
16710	 => std_logic_vector(to_unsigned(122,8) ,
16711	 => std_logic_vector(to_unsigned(139,8) ,
16712	 => std_logic_vector(to_unsigned(152,8) ,
16713	 => std_logic_vector(to_unsigned(157,8) ,
16714	 => std_logic_vector(to_unsigned(141,8) ,
16715	 => std_logic_vector(to_unsigned(139,8) ,
16716	 => std_logic_vector(to_unsigned(154,8) ,
16717	 => std_logic_vector(to_unsigned(152,8) ,
16718	 => std_logic_vector(to_unsigned(147,8) ,
16719	 => std_logic_vector(to_unsigned(127,8) ,
16720	 => std_logic_vector(to_unsigned(128,8) ,
16721	 => std_logic_vector(to_unsigned(131,8) ,
16722	 => std_logic_vector(to_unsigned(121,8) ,
16723	 => std_logic_vector(to_unsigned(138,8) ,
16724	 => std_logic_vector(to_unsigned(156,8) ,
16725	 => std_logic_vector(to_unsigned(159,8) ,
16726	 => std_logic_vector(to_unsigned(159,8) ,
16727	 => std_logic_vector(to_unsigned(161,8) ,
16728	 => std_logic_vector(to_unsigned(161,8) ,
16729	 => std_logic_vector(to_unsigned(168,8) ,
16730	 => std_logic_vector(to_unsigned(173,8) ,
16731	 => std_logic_vector(to_unsigned(84,8) ,
16732	 => std_logic_vector(to_unsigned(14,8) ,
16733	 => std_logic_vector(to_unsigned(1,8) ,
16734	 => std_logic_vector(to_unsigned(1,8) ,
16735	 => std_logic_vector(to_unsigned(0,8) ,
16736	 => std_logic_vector(to_unsigned(0,8) ,
16737	 => std_logic_vector(to_unsigned(1,8) ,
16738	 => std_logic_vector(to_unsigned(4,8) ,
16739	 => std_logic_vector(to_unsigned(25,8) ,
16740	 => std_logic_vector(to_unsigned(112,8) ,
16741	 => std_logic_vector(to_unsigned(188,8) ,
16742	 => std_logic_vector(to_unsigned(170,8) ,
16743	 => std_logic_vector(to_unsigned(161,8) ,
16744	 => std_logic_vector(to_unsigned(164,8) ,
16745	 => std_logic_vector(to_unsigned(164,8) ,
16746	 => std_logic_vector(to_unsigned(163,8) ,
16747	 => std_logic_vector(to_unsigned(163,8) ,
16748	 => std_logic_vector(to_unsigned(156,8) ,
16749	 => std_logic_vector(to_unsigned(156,8) ,
16750	 => std_logic_vector(to_unsigned(144,8) ,
16751	 => std_logic_vector(to_unsigned(144,8) ,
16752	 => std_logic_vector(to_unsigned(163,8) ,
16753	 => std_logic_vector(to_unsigned(170,8) ,
16754	 => std_logic_vector(to_unsigned(149,8) ,
16755	 => std_logic_vector(to_unsigned(118,8) ,
16756	 => std_logic_vector(to_unsigned(111,8) ,
16757	 => std_logic_vector(to_unsigned(107,8) ,
16758	 => std_logic_vector(to_unsigned(116,8) ,
16759	 => std_logic_vector(to_unsigned(127,8) ,
16760	 => std_logic_vector(to_unsigned(108,8) ,
16761	 => std_logic_vector(to_unsigned(118,8) ,
16762	 => std_logic_vector(to_unsigned(107,8) ,
16763	 => std_logic_vector(to_unsigned(116,8) ,
16764	 => std_logic_vector(to_unsigned(116,8) ,
16765	 => std_logic_vector(to_unsigned(116,8) ,
16766	 => std_logic_vector(to_unsigned(105,8) ,
16767	 => std_logic_vector(to_unsigned(116,8) ,
16768	 => std_logic_vector(to_unsigned(133,8) ,
16769	 => std_logic_vector(to_unsigned(119,8) ,
16770	 => std_logic_vector(to_unsigned(115,8) ,
16771	 => std_logic_vector(to_unsigned(111,8) ,
16772	 => std_logic_vector(to_unsigned(108,8) ,
16773	 => std_logic_vector(to_unsigned(111,8) ,
16774	 => std_logic_vector(to_unsigned(125,8) ,
16775	 => std_logic_vector(to_unsigned(139,8) ,
16776	 => std_logic_vector(to_unsigned(144,8) ,
16777	 => std_logic_vector(to_unsigned(146,8) ,
16778	 => std_logic_vector(to_unsigned(142,8) ,
16779	 => std_logic_vector(to_unsigned(139,8) ,
16780	 => std_logic_vector(to_unsigned(142,8) ,
16781	 => std_logic_vector(to_unsigned(133,8) ,
16782	 => std_logic_vector(to_unsigned(118,8) ,
16783	 => std_logic_vector(to_unsigned(125,8) ,
16784	 => std_logic_vector(to_unsigned(121,8) ,
16785	 => std_logic_vector(to_unsigned(124,8) ,
16786	 => std_logic_vector(to_unsigned(114,8) ,
16787	 => std_logic_vector(to_unsigned(90,8) ,
16788	 => std_logic_vector(to_unsigned(79,8) ,
16789	 => std_logic_vector(to_unsigned(95,8) ,
16790	 => std_logic_vector(to_unsigned(87,8) ,
16791	 => std_logic_vector(to_unsigned(68,8) ,
16792	 => std_logic_vector(to_unsigned(77,8) ,
16793	 => std_logic_vector(to_unsigned(88,8) ,
16794	 => std_logic_vector(to_unsigned(101,8) ,
16795	 => std_logic_vector(to_unsigned(105,8) ,
16796	 => std_logic_vector(to_unsigned(99,8) ,
16797	 => std_logic_vector(to_unsigned(96,8) ,
16798	 => std_logic_vector(to_unsigned(90,8) ,
16799	 => std_logic_vector(to_unsigned(81,8) ,
16800	 => std_logic_vector(to_unsigned(80,8) ,
16801	 => std_logic_vector(to_unsigned(79,8) ,
16802	 => std_logic_vector(to_unsigned(85,8) ,
16803	 => std_logic_vector(to_unsigned(90,8) ,
16804	 => std_logic_vector(to_unsigned(96,8) ,
16805	 => std_logic_vector(to_unsigned(104,8) ,
16806	 => std_logic_vector(to_unsigned(100,8) ,
16807	 => std_logic_vector(to_unsigned(93,8) ,
16808	 => std_logic_vector(to_unsigned(93,8) ,
16809	 => std_logic_vector(to_unsigned(115,8) ,
16810	 => std_logic_vector(to_unsigned(109,8) ,
16811	 => std_logic_vector(to_unsigned(118,8) ,
16812	 => std_logic_vector(to_unsigned(93,8) ,
16813	 => std_logic_vector(to_unsigned(104,8) ,
16814	 => std_logic_vector(to_unsigned(115,8) ,
16815	 => std_logic_vector(to_unsigned(88,8) ,
16816	 => std_logic_vector(to_unsigned(93,8) ,
16817	 => std_logic_vector(to_unsigned(99,8) ,
16818	 => std_logic_vector(to_unsigned(97,8) ,
16819	 => std_logic_vector(to_unsigned(108,8) ,
16820	 => std_logic_vector(to_unsigned(115,8) ,
16821	 => std_logic_vector(to_unsigned(116,8) ,
16822	 => std_logic_vector(to_unsigned(114,8) ,
16823	 => std_logic_vector(to_unsigned(108,8) ,
16824	 => std_logic_vector(to_unsigned(74,8) ,
16825	 => std_logic_vector(to_unsigned(69,8) ,
16826	 => std_logic_vector(to_unsigned(81,8) ,
16827	 => std_logic_vector(to_unsigned(90,8) ,
16828	 => std_logic_vector(to_unsigned(90,8) ,
16829	 => std_logic_vector(to_unsigned(88,8) ,
16830	 => std_logic_vector(to_unsigned(93,8) ,
16831	 => std_logic_vector(to_unsigned(109,8) ,
16832	 => std_logic_vector(to_unsigned(119,8) ,
16833	 => std_logic_vector(to_unsigned(127,8) ,
16834	 => std_logic_vector(to_unsigned(131,8) ,
16835	 => std_logic_vector(to_unsigned(116,8) ,
16836	 => std_logic_vector(to_unsigned(112,8) ,
16837	 => std_logic_vector(to_unsigned(121,8) ,
16838	 => std_logic_vector(to_unsigned(112,8) ,
16839	 => std_logic_vector(to_unsigned(121,8) ,
16840	 => std_logic_vector(to_unsigned(130,8) ,
16841	 => std_logic_vector(to_unsigned(122,8) ,
16842	 => std_logic_vector(to_unsigned(119,8) ,
16843	 => std_logic_vector(to_unsigned(124,8) ,
16844	 => std_logic_vector(to_unsigned(121,8) ,
16845	 => std_logic_vector(to_unsigned(115,8) ,
16846	 => std_logic_vector(to_unsigned(105,8) ,
16847	 => std_logic_vector(to_unsigned(84,8) ,
16848	 => std_logic_vector(to_unsigned(85,8) ,
16849	 => std_logic_vector(to_unsigned(82,8) ,
16850	 => std_logic_vector(to_unsigned(68,8) ,
16851	 => std_logic_vector(to_unsigned(44,8) ,
16852	 => std_logic_vector(to_unsigned(45,8) ,
16853	 => std_logic_vector(to_unsigned(51,8) ,
16854	 => std_logic_vector(to_unsigned(46,8) ,
16855	 => std_logic_vector(to_unsigned(47,8) ,
16856	 => std_logic_vector(to_unsigned(46,8) ,
16857	 => std_logic_vector(to_unsigned(56,8) ,
16858	 => std_logic_vector(to_unsigned(65,8) ,
16859	 => std_logic_vector(to_unsigned(66,8) ,
16860	 => std_logic_vector(to_unsigned(68,8) ,
16861	 => std_logic_vector(to_unsigned(65,8) ,
16862	 => std_logic_vector(to_unsigned(74,8) ,
16863	 => std_logic_vector(to_unsigned(66,8) ,
16864	 => std_logic_vector(to_unsigned(53,8) ,
16865	 => std_logic_vector(to_unsigned(58,8) ,
16866	 => std_logic_vector(to_unsigned(73,8) ,
16867	 => std_logic_vector(to_unsigned(77,8) ,
16868	 => std_logic_vector(to_unsigned(67,8) ,
16869	 => std_logic_vector(to_unsigned(70,8) ,
16870	 => std_logic_vector(to_unsigned(63,8) ,
16871	 => std_logic_vector(to_unsigned(51,8) ,
16872	 => std_logic_vector(to_unsigned(55,8) ,
16873	 => std_logic_vector(to_unsigned(56,8) ,
16874	 => std_logic_vector(to_unsigned(62,8) ,
16875	 => std_logic_vector(to_unsigned(67,8) ,
16876	 => std_logic_vector(to_unsigned(62,8) ,
16877	 => std_logic_vector(to_unsigned(59,8) ,
16878	 => std_logic_vector(to_unsigned(71,8) ,
16879	 => std_logic_vector(to_unsigned(73,8) ,
16880	 => std_logic_vector(to_unsigned(67,8) ,
16881	 => std_logic_vector(to_unsigned(72,8) ,
16882	 => std_logic_vector(to_unsigned(73,8) ,
16883	 => std_logic_vector(to_unsigned(74,8) ,
16884	 => std_logic_vector(to_unsigned(80,8) ,
16885	 => std_logic_vector(to_unsigned(71,8) ,
16886	 => std_logic_vector(to_unsigned(68,8) ,
16887	 => std_logic_vector(to_unsigned(68,8) ,
16888	 => std_logic_vector(to_unsigned(21,8) ,
16889	 => std_logic_vector(to_unsigned(1,8) ,
16890	 => std_logic_vector(to_unsigned(0,8) ,
16891	 => std_logic_vector(to_unsigned(5,8) ,
16892	 => std_logic_vector(to_unsigned(73,8) ,
16893	 => std_logic_vector(to_unsigned(82,8) ,
16894	 => std_logic_vector(to_unsigned(71,8) ,
16895	 => std_logic_vector(to_unsigned(78,8) ,
16896	 => std_logic_vector(to_unsigned(81,8) ,
16897	 => std_logic_vector(to_unsigned(77,8) ,
16898	 => std_logic_vector(to_unsigned(73,8) ,
16899	 => std_logic_vector(to_unsigned(85,8) ,
16900	 => std_logic_vector(to_unsigned(88,8) ,
16901	 => std_logic_vector(to_unsigned(77,8) ,
16902	 => std_logic_vector(to_unsigned(84,8) ,
16903	 => std_logic_vector(to_unsigned(81,8) ,
16904	 => std_logic_vector(to_unsigned(72,8) ,
16905	 => std_logic_vector(to_unsigned(84,8) ,
16906	 => std_logic_vector(to_unsigned(86,8) ,
16907	 => std_logic_vector(to_unsigned(81,8) ,
16908	 => std_logic_vector(to_unsigned(81,8) ,
16909	 => std_logic_vector(to_unsigned(88,8) ,
16910	 => std_logic_vector(to_unsigned(87,8) ,
16911	 => std_logic_vector(to_unsigned(72,8) ,
16912	 => std_logic_vector(to_unsigned(76,8) ,
16913	 => std_logic_vector(to_unsigned(78,8) ,
16914	 => std_logic_vector(to_unsigned(65,8) ,
16915	 => std_logic_vector(to_unsigned(63,8) ,
16916	 => std_logic_vector(to_unsigned(66,8) ,
16917	 => std_logic_vector(to_unsigned(78,8) ,
16918	 => std_logic_vector(to_unsigned(71,8) ,
16919	 => std_logic_vector(to_unsigned(61,8) ,
16920	 => std_logic_vector(to_unsigned(65,8) ,
16921	 => std_logic_vector(to_unsigned(66,8) ,
16922	 => std_logic_vector(to_unsigned(69,8) ,
16923	 => std_logic_vector(to_unsigned(74,8) ,
16924	 => std_logic_vector(to_unsigned(72,8) ,
16925	 => std_logic_vector(to_unsigned(72,8) ,
16926	 => std_logic_vector(to_unsigned(74,8) ,
16927	 => std_logic_vector(to_unsigned(71,8) ,
16928	 => std_logic_vector(to_unsigned(76,8) ,
16929	 => std_logic_vector(to_unsigned(84,8) ,
16930	 => std_logic_vector(to_unsigned(77,8) ,
16931	 => std_logic_vector(to_unsigned(73,8) ,
16932	 => std_logic_vector(to_unsigned(67,8) ,
16933	 => std_logic_vector(to_unsigned(74,8) ,
16934	 => std_logic_vector(to_unsigned(77,8) ,
16935	 => std_logic_vector(to_unsigned(70,8) ,
16936	 => std_logic_vector(to_unsigned(78,8) ,
16937	 => std_logic_vector(to_unsigned(73,8) ,
16938	 => std_logic_vector(to_unsigned(68,8) ,
16939	 => std_logic_vector(to_unsigned(70,8) ,
16940	 => std_logic_vector(to_unsigned(74,8) ,
16941	 => std_logic_vector(to_unsigned(81,8) ,
16942	 => std_logic_vector(to_unsigned(79,8) ,
16943	 => std_logic_vector(to_unsigned(88,8) ,
16944	 => std_logic_vector(to_unsigned(82,8) ,
16945	 => std_logic_vector(to_unsigned(85,8) ,
16946	 => std_logic_vector(to_unsigned(93,8) ,
16947	 => std_logic_vector(to_unsigned(91,8) ,
16948	 => std_logic_vector(to_unsigned(82,8) ,
16949	 => std_logic_vector(to_unsigned(78,8) ,
16950	 => std_logic_vector(to_unsigned(74,8) ,
16951	 => std_logic_vector(to_unsigned(86,8) ,
16952	 => std_logic_vector(to_unsigned(77,8) ,
16953	 => std_logic_vector(to_unsigned(68,8) ,
16954	 => std_logic_vector(to_unsigned(68,8) ,
16955	 => std_logic_vector(to_unsigned(74,8) ,
16956	 => std_logic_vector(to_unsigned(80,8) ,
16957	 => std_logic_vector(to_unsigned(78,8) ,
16958	 => std_logic_vector(to_unsigned(84,8) ,
16959	 => std_logic_vector(to_unsigned(90,8) ,
16960	 => std_logic_vector(to_unsigned(88,8) ,
16961	 => std_logic_vector(to_unsigned(144,8) ,
16962	 => std_logic_vector(to_unsigned(157,8) ,
16963	 => std_logic_vector(to_unsigned(152,8) ,
16964	 => std_logic_vector(to_unsigned(147,8) ,
16965	 => std_logic_vector(to_unsigned(154,8) ,
16966	 => std_logic_vector(to_unsigned(156,8) ,
16967	 => std_logic_vector(to_unsigned(157,8) ,
16968	 => std_logic_vector(to_unsigned(159,8) ,
16969	 => std_logic_vector(to_unsigned(161,8) ,
16970	 => std_logic_vector(to_unsigned(157,8) ,
16971	 => std_logic_vector(to_unsigned(157,8) ,
16972	 => std_logic_vector(to_unsigned(163,8) ,
16973	 => std_logic_vector(to_unsigned(159,8) ,
16974	 => std_logic_vector(to_unsigned(154,8) ,
16975	 => std_logic_vector(to_unsigned(151,8) ,
16976	 => std_logic_vector(to_unsigned(149,8) ,
16977	 => std_logic_vector(to_unsigned(151,8) ,
16978	 => std_logic_vector(to_unsigned(151,8) ,
16979	 => std_logic_vector(to_unsigned(149,8) ,
16980	 => std_logic_vector(to_unsigned(152,8) ,
16981	 => std_logic_vector(to_unsigned(151,8) ,
16982	 => std_logic_vector(to_unsigned(152,8) ,
16983	 => std_logic_vector(to_unsigned(157,8) ,
16984	 => std_logic_vector(to_unsigned(157,8) ,
16985	 => std_logic_vector(to_unsigned(161,8) ,
16986	 => std_logic_vector(to_unsigned(159,8) ,
16987	 => std_logic_vector(to_unsigned(154,8) ,
16988	 => std_logic_vector(to_unsigned(152,8) ,
16989	 => std_logic_vector(to_unsigned(151,8) ,
16990	 => std_logic_vector(to_unsigned(156,8) ,
16991	 => std_logic_vector(to_unsigned(146,8) ,
16992	 => std_logic_vector(to_unsigned(76,8) ,
16993	 => std_logic_vector(to_unsigned(69,8) ,
16994	 => std_logic_vector(to_unsigned(131,8) ,
16995	 => std_logic_vector(to_unsigned(151,8) ,
16996	 => std_logic_vector(to_unsigned(139,8) ,
16997	 => std_logic_vector(to_unsigned(151,8) ,
16998	 => std_logic_vector(to_unsigned(147,8) ,
16999	 => std_logic_vector(to_unsigned(147,8) ,
17000	 => std_logic_vector(to_unsigned(147,8) ,
17001	 => std_logic_vector(to_unsigned(149,8) ,
17002	 => std_logic_vector(to_unsigned(152,8) ,
17003	 => std_logic_vector(to_unsigned(149,8) ,
17004	 => std_logic_vector(to_unsigned(149,8) ,
17005	 => std_logic_vector(to_unsigned(152,8) ,
17006	 => std_logic_vector(to_unsigned(156,8) ,
17007	 => std_logic_vector(to_unsigned(149,8) ,
17008	 => std_logic_vector(to_unsigned(144,8) ,
17009	 => std_logic_vector(to_unsigned(142,8) ,
17010	 => std_logic_vector(to_unsigned(151,8) ,
17011	 => std_logic_vector(to_unsigned(156,8) ,
17012	 => std_logic_vector(to_unsigned(154,8) ,
17013	 => std_logic_vector(to_unsigned(152,8) ,
17014	 => std_logic_vector(to_unsigned(156,8) ,
17015	 => std_logic_vector(to_unsigned(168,8) ,
17016	 => std_logic_vector(to_unsigned(179,8) ,
17017	 => std_logic_vector(to_unsigned(173,8) ,
17018	 => std_logic_vector(to_unsigned(115,8) ,
17019	 => std_logic_vector(to_unsigned(104,8) ,
17020	 => std_logic_vector(to_unsigned(97,8) ,
17021	 => std_logic_vector(to_unsigned(81,8) ,
17022	 => std_logic_vector(to_unsigned(67,8) ,
17023	 => std_logic_vector(to_unsigned(92,8) ,
17024	 => std_logic_vector(to_unsigned(91,8) ,
17025	 => std_logic_vector(to_unsigned(109,8) ,
17026	 => std_logic_vector(to_unsigned(139,8) ,
17027	 => std_logic_vector(to_unsigned(154,8) ,
17028	 => std_logic_vector(to_unsigned(138,8) ,
17029	 => std_logic_vector(to_unsigned(133,8) ,
17030	 => std_logic_vector(to_unsigned(142,8) ,
17031	 => std_logic_vector(to_unsigned(149,8) ,
17032	 => std_logic_vector(to_unsigned(151,8) ,
17033	 => std_logic_vector(to_unsigned(154,8) ,
17034	 => std_logic_vector(to_unsigned(139,8) ,
17035	 => std_logic_vector(to_unsigned(138,8) ,
17036	 => std_logic_vector(to_unsigned(159,8) ,
17037	 => std_logic_vector(to_unsigned(166,8) ,
17038	 => std_logic_vector(to_unsigned(147,8) ,
17039	 => std_logic_vector(to_unsigned(121,8) ,
17040	 => std_logic_vector(to_unsigned(139,8) ,
17041	 => std_logic_vector(to_unsigned(141,8) ,
17042	 => std_logic_vector(to_unsigned(121,8) ,
17043	 => std_logic_vector(to_unsigned(142,8) ,
17044	 => std_logic_vector(to_unsigned(156,8) ,
17045	 => std_logic_vector(to_unsigned(156,8) ,
17046	 => std_logic_vector(to_unsigned(157,8) ,
17047	 => std_logic_vector(to_unsigned(159,8) ,
17048	 => std_logic_vector(to_unsigned(173,8) ,
17049	 => std_logic_vector(to_unsigned(161,8) ,
17050	 => std_logic_vector(to_unsigned(38,8) ,
17051	 => std_logic_vector(to_unsigned(2,8) ,
17052	 => std_logic_vector(to_unsigned(0,8) ,
17053	 => std_logic_vector(to_unsigned(2,8) ,
17054	 => std_logic_vector(to_unsigned(2,8) ,
17055	 => std_logic_vector(to_unsigned(2,8) ,
17056	 => std_logic_vector(to_unsigned(2,8) ,
17057	 => std_logic_vector(to_unsigned(2,8) ,
17058	 => std_logic_vector(to_unsigned(2,8) ,
17059	 => std_logic_vector(to_unsigned(2,8) ,
17060	 => std_logic_vector(to_unsigned(5,8) ,
17061	 => std_logic_vector(to_unsigned(92,8) ,
17062	 => std_logic_vector(to_unsigned(188,8) ,
17063	 => std_logic_vector(to_unsigned(159,8) ,
17064	 => std_logic_vector(to_unsigned(161,8) ,
17065	 => std_logic_vector(to_unsigned(163,8) ,
17066	 => std_logic_vector(to_unsigned(161,8) ,
17067	 => std_logic_vector(to_unsigned(156,8) ,
17068	 => std_logic_vector(to_unsigned(159,8) ,
17069	 => std_logic_vector(to_unsigned(164,8) ,
17070	 => std_logic_vector(to_unsigned(159,8) ,
17071	 => std_logic_vector(to_unsigned(166,8) ,
17072	 => std_logic_vector(to_unsigned(163,8) ,
17073	 => std_logic_vector(to_unsigned(159,8) ,
17074	 => std_logic_vector(to_unsigned(157,8) ,
17075	 => std_logic_vector(to_unsigned(127,8) ,
17076	 => std_logic_vector(to_unsigned(119,8) ,
17077	 => std_logic_vector(to_unsigned(114,8) ,
17078	 => std_logic_vector(to_unsigned(127,8) ,
17079	 => std_logic_vector(to_unsigned(134,8) ,
17080	 => std_logic_vector(to_unsigned(112,8) ,
17081	 => std_logic_vector(to_unsigned(116,8) ,
17082	 => std_logic_vector(to_unsigned(116,8) ,
17083	 => std_logic_vector(to_unsigned(127,8) ,
17084	 => std_logic_vector(to_unsigned(118,8) ,
17085	 => std_logic_vector(to_unsigned(115,8) ,
17086	 => std_logic_vector(to_unsigned(111,8) ,
17087	 => std_logic_vector(to_unsigned(130,8) ,
17088	 => std_logic_vector(to_unsigned(133,8) ,
17089	 => std_logic_vector(to_unsigned(116,8) ,
17090	 => std_logic_vector(to_unsigned(121,8) ,
17091	 => std_logic_vector(to_unsigned(118,8) ,
17092	 => std_logic_vector(to_unsigned(119,8) ,
17093	 => std_logic_vector(to_unsigned(127,8) ,
17094	 => std_logic_vector(to_unsigned(130,8) ,
17095	 => std_logic_vector(to_unsigned(136,8) ,
17096	 => std_logic_vector(to_unsigned(147,8) ,
17097	 => std_logic_vector(to_unsigned(146,8) ,
17098	 => std_logic_vector(to_unsigned(142,8) ,
17099	 => std_logic_vector(to_unsigned(152,8) ,
17100	 => std_logic_vector(to_unsigned(159,8) ,
17101	 => std_logic_vector(to_unsigned(146,8) ,
17102	 => std_logic_vector(to_unsigned(116,8) ,
17103	 => std_logic_vector(to_unsigned(116,8) ,
17104	 => std_logic_vector(to_unsigned(124,8) ,
17105	 => std_logic_vector(to_unsigned(130,8) ,
17106	 => std_logic_vector(to_unsigned(146,8) ,
17107	 => std_logic_vector(to_unsigned(116,8) ,
17108	 => std_logic_vector(to_unsigned(100,8) ,
17109	 => std_logic_vector(to_unsigned(127,8) ,
17110	 => std_logic_vector(to_unsigned(112,8) ,
17111	 => std_logic_vector(to_unsigned(87,8) ,
17112	 => std_logic_vector(to_unsigned(85,8) ,
17113	 => std_logic_vector(to_unsigned(95,8) ,
17114	 => std_logic_vector(to_unsigned(95,8) ,
17115	 => std_logic_vector(to_unsigned(93,8) ,
17116	 => std_logic_vector(to_unsigned(92,8) ,
17117	 => std_logic_vector(to_unsigned(88,8) ,
17118	 => std_logic_vector(to_unsigned(81,8) ,
17119	 => std_logic_vector(to_unsigned(82,8) ,
17120	 => std_logic_vector(to_unsigned(90,8) ,
17121	 => std_logic_vector(to_unsigned(72,8) ,
17122	 => std_logic_vector(to_unsigned(72,8) ,
17123	 => std_logic_vector(to_unsigned(87,8) ,
17124	 => std_logic_vector(to_unsigned(112,8) ,
17125	 => std_logic_vector(to_unsigned(112,8) ,
17126	 => std_logic_vector(to_unsigned(93,8) ,
17127	 => std_logic_vector(to_unsigned(97,8) ,
17128	 => std_logic_vector(to_unsigned(107,8) ,
17129	 => std_logic_vector(to_unsigned(118,8) ,
17130	 => std_logic_vector(to_unsigned(115,8) ,
17131	 => std_logic_vector(to_unsigned(118,8) ,
17132	 => std_logic_vector(to_unsigned(99,8) ,
17133	 => std_logic_vector(to_unsigned(99,8) ,
17134	 => std_logic_vector(to_unsigned(105,8) ,
17135	 => std_logic_vector(to_unsigned(91,8) ,
17136	 => std_logic_vector(to_unsigned(90,8) ,
17137	 => std_logic_vector(to_unsigned(99,8) ,
17138	 => std_logic_vector(to_unsigned(107,8) ,
17139	 => std_logic_vector(to_unsigned(114,8) ,
17140	 => std_logic_vector(to_unsigned(116,8) ,
17141	 => std_logic_vector(to_unsigned(121,8) ,
17142	 => std_logic_vector(to_unsigned(115,8) ,
17143	 => std_logic_vector(to_unsigned(111,8) ,
17144	 => std_logic_vector(to_unsigned(85,8) ,
17145	 => std_logic_vector(to_unsigned(78,8) ,
17146	 => std_logic_vector(to_unsigned(95,8) ,
17147	 => std_logic_vector(to_unsigned(99,8) ,
17148	 => std_logic_vector(to_unsigned(93,8) ,
17149	 => std_logic_vector(to_unsigned(88,8) ,
17150	 => std_logic_vector(to_unsigned(90,8) ,
17151	 => std_logic_vector(to_unsigned(87,8) ,
17152	 => std_logic_vector(to_unsigned(111,8) ,
17153	 => std_logic_vector(to_unsigned(127,8) ,
17154	 => std_logic_vector(to_unsigned(128,8) ,
17155	 => std_logic_vector(to_unsigned(116,8) ,
17156	 => std_logic_vector(to_unsigned(109,8) ,
17157	 => std_logic_vector(to_unsigned(115,8) ,
17158	 => std_logic_vector(to_unsigned(116,8) ,
17159	 => std_logic_vector(to_unsigned(122,8) ,
17160	 => std_logic_vector(to_unsigned(133,8) ,
17161	 => std_logic_vector(to_unsigned(130,8) ,
17162	 => std_logic_vector(to_unsigned(124,8) ,
17163	 => std_logic_vector(to_unsigned(121,8) ,
17164	 => std_logic_vector(to_unsigned(99,8) ,
17165	 => std_logic_vector(to_unsigned(96,8) ,
17166	 => std_logic_vector(to_unsigned(77,8) ,
17167	 => std_logic_vector(to_unsigned(52,8) ,
17168	 => std_logic_vector(to_unsigned(74,8) ,
17169	 => std_logic_vector(to_unsigned(79,8) ,
17170	 => std_logic_vector(to_unsigned(67,8) ,
17171	 => std_logic_vector(to_unsigned(44,8) ,
17172	 => std_logic_vector(to_unsigned(43,8) ,
17173	 => std_logic_vector(to_unsigned(46,8) ,
17174	 => std_logic_vector(to_unsigned(48,8) ,
17175	 => std_logic_vector(to_unsigned(50,8) ,
17176	 => std_logic_vector(to_unsigned(54,8) ,
17177	 => std_logic_vector(to_unsigned(69,8) ,
17178	 => std_logic_vector(to_unsigned(63,8) ,
17179	 => std_logic_vector(to_unsigned(65,8) ,
17180	 => std_logic_vector(to_unsigned(70,8) ,
17181	 => std_logic_vector(to_unsigned(67,8) ,
17182	 => std_logic_vector(to_unsigned(74,8) ,
17183	 => std_logic_vector(to_unsigned(74,8) ,
17184	 => std_logic_vector(to_unsigned(61,8) ,
17185	 => std_logic_vector(to_unsigned(60,8) ,
17186	 => std_logic_vector(to_unsigned(72,8) ,
17187	 => std_logic_vector(to_unsigned(74,8) ,
17188	 => std_logic_vector(to_unsigned(69,8) ,
17189	 => std_logic_vector(to_unsigned(69,8) ,
17190	 => std_logic_vector(to_unsigned(74,8) ,
17191	 => std_logic_vector(to_unsigned(69,8) ,
17192	 => std_logic_vector(to_unsigned(68,8) ,
17193	 => std_logic_vector(to_unsigned(64,8) ,
17194	 => std_logic_vector(to_unsigned(55,8) ,
17195	 => std_logic_vector(to_unsigned(63,8) ,
17196	 => std_logic_vector(to_unsigned(68,8) ,
17197	 => std_logic_vector(to_unsigned(71,8) ,
17198	 => std_logic_vector(to_unsigned(81,8) ,
17199	 => std_logic_vector(to_unsigned(71,8) ,
17200	 => std_logic_vector(to_unsigned(59,8) ,
17201	 => std_logic_vector(to_unsigned(69,8) ,
17202	 => std_logic_vector(to_unsigned(67,8) ,
17203	 => std_logic_vector(to_unsigned(71,8) ,
17204	 => std_logic_vector(to_unsigned(77,8) ,
17205	 => std_logic_vector(to_unsigned(70,8) ,
17206	 => std_logic_vector(to_unsigned(66,8) ,
17207	 => std_logic_vector(to_unsigned(73,8) ,
17208	 => std_logic_vector(to_unsigned(51,8) ,
17209	 => std_logic_vector(to_unsigned(2,8) ,
17210	 => std_logic_vector(to_unsigned(0,8) ,
17211	 => std_logic_vector(to_unsigned(2,8) ,
17212	 => std_logic_vector(to_unsigned(59,8) ,
17213	 => std_logic_vector(to_unsigned(90,8) ,
17214	 => std_logic_vector(to_unsigned(64,8) ,
17215	 => std_logic_vector(to_unsigned(70,8) ,
17216	 => std_logic_vector(to_unsigned(72,8) ,
17217	 => std_logic_vector(to_unsigned(72,8) ,
17218	 => std_logic_vector(to_unsigned(77,8) ,
17219	 => std_logic_vector(to_unsigned(87,8) ,
17220	 => std_logic_vector(to_unsigned(87,8) ,
17221	 => std_logic_vector(to_unsigned(81,8) ,
17222	 => std_logic_vector(to_unsigned(85,8) ,
17223	 => std_logic_vector(to_unsigned(81,8) ,
17224	 => std_logic_vector(to_unsigned(78,8) ,
17225	 => std_logic_vector(to_unsigned(81,8) ,
17226	 => std_logic_vector(to_unsigned(85,8) ,
17227	 => std_logic_vector(to_unsigned(84,8) ,
17228	 => std_logic_vector(to_unsigned(76,8) ,
17229	 => std_logic_vector(to_unsigned(77,8) ,
17230	 => std_logic_vector(to_unsigned(82,8) ,
17231	 => std_logic_vector(to_unsigned(80,8) ,
17232	 => std_logic_vector(to_unsigned(76,8) ,
17233	 => std_logic_vector(to_unsigned(71,8) ,
17234	 => std_logic_vector(to_unsigned(72,8) ,
17235	 => std_logic_vector(to_unsigned(76,8) ,
17236	 => std_logic_vector(to_unsigned(71,8) ,
17237	 => std_logic_vector(to_unsigned(74,8) ,
17238	 => std_logic_vector(to_unsigned(70,8) ,
17239	 => std_logic_vector(to_unsigned(67,8) ,
17240	 => std_logic_vector(to_unsigned(68,8) ,
17241	 => std_logic_vector(to_unsigned(67,8) ,
17242	 => std_logic_vector(to_unsigned(72,8) ,
17243	 => std_logic_vector(to_unsigned(72,8) ,
17244	 => std_logic_vector(to_unsigned(66,8) ,
17245	 => std_logic_vector(to_unsigned(73,8) ,
17246	 => std_logic_vector(to_unsigned(74,8) ,
17247	 => std_logic_vector(to_unsigned(72,8) ,
17248	 => std_logic_vector(to_unsigned(78,8) ,
17249	 => std_logic_vector(to_unsigned(86,8) ,
17250	 => std_logic_vector(to_unsigned(85,8) ,
17251	 => std_logic_vector(to_unsigned(73,8) ,
17252	 => std_logic_vector(to_unsigned(73,8) ,
17253	 => std_logic_vector(to_unsigned(79,8) ,
17254	 => std_logic_vector(to_unsigned(78,8) ,
17255	 => std_logic_vector(to_unsigned(74,8) ,
17256	 => std_logic_vector(to_unsigned(80,8) ,
17257	 => std_logic_vector(to_unsigned(79,8) ,
17258	 => std_logic_vector(to_unsigned(73,8) ,
17259	 => std_logic_vector(to_unsigned(69,8) ,
17260	 => std_logic_vector(to_unsigned(81,8) ,
17261	 => std_logic_vector(to_unsigned(91,8) ,
17262	 => std_logic_vector(to_unsigned(86,8) ,
17263	 => std_logic_vector(to_unsigned(93,8) ,
17264	 => std_logic_vector(to_unsigned(90,8) ,
17265	 => std_logic_vector(to_unsigned(81,8) ,
17266	 => std_logic_vector(to_unsigned(78,8) ,
17267	 => std_logic_vector(to_unsigned(86,8) ,
17268	 => std_logic_vector(to_unsigned(85,8) ,
17269	 => std_logic_vector(to_unsigned(82,8) ,
17270	 => std_logic_vector(to_unsigned(81,8) ,
17271	 => std_logic_vector(to_unsigned(91,8) ,
17272	 => std_logic_vector(to_unsigned(78,8) ,
17273	 => std_logic_vector(to_unsigned(67,8) ,
17274	 => std_logic_vector(to_unsigned(79,8) ,
17275	 => std_logic_vector(to_unsigned(90,8) ,
17276	 => std_logic_vector(to_unsigned(93,8) ,
17277	 => std_logic_vector(to_unsigned(90,8) ,
17278	 => std_logic_vector(to_unsigned(92,8) ,
17279	 => std_logic_vector(to_unsigned(93,8) ,
17280	 => std_logic_vector(to_unsigned(95,8) ,
17281	 => std_logic_vector(to_unsigned(147,8) ,
17282	 => std_logic_vector(to_unsigned(152,8) ,
17283	 => std_logic_vector(to_unsigned(144,8) ,
17284	 => std_logic_vector(to_unsigned(138,8) ,
17285	 => std_logic_vector(to_unsigned(147,8) ,
17286	 => std_logic_vector(to_unsigned(159,8) ,
17287	 => std_logic_vector(to_unsigned(161,8) ,
17288	 => std_logic_vector(to_unsigned(156,8) ,
17289	 => std_logic_vector(to_unsigned(157,8) ,
17290	 => std_logic_vector(to_unsigned(154,8) ,
17291	 => std_logic_vector(to_unsigned(149,8) ,
17292	 => std_logic_vector(to_unsigned(154,8) ,
17293	 => std_logic_vector(to_unsigned(157,8) ,
17294	 => std_logic_vector(to_unsigned(154,8) ,
17295	 => std_logic_vector(to_unsigned(152,8) ,
17296	 => std_logic_vector(to_unsigned(156,8) ,
17297	 => std_logic_vector(to_unsigned(154,8) ,
17298	 => std_logic_vector(to_unsigned(152,8) ,
17299	 => std_logic_vector(to_unsigned(149,8) ,
17300	 => std_logic_vector(to_unsigned(149,8) ,
17301	 => std_logic_vector(to_unsigned(146,8) ,
17302	 => std_logic_vector(to_unsigned(151,8) ,
17303	 => std_logic_vector(to_unsigned(157,8) ,
17304	 => std_logic_vector(to_unsigned(154,8) ,
17305	 => std_logic_vector(to_unsigned(156,8) ,
17306	 => std_logic_vector(to_unsigned(159,8) ,
17307	 => std_logic_vector(to_unsigned(149,8) ,
17308	 => std_logic_vector(to_unsigned(151,8) ,
17309	 => std_logic_vector(to_unsigned(151,8) ,
17310	 => std_logic_vector(to_unsigned(149,8) ,
17311	 => std_logic_vector(to_unsigned(108,8) ,
17312	 => std_logic_vector(to_unsigned(35,8) ,
17313	 => std_logic_vector(to_unsigned(29,8) ,
17314	 => std_logic_vector(to_unsigned(41,8) ,
17315	 => std_logic_vector(to_unsigned(108,8) ,
17316	 => std_logic_vector(to_unsigned(154,8) ,
17317	 => std_logic_vector(to_unsigned(144,8) ,
17318	 => std_logic_vector(to_unsigned(151,8) ,
17319	 => std_logic_vector(to_unsigned(147,8) ,
17320	 => std_logic_vector(to_unsigned(141,8) ,
17321	 => std_logic_vector(to_unsigned(147,8) ,
17322	 => std_logic_vector(to_unsigned(151,8) ,
17323	 => std_logic_vector(to_unsigned(151,8) ,
17324	 => std_logic_vector(to_unsigned(147,8) ,
17325	 => std_logic_vector(to_unsigned(147,8) ,
17326	 => std_logic_vector(to_unsigned(151,8) ,
17327	 => std_logic_vector(to_unsigned(146,8) ,
17328	 => std_logic_vector(to_unsigned(146,8) ,
17329	 => std_logic_vector(to_unsigned(147,8) ,
17330	 => std_logic_vector(to_unsigned(149,8) ,
17331	 => std_logic_vector(to_unsigned(151,8) ,
17332	 => std_logic_vector(to_unsigned(147,8) ,
17333	 => std_logic_vector(to_unsigned(152,8) ,
17334	 => std_logic_vector(to_unsigned(147,8) ,
17335	 => std_logic_vector(to_unsigned(146,8) ,
17336	 => std_logic_vector(to_unsigned(159,8) ,
17337	 => std_logic_vector(to_unsigned(116,8) ,
17338	 => std_logic_vector(to_unsigned(46,8) ,
17339	 => std_logic_vector(to_unsigned(58,8) ,
17340	 => std_logic_vector(to_unsigned(64,8) ,
17341	 => std_logic_vector(to_unsigned(65,8) ,
17342	 => std_logic_vector(to_unsigned(41,8) ,
17343	 => std_logic_vector(to_unsigned(55,8) ,
17344	 => std_logic_vector(to_unsigned(61,8) ,
17345	 => std_logic_vector(to_unsigned(64,8) ,
17346	 => std_logic_vector(to_unsigned(103,8) ,
17347	 => std_logic_vector(to_unsigned(138,8) ,
17348	 => std_logic_vector(to_unsigned(139,8) ,
17349	 => std_logic_vector(to_unsigned(141,8) ,
17350	 => std_logic_vector(to_unsigned(151,8) ,
17351	 => std_logic_vector(to_unsigned(156,8) ,
17352	 => std_logic_vector(to_unsigned(159,8) ,
17353	 => std_logic_vector(to_unsigned(163,8) ,
17354	 => std_logic_vector(to_unsigned(154,8) ,
17355	 => std_logic_vector(to_unsigned(147,8) ,
17356	 => std_logic_vector(to_unsigned(163,8) ,
17357	 => std_logic_vector(to_unsigned(164,8) ,
17358	 => std_logic_vector(to_unsigned(146,8) ,
17359	 => std_logic_vector(to_unsigned(130,8) ,
17360	 => std_logic_vector(to_unsigned(144,8) ,
17361	 => std_logic_vector(to_unsigned(131,8) ,
17362	 => std_logic_vector(to_unsigned(116,8) ,
17363	 => std_logic_vector(to_unsigned(138,8) ,
17364	 => std_logic_vector(to_unsigned(142,8) ,
17365	 => std_logic_vector(to_unsigned(144,8) ,
17366	 => std_logic_vector(to_unsigned(152,8) ,
17367	 => std_logic_vector(to_unsigned(175,8) ,
17368	 => std_logic_vector(to_unsigned(141,8) ,
17369	 => std_logic_vector(to_unsigned(24,8) ,
17370	 => std_logic_vector(to_unsigned(1,8) ,
17371	 => std_logic_vector(to_unsigned(1,8) ,
17372	 => std_logic_vector(to_unsigned(1,8) ,
17373	 => std_logic_vector(to_unsigned(2,8) ,
17374	 => std_logic_vector(to_unsigned(2,8) ,
17375	 => std_logic_vector(to_unsigned(3,8) ,
17376	 => std_logic_vector(to_unsigned(2,8) ,
17377	 => std_logic_vector(to_unsigned(2,8) ,
17378	 => std_logic_vector(to_unsigned(2,8) ,
17379	 => std_logic_vector(to_unsigned(6,8) ,
17380	 => std_logic_vector(to_unsigned(1,8) ,
17381	 => std_logic_vector(to_unsigned(4,8) ,
17382	 => std_logic_vector(to_unsigned(109,8) ,
17383	 => std_logic_vector(to_unsigned(175,8) ,
17384	 => std_logic_vector(to_unsigned(157,8) ,
17385	 => std_logic_vector(to_unsigned(161,8) ,
17386	 => std_logic_vector(to_unsigned(171,8) ,
17387	 => std_logic_vector(to_unsigned(166,8) ,
17388	 => std_logic_vector(to_unsigned(163,8) ,
17389	 => std_logic_vector(to_unsigned(163,8) ,
17390	 => std_logic_vector(to_unsigned(157,8) ,
17391	 => std_logic_vector(to_unsigned(163,8) ,
17392	 => std_logic_vector(to_unsigned(163,8) ,
17393	 => std_logic_vector(to_unsigned(159,8) ,
17394	 => std_logic_vector(to_unsigned(157,8) ,
17395	 => std_logic_vector(to_unsigned(138,8) ,
17396	 => std_logic_vector(to_unsigned(125,8) ,
17397	 => std_logic_vector(to_unsigned(124,8) ,
17398	 => std_logic_vector(to_unsigned(141,8) ,
17399	 => std_logic_vector(to_unsigned(147,8) ,
17400	 => std_logic_vector(to_unsigned(130,8) ,
17401	 => std_logic_vector(to_unsigned(124,8) ,
17402	 => std_logic_vector(to_unsigned(118,8) ,
17403	 => std_logic_vector(to_unsigned(124,8) ,
17404	 => std_logic_vector(to_unsigned(122,8) ,
17405	 => std_logic_vector(to_unsigned(119,8) ,
17406	 => std_logic_vector(to_unsigned(116,8) ,
17407	 => std_logic_vector(to_unsigned(122,8) ,
17408	 => std_logic_vector(to_unsigned(114,8) ,
17409	 => std_logic_vector(to_unsigned(104,8) ,
17410	 => std_logic_vector(to_unsigned(112,8) ,
17411	 => std_logic_vector(to_unsigned(111,8) ,
17412	 => std_logic_vector(to_unsigned(111,8) ,
17413	 => std_logic_vector(to_unsigned(124,8) ,
17414	 => std_logic_vector(to_unsigned(134,8) ,
17415	 => std_logic_vector(to_unsigned(136,8) ,
17416	 => std_logic_vector(to_unsigned(134,8) ,
17417	 => std_logic_vector(to_unsigned(138,8) ,
17418	 => std_logic_vector(to_unsigned(136,8) ,
17419	 => std_logic_vector(to_unsigned(147,8) ,
17420	 => std_logic_vector(to_unsigned(147,8) ,
17421	 => std_logic_vector(to_unsigned(139,8) ,
17422	 => std_logic_vector(to_unsigned(118,8) ,
17423	 => std_logic_vector(to_unsigned(111,8) ,
17424	 => std_logic_vector(to_unsigned(112,8) ,
17425	 => std_logic_vector(to_unsigned(130,8) ,
17426	 => std_logic_vector(to_unsigned(159,8) ,
17427	 => std_logic_vector(to_unsigned(122,8) ,
17428	 => std_logic_vector(to_unsigned(95,8) ,
17429	 => std_logic_vector(to_unsigned(111,8) ,
17430	 => std_logic_vector(to_unsigned(99,8) ,
17431	 => std_logic_vector(to_unsigned(77,8) ,
17432	 => std_logic_vector(to_unsigned(82,8) ,
17433	 => std_logic_vector(to_unsigned(92,8) ,
17434	 => std_logic_vector(to_unsigned(88,8) ,
17435	 => std_logic_vector(to_unsigned(84,8) ,
17436	 => std_logic_vector(to_unsigned(84,8) ,
17437	 => std_logic_vector(to_unsigned(97,8) ,
17438	 => std_logic_vector(to_unsigned(91,8) ,
17439	 => std_logic_vector(to_unsigned(86,8) ,
17440	 => std_logic_vector(to_unsigned(86,8) ,
17441	 => std_logic_vector(to_unsigned(87,8) ,
17442	 => std_logic_vector(to_unsigned(91,8) ,
17443	 => std_logic_vector(to_unsigned(100,8) ,
17444	 => std_logic_vector(to_unsigned(116,8) ,
17445	 => std_logic_vector(to_unsigned(114,8) ,
17446	 => std_logic_vector(to_unsigned(93,8) ,
17447	 => std_logic_vector(to_unsigned(95,8) ,
17448	 => std_logic_vector(to_unsigned(97,8) ,
17449	 => std_logic_vector(to_unsigned(93,8) ,
17450	 => std_logic_vector(to_unsigned(95,8) ,
17451	 => std_logic_vector(to_unsigned(105,8) ,
17452	 => std_logic_vector(to_unsigned(95,8) ,
17453	 => std_logic_vector(to_unsigned(93,8) ,
17454	 => std_logic_vector(to_unsigned(93,8) ,
17455	 => std_logic_vector(to_unsigned(90,8) ,
17456	 => std_logic_vector(to_unsigned(88,8) ,
17457	 => std_logic_vector(to_unsigned(92,8) ,
17458	 => std_logic_vector(to_unsigned(105,8) ,
17459	 => std_logic_vector(to_unsigned(115,8) ,
17460	 => std_logic_vector(to_unsigned(115,8) ,
17461	 => std_logic_vector(to_unsigned(118,8) ,
17462	 => std_logic_vector(to_unsigned(114,8) ,
17463	 => std_logic_vector(to_unsigned(109,8) ,
17464	 => std_logic_vector(to_unsigned(84,8) ,
17465	 => std_logic_vector(to_unsigned(84,8) ,
17466	 => std_logic_vector(to_unsigned(107,8) ,
17467	 => std_logic_vector(to_unsigned(93,8) ,
17468	 => std_logic_vector(to_unsigned(85,8) ,
17469	 => std_logic_vector(to_unsigned(87,8) ,
17470	 => std_logic_vector(to_unsigned(90,8) ,
17471	 => std_logic_vector(to_unsigned(88,8) ,
17472	 => std_logic_vector(to_unsigned(118,8) ,
17473	 => std_logic_vector(to_unsigned(128,8) ,
17474	 => std_logic_vector(to_unsigned(122,8) ,
17475	 => std_logic_vector(to_unsigned(119,8) ,
17476	 => std_logic_vector(to_unsigned(111,8) ,
17477	 => std_logic_vector(to_unsigned(112,8) ,
17478	 => std_logic_vector(to_unsigned(112,8) ,
17479	 => std_logic_vector(to_unsigned(116,8) ,
17480	 => std_logic_vector(to_unsigned(121,8) ,
17481	 => std_logic_vector(to_unsigned(115,8) ,
17482	 => std_logic_vector(to_unsigned(96,8) ,
17483	 => std_logic_vector(to_unsigned(85,8) ,
17484	 => std_logic_vector(to_unsigned(84,8) ,
17485	 => std_logic_vector(to_unsigned(68,8) ,
17486	 => std_logic_vector(to_unsigned(60,8) ,
17487	 => std_logic_vector(to_unsigned(54,8) ,
17488	 => std_logic_vector(to_unsigned(66,8) ,
17489	 => std_logic_vector(to_unsigned(78,8) ,
17490	 => std_logic_vector(to_unsigned(68,8) ,
17491	 => std_logic_vector(to_unsigned(61,8) ,
17492	 => std_logic_vector(to_unsigned(51,8) ,
17493	 => std_logic_vector(to_unsigned(45,8) ,
17494	 => std_logic_vector(to_unsigned(47,8) ,
17495	 => std_logic_vector(to_unsigned(55,8) ,
17496	 => std_logic_vector(to_unsigned(68,8) ,
17497	 => std_logic_vector(to_unsigned(65,8) ,
17498	 => std_logic_vector(to_unsigned(65,8) ,
17499	 => std_logic_vector(to_unsigned(68,8) ,
17500	 => std_logic_vector(to_unsigned(66,8) ,
17501	 => std_logic_vector(to_unsigned(61,8) ,
17502	 => std_logic_vector(to_unsigned(59,8) ,
17503	 => std_logic_vector(to_unsigned(72,8) ,
17504	 => std_logic_vector(to_unsigned(66,8) ,
17505	 => std_logic_vector(to_unsigned(58,8) ,
17506	 => std_logic_vector(to_unsigned(69,8) ,
17507	 => std_logic_vector(to_unsigned(85,8) ,
17508	 => std_logic_vector(to_unsigned(80,8) ,
17509	 => std_logic_vector(to_unsigned(73,8) ,
17510	 => std_logic_vector(to_unsigned(74,8) ,
17511	 => std_logic_vector(to_unsigned(70,8) ,
17512	 => std_logic_vector(to_unsigned(69,8) ,
17513	 => std_logic_vector(to_unsigned(72,8) ,
17514	 => std_logic_vector(to_unsigned(66,8) ,
17515	 => std_logic_vector(to_unsigned(71,8) ,
17516	 => std_logic_vector(to_unsigned(74,8) ,
17517	 => std_logic_vector(to_unsigned(73,8) ,
17518	 => std_logic_vector(to_unsigned(76,8) ,
17519	 => std_logic_vector(to_unsigned(72,8) ,
17520	 => std_logic_vector(to_unsigned(65,8) ,
17521	 => std_logic_vector(to_unsigned(72,8) ,
17522	 => std_logic_vector(to_unsigned(74,8) ,
17523	 => std_logic_vector(to_unsigned(90,8) ,
17524	 => std_logic_vector(to_unsigned(81,8) ,
17525	 => std_logic_vector(to_unsigned(79,8) ,
17526	 => std_logic_vector(to_unsigned(78,8) ,
17527	 => std_logic_vector(to_unsigned(81,8) ,
17528	 => std_logic_vector(to_unsigned(82,8) ,
17529	 => std_logic_vector(to_unsigned(8,8) ,
17530	 => std_logic_vector(to_unsigned(0,8) ,
17531	 => std_logic_vector(to_unsigned(1,8) ,
17532	 => std_logic_vector(to_unsigned(41,8) ,
17533	 => std_logic_vector(to_unsigned(111,8) ,
17534	 => std_logic_vector(to_unsigned(76,8) ,
17535	 => std_logic_vector(to_unsigned(71,8) ,
17536	 => std_logic_vector(to_unsigned(72,8) ,
17537	 => std_logic_vector(to_unsigned(79,8) ,
17538	 => std_logic_vector(to_unsigned(87,8) ,
17539	 => std_logic_vector(to_unsigned(88,8) ,
17540	 => std_logic_vector(to_unsigned(87,8) ,
17541	 => std_logic_vector(to_unsigned(90,8) ,
17542	 => std_logic_vector(to_unsigned(80,8) ,
17543	 => std_logic_vector(to_unsigned(82,8) ,
17544	 => std_logic_vector(to_unsigned(97,8) ,
17545	 => std_logic_vector(to_unsigned(92,8) ,
17546	 => std_logic_vector(to_unsigned(81,8) ,
17547	 => std_logic_vector(to_unsigned(73,8) ,
17548	 => std_logic_vector(to_unsigned(74,8) ,
17549	 => std_logic_vector(to_unsigned(81,8) ,
17550	 => std_logic_vector(to_unsigned(85,8) ,
17551	 => std_logic_vector(to_unsigned(74,8) ,
17552	 => std_logic_vector(to_unsigned(72,8) ,
17553	 => std_logic_vector(to_unsigned(76,8) ,
17554	 => std_logic_vector(to_unsigned(74,8) ,
17555	 => std_logic_vector(to_unsigned(80,8) ,
17556	 => std_logic_vector(to_unsigned(78,8) ,
17557	 => std_logic_vector(to_unsigned(77,8) ,
17558	 => std_logic_vector(to_unsigned(71,8) ,
17559	 => std_logic_vector(to_unsigned(69,8) ,
17560	 => std_logic_vector(to_unsigned(69,8) ,
17561	 => std_logic_vector(to_unsigned(67,8) ,
17562	 => std_logic_vector(to_unsigned(71,8) ,
17563	 => std_logic_vector(to_unsigned(70,8) ,
17564	 => std_logic_vector(to_unsigned(71,8) ,
17565	 => std_logic_vector(to_unsigned(85,8) ,
17566	 => std_logic_vector(to_unsigned(82,8) ,
17567	 => std_logic_vector(to_unsigned(77,8) ,
17568	 => std_logic_vector(to_unsigned(77,8) ,
17569	 => std_logic_vector(to_unsigned(84,8) ,
17570	 => std_logic_vector(to_unsigned(82,8) ,
17571	 => std_logic_vector(to_unsigned(73,8) ,
17572	 => std_logic_vector(to_unsigned(81,8) ,
17573	 => std_logic_vector(to_unsigned(80,8) ,
17574	 => std_logic_vector(to_unsigned(78,8) ,
17575	 => std_logic_vector(to_unsigned(84,8) ,
17576	 => std_logic_vector(to_unsigned(77,8) ,
17577	 => std_logic_vector(to_unsigned(84,8) ,
17578	 => std_logic_vector(to_unsigned(88,8) ,
17579	 => std_logic_vector(to_unsigned(79,8) ,
17580	 => std_logic_vector(to_unsigned(79,8) ,
17581	 => std_logic_vector(to_unsigned(85,8) ,
17582	 => std_logic_vector(to_unsigned(86,8) ,
17583	 => std_logic_vector(to_unsigned(87,8) ,
17584	 => std_logic_vector(to_unsigned(91,8) ,
17585	 => std_logic_vector(to_unsigned(86,8) ,
17586	 => std_logic_vector(to_unsigned(79,8) ,
17587	 => std_logic_vector(to_unsigned(87,8) ,
17588	 => std_logic_vector(to_unsigned(90,8) ,
17589	 => std_logic_vector(to_unsigned(85,8) ,
17590	 => std_logic_vector(to_unsigned(87,8) ,
17591	 => std_logic_vector(to_unsigned(87,8) ,
17592	 => std_logic_vector(to_unsigned(81,8) ,
17593	 => std_logic_vector(to_unsigned(80,8) ,
17594	 => std_logic_vector(to_unsigned(82,8) ,
17595	 => std_logic_vector(to_unsigned(88,8) ,
17596	 => std_logic_vector(to_unsigned(95,8) ,
17597	 => std_logic_vector(to_unsigned(87,8) ,
17598	 => std_logic_vector(to_unsigned(86,8) ,
17599	 => std_logic_vector(to_unsigned(90,8) ,
17600	 => std_logic_vector(to_unsigned(90,8) ,
17601	 => std_logic_vector(to_unsigned(144,8) ,
17602	 => std_logic_vector(to_unsigned(142,8) ,
17603	 => std_logic_vector(to_unsigned(142,8) ,
17604	 => std_logic_vector(to_unsigned(144,8) ,
17605	 => std_logic_vector(to_unsigned(147,8) ,
17606	 => std_logic_vector(to_unsigned(152,8) ,
17607	 => std_logic_vector(to_unsigned(154,8) ,
17608	 => std_logic_vector(to_unsigned(154,8) ,
17609	 => std_logic_vector(to_unsigned(156,8) ,
17610	 => std_logic_vector(to_unsigned(154,8) ,
17611	 => std_logic_vector(to_unsigned(146,8) ,
17612	 => std_logic_vector(to_unsigned(149,8) ,
17613	 => std_logic_vector(to_unsigned(154,8) ,
17614	 => std_logic_vector(to_unsigned(157,8) ,
17615	 => std_logic_vector(to_unsigned(152,8) ,
17616	 => std_logic_vector(to_unsigned(156,8) ,
17617	 => std_logic_vector(to_unsigned(159,8) ,
17618	 => std_logic_vector(to_unsigned(152,8) ,
17619	 => std_logic_vector(to_unsigned(149,8) ,
17620	 => std_logic_vector(to_unsigned(151,8) ,
17621	 => std_logic_vector(to_unsigned(144,8) ,
17622	 => std_logic_vector(to_unsigned(147,8) ,
17623	 => std_logic_vector(to_unsigned(156,8) ,
17624	 => std_logic_vector(to_unsigned(154,8) ,
17625	 => std_logic_vector(to_unsigned(156,8) ,
17626	 => std_logic_vector(to_unsigned(151,8) ,
17627	 => std_logic_vector(to_unsigned(151,8) ,
17628	 => std_logic_vector(to_unsigned(164,8) ,
17629	 => std_logic_vector(to_unsigned(79,8) ,
17630	 => std_logic_vector(to_unsigned(45,8) ,
17631	 => std_logic_vector(to_unsigned(46,8) ,
17632	 => std_logic_vector(to_unsigned(18,8) ,
17633	 => std_logic_vector(to_unsigned(12,8) ,
17634	 => std_logic_vector(to_unsigned(7,8) ,
17635	 => std_logic_vector(to_unsigned(79,8) ,
17636	 => std_logic_vector(to_unsigned(173,8) ,
17637	 => std_logic_vector(to_unsigned(147,8) ,
17638	 => std_logic_vector(to_unsigned(151,8) ,
17639	 => std_logic_vector(to_unsigned(152,8) ,
17640	 => std_logic_vector(to_unsigned(141,8) ,
17641	 => std_logic_vector(to_unsigned(144,8) ,
17642	 => std_logic_vector(to_unsigned(151,8) ,
17643	 => std_logic_vector(to_unsigned(152,8) ,
17644	 => std_logic_vector(to_unsigned(149,8) ,
17645	 => std_logic_vector(to_unsigned(152,8) ,
17646	 => std_logic_vector(to_unsigned(154,8) ,
17647	 => std_logic_vector(to_unsigned(146,8) ,
17648	 => std_logic_vector(to_unsigned(154,8) ,
17649	 => std_logic_vector(to_unsigned(157,8) ,
17650	 => std_logic_vector(to_unsigned(156,8) ,
17651	 => std_logic_vector(to_unsigned(154,8) ,
17652	 => std_logic_vector(to_unsigned(152,8) ,
17653	 => std_logic_vector(to_unsigned(147,8) ,
17654	 => std_logic_vector(to_unsigned(146,8) ,
17655	 => std_logic_vector(to_unsigned(146,8) ,
17656	 => std_logic_vector(to_unsigned(100,8) ,
17657	 => std_logic_vector(to_unsigned(63,8) ,
17658	 => std_logic_vector(to_unsigned(72,8) ,
17659	 => std_logic_vector(to_unsigned(77,8) ,
17660	 => std_logic_vector(to_unsigned(72,8) ,
17661	 => std_logic_vector(to_unsigned(74,8) ,
17662	 => std_logic_vector(to_unsigned(71,8) ,
17663	 => std_logic_vector(to_unsigned(56,8) ,
17664	 => std_logic_vector(to_unsigned(51,8) ,
17665	 => std_logic_vector(to_unsigned(52,8) ,
17666	 => std_logic_vector(to_unsigned(45,8) ,
17667	 => std_logic_vector(to_unsigned(76,8) ,
17668	 => std_logic_vector(to_unsigned(139,8) ,
17669	 => std_logic_vector(to_unsigned(156,8) ,
17670	 => std_logic_vector(to_unsigned(154,8) ,
17671	 => std_logic_vector(to_unsigned(159,8) ,
17672	 => std_logic_vector(to_unsigned(159,8) ,
17673	 => std_logic_vector(to_unsigned(166,8) ,
17674	 => std_logic_vector(to_unsigned(163,8) ,
17675	 => std_logic_vector(to_unsigned(147,8) ,
17676	 => std_logic_vector(to_unsigned(149,8) ,
17677	 => std_logic_vector(to_unsigned(151,8) ,
17678	 => std_logic_vector(to_unsigned(142,8) ,
17679	 => std_logic_vector(to_unsigned(134,8) ,
17680	 => std_logic_vector(to_unsigned(139,8) ,
17681	 => std_logic_vector(to_unsigned(128,8) ,
17682	 => std_logic_vector(to_unsigned(133,8) ,
17683	 => std_logic_vector(to_unsigned(149,8) ,
17684	 => std_logic_vector(to_unsigned(142,8) ,
17685	 => std_logic_vector(to_unsigned(154,8) ,
17686	 => std_logic_vector(to_unsigned(166,8) ,
17687	 => std_logic_vector(to_unsigned(146,8) ,
17688	 => std_logic_vector(to_unsigned(20,8) ,
17689	 => std_logic_vector(to_unsigned(0,8) ,
17690	 => std_logic_vector(to_unsigned(1,8) ,
17691	 => std_logic_vector(to_unsigned(2,8) ,
17692	 => std_logic_vector(to_unsigned(2,8) ,
17693	 => std_logic_vector(to_unsigned(1,8) ,
17694	 => std_logic_vector(to_unsigned(1,8) ,
17695	 => std_logic_vector(to_unsigned(2,8) ,
17696	 => std_logic_vector(to_unsigned(3,8) ,
17697	 => std_logic_vector(to_unsigned(2,8) ,
17698	 => std_logic_vector(to_unsigned(2,8) ,
17699	 => std_logic_vector(to_unsigned(2,8) ,
17700	 => std_logic_vector(to_unsigned(4,8) ,
17701	 => std_logic_vector(to_unsigned(1,8) ,
17702	 => std_logic_vector(to_unsigned(43,8) ,
17703	 => std_logic_vector(to_unsigned(181,8) ,
17704	 => std_logic_vector(to_unsigned(163,8) ,
17705	 => std_logic_vector(to_unsigned(170,8) ,
17706	 => std_logic_vector(to_unsigned(170,8) ,
17707	 => std_logic_vector(to_unsigned(168,8) ,
17708	 => std_logic_vector(to_unsigned(163,8) ,
17709	 => std_logic_vector(to_unsigned(161,8) ,
17710	 => std_logic_vector(to_unsigned(159,8) ,
17711	 => std_logic_vector(to_unsigned(159,8) ,
17712	 => std_logic_vector(to_unsigned(163,8) ,
17713	 => std_logic_vector(to_unsigned(156,8) ,
17714	 => std_logic_vector(to_unsigned(154,8) ,
17715	 => std_logic_vector(to_unsigned(154,8) ,
17716	 => std_logic_vector(to_unsigned(130,8) ,
17717	 => std_logic_vector(to_unsigned(122,8) ,
17718	 => std_logic_vector(to_unsigned(134,8) ,
17719	 => std_logic_vector(to_unsigned(146,8) ,
17720	 => std_logic_vector(to_unsigned(131,8) ,
17721	 => std_logic_vector(to_unsigned(131,8) ,
17722	 => std_logic_vector(to_unsigned(133,8) ,
17723	 => std_logic_vector(to_unsigned(128,8) ,
17724	 => std_logic_vector(to_unsigned(147,8) ,
17725	 => std_logic_vector(to_unsigned(151,8) ,
17726	 => std_logic_vector(to_unsigned(142,8) ,
17727	 => std_logic_vector(to_unsigned(133,8) ,
17728	 => std_logic_vector(to_unsigned(139,8) ,
17729	 => std_logic_vector(to_unsigned(131,8) ,
17730	 => std_logic_vector(to_unsigned(119,8) ,
17731	 => std_logic_vector(to_unsigned(116,8) ,
17732	 => std_logic_vector(to_unsigned(112,8) ,
17733	 => std_logic_vector(to_unsigned(124,8) ,
17734	 => std_logic_vector(to_unsigned(146,8) ,
17735	 => std_logic_vector(to_unsigned(142,8) ,
17736	 => std_logic_vector(to_unsigned(133,8) ,
17737	 => std_logic_vector(to_unsigned(141,8) ,
17738	 => std_logic_vector(to_unsigned(133,8) ,
17739	 => std_logic_vector(to_unsigned(138,8) ,
17740	 => std_logic_vector(to_unsigned(136,8) ,
17741	 => std_logic_vector(to_unsigned(128,8) ,
17742	 => std_logic_vector(to_unsigned(128,8) ,
17743	 => std_logic_vector(to_unsigned(118,8) ,
17744	 => std_logic_vector(to_unsigned(119,8) ,
17745	 => std_logic_vector(to_unsigned(142,8) ,
17746	 => std_logic_vector(to_unsigned(161,8) ,
17747	 => std_logic_vector(to_unsigned(119,8) ,
17748	 => std_logic_vector(to_unsigned(100,8) ,
17749	 => std_logic_vector(to_unsigned(141,8) ,
17750	 => std_logic_vector(to_unsigned(115,8) ,
17751	 => std_logic_vector(to_unsigned(84,8) ,
17752	 => std_logic_vector(to_unsigned(111,8) ,
17753	 => std_logic_vector(to_unsigned(131,8) ,
17754	 => std_logic_vector(to_unsigned(112,8) ,
17755	 => std_logic_vector(to_unsigned(95,8) ,
17756	 => std_logic_vector(to_unsigned(86,8) ,
17757	 => std_logic_vector(to_unsigned(86,8) ,
17758	 => std_logic_vector(to_unsigned(85,8) ,
17759	 => std_logic_vector(to_unsigned(70,8) ,
17760	 => std_logic_vector(to_unsigned(77,8) ,
17761	 => std_logic_vector(to_unsigned(81,8) ,
17762	 => std_logic_vector(to_unsigned(84,8) ,
17763	 => std_logic_vector(to_unsigned(95,8) ,
17764	 => std_logic_vector(to_unsigned(107,8) ,
17765	 => std_logic_vector(to_unsigned(116,8) ,
17766	 => std_logic_vector(to_unsigned(100,8) ,
17767	 => std_logic_vector(to_unsigned(93,8) ,
17768	 => std_logic_vector(to_unsigned(100,8) ,
17769	 => std_logic_vector(to_unsigned(96,8) ,
17770	 => std_logic_vector(to_unsigned(86,8) ,
17771	 => std_logic_vector(to_unsigned(97,8) ,
17772	 => std_logic_vector(to_unsigned(131,8) ,
17773	 => std_logic_vector(to_unsigned(130,8) ,
17774	 => std_logic_vector(to_unsigned(104,8) ,
17775	 => std_logic_vector(to_unsigned(93,8) ,
17776	 => std_logic_vector(to_unsigned(95,8) ,
17777	 => std_logic_vector(to_unsigned(96,8) ,
17778	 => std_logic_vector(to_unsigned(105,8) ,
17779	 => std_logic_vector(to_unsigned(119,8) ,
17780	 => std_logic_vector(to_unsigned(125,8) ,
17781	 => std_logic_vector(to_unsigned(131,8) ,
17782	 => std_logic_vector(to_unsigned(124,8) ,
17783	 => std_logic_vector(to_unsigned(118,8) ,
17784	 => std_logic_vector(to_unsigned(86,8) ,
17785	 => std_logic_vector(to_unsigned(72,8) ,
17786	 => std_logic_vector(to_unsigned(90,8) ,
17787	 => std_logic_vector(to_unsigned(90,8) ,
17788	 => std_logic_vector(to_unsigned(92,8) ,
17789	 => std_logic_vector(to_unsigned(92,8) ,
17790	 => std_logic_vector(to_unsigned(86,8) ,
17791	 => std_logic_vector(to_unsigned(88,8) ,
17792	 => std_logic_vector(to_unsigned(104,8) ,
17793	 => std_logic_vector(to_unsigned(133,8) ,
17794	 => std_logic_vector(to_unsigned(138,8) ,
17795	 => std_logic_vector(to_unsigned(118,8) ,
17796	 => std_logic_vector(to_unsigned(96,8) ,
17797	 => std_logic_vector(to_unsigned(92,8) ,
17798	 => std_logic_vector(to_unsigned(99,8) ,
17799	 => std_logic_vector(to_unsigned(92,8) ,
17800	 => std_logic_vector(to_unsigned(74,8) ,
17801	 => std_logic_vector(to_unsigned(70,8) ,
17802	 => std_logic_vector(to_unsigned(77,8) ,
17803	 => std_logic_vector(to_unsigned(72,8) ,
17804	 => std_logic_vector(to_unsigned(71,8) ,
17805	 => std_logic_vector(to_unsigned(64,8) ,
17806	 => std_logic_vector(to_unsigned(56,8) ,
17807	 => std_logic_vector(to_unsigned(56,8) ,
17808	 => std_logic_vector(to_unsigned(61,8) ,
17809	 => std_logic_vector(to_unsigned(69,8) ,
17810	 => std_logic_vector(to_unsigned(67,8) ,
17811	 => std_logic_vector(to_unsigned(72,8) ,
17812	 => std_logic_vector(to_unsigned(67,8) ,
17813	 => std_logic_vector(to_unsigned(56,8) ,
17814	 => std_logic_vector(to_unsigned(58,8) ,
17815	 => std_logic_vector(to_unsigned(70,8) ,
17816	 => std_logic_vector(to_unsigned(79,8) ,
17817	 => std_logic_vector(to_unsigned(72,8) ,
17818	 => std_logic_vector(to_unsigned(77,8) ,
17819	 => std_logic_vector(to_unsigned(72,8) ,
17820	 => std_logic_vector(to_unsigned(70,8) ,
17821	 => std_logic_vector(to_unsigned(62,8) ,
17822	 => std_logic_vector(to_unsigned(55,8) ,
17823	 => std_logic_vector(to_unsigned(66,8) ,
17824	 => std_logic_vector(to_unsigned(66,8) ,
17825	 => std_logic_vector(to_unsigned(67,8) ,
17826	 => std_logic_vector(to_unsigned(74,8) ,
17827	 => std_logic_vector(to_unsigned(77,8) ,
17828	 => std_logic_vector(to_unsigned(66,8) ,
17829	 => std_logic_vector(to_unsigned(72,8) ,
17830	 => std_logic_vector(to_unsigned(71,8) ,
17831	 => std_logic_vector(to_unsigned(61,8) ,
17832	 => std_logic_vector(to_unsigned(63,8) ,
17833	 => std_logic_vector(to_unsigned(62,8) ,
17834	 => std_logic_vector(to_unsigned(67,8) ,
17835	 => std_logic_vector(to_unsigned(71,8) ,
17836	 => std_logic_vector(to_unsigned(71,8) ,
17837	 => std_logic_vector(to_unsigned(64,8) ,
17838	 => std_logic_vector(to_unsigned(69,8) ,
17839	 => std_logic_vector(to_unsigned(79,8) ,
17840	 => std_logic_vector(to_unsigned(76,8) ,
17841	 => std_logic_vector(to_unsigned(76,8) ,
17842	 => std_logic_vector(to_unsigned(78,8) ,
17843	 => std_logic_vector(to_unsigned(96,8) ,
17844	 => std_logic_vector(to_unsigned(112,8) ,
17845	 => std_logic_vector(to_unsigned(108,8) ,
17846	 => std_logic_vector(to_unsigned(105,8) ,
17847	 => std_logic_vector(to_unsigned(97,8) ,
17848	 => std_logic_vector(to_unsigned(115,8) ,
17849	 => std_logic_vector(to_unsigned(33,8) ,
17850	 => std_logic_vector(to_unsigned(0,8) ,
17851	 => std_logic_vector(to_unsigned(0,8) ,
17852	 => std_logic_vector(to_unsigned(22,8) ,
17853	 => std_logic_vector(to_unsigned(138,8) ,
17854	 => std_logic_vector(to_unsigned(101,8) ,
17855	 => std_logic_vector(to_unsigned(84,8) ,
17856	 => std_logic_vector(to_unsigned(88,8) ,
17857	 => std_logic_vector(to_unsigned(91,8) ,
17858	 => std_logic_vector(to_unsigned(96,8) ,
17859	 => std_logic_vector(to_unsigned(112,8) ,
17860	 => std_logic_vector(to_unsigned(97,8) ,
17861	 => std_logic_vector(to_unsigned(81,8) ,
17862	 => std_logic_vector(to_unsigned(87,8) ,
17863	 => std_logic_vector(to_unsigned(90,8) ,
17864	 => std_logic_vector(to_unsigned(100,8) ,
17865	 => std_logic_vector(to_unsigned(104,8) ,
17866	 => std_logic_vector(to_unsigned(91,8) ,
17867	 => std_logic_vector(to_unsigned(79,8) ,
17868	 => std_logic_vector(to_unsigned(79,8) ,
17869	 => std_logic_vector(to_unsigned(82,8) ,
17870	 => std_logic_vector(to_unsigned(78,8) ,
17871	 => std_logic_vector(to_unsigned(71,8) ,
17872	 => std_logic_vector(to_unsigned(74,8) ,
17873	 => std_logic_vector(to_unsigned(77,8) ,
17874	 => std_logic_vector(to_unsigned(81,8) ,
17875	 => std_logic_vector(to_unsigned(84,8) ,
17876	 => std_logic_vector(to_unsigned(78,8) ,
17877	 => std_logic_vector(to_unsigned(76,8) ,
17878	 => std_logic_vector(to_unsigned(73,8) ,
17879	 => std_logic_vector(to_unsigned(77,8) ,
17880	 => std_logic_vector(to_unsigned(76,8) ,
17881	 => std_logic_vector(to_unsigned(74,8) ,
17882	 => std_logic_vector(to_unsigned(74,8) ,
17883	 => std_logic_vector(to_unsigned(67,8) ,
17884	 => std_logic_vector(to_unsigned(72,8) ,
17885	 => std_logic_vector(to_unsigned(84,8) ,
17886	 => std_logic_vector(to_unsigned(87,8) ,
17887	 => std_logic_vector(to_unsigned(82,8) ,
17888	 => std_logic_vector(to_unsigned(78,8) ,
17889	 => std_logic_vector(to_unsigned(84,8) ,
17890	 => std_logic_vector(to_unsigned(88,8) ,
17891	 => std_logic_vector(to_unsigned(87,8) ,
17892	 => std_logic_vector(to_unsigned(82,8) ,
17893	 => std_logic_vector(to_unsigned(78,8) ,
17894	 => std_logic_vector(to_unsigned(81,8) ,
17895	 => std_logic_vector(to_unsigned(81,8) ,
17896	 => std_logic_vector(to_unsigned(79,8) ,
17897	 => std_logic_vector(to_unsigned(82,8) ,
17898	 => std_logic_vector(to_unsigned(88,8) ,
17899	 => std_logic_vector(to_unsigned(84,8) ,
17900	 => std_logic_vector(to_unsigned(74,8) ,
17901	 => std_logic_vector(to_unsigned(73,8) ,
17902	 => std_logic_vector(to_unsigned(85,8) ,
17903	 => std_logic_vector(to_unsigned(88,8) ,
17904	 => std_logic_vector(to_unsigned(84,8) ,
17905	 => std_logic_vector(to_unsigned(87,8) ,
17906	 => std_logic_vector(to_unsigned(86,8) ,
17907	 => std_logic_vector(to_unsigned(87,8) ,
17908	 => std_logic_vector(to_unsigned(88,8) ,
17909	 => std_logic_vector(to_unsigned(84,8) ,
17910	 => std_logic_vector(to_unsigned(86,8) ,
17911	 => std_logic_vector(to_unsigned(86,8) ,
17912	 => std_logic_vector(to_unsigned(84,8) ,
17913	 => std_logic_vector(to_unsigned(85,8) ,
17914	 => std_logic_vector(to_unsigned(80,8) ,
17915	 => std_logic_vector(to_unsigned(84,8) ,
17916	 => std_logic_vector(to_unsigned(91,8) ,
17917	 => std_logic_vector(to_unsigned(84,8) ,
17918	 => std_logic_vector(to_unsigned(84,8) ,
17919	 => std_logic_vector(to_unsigned(90,8) ,
17920	 => std_logic_vector(to_unsigned(87,8) ,
17921	 => std_logic_vector(to_unsigned(144,8) ,
17922	 => std_logic_vector(to_unsigned(149,8) ,
17923	 => std_logic_vector(to_unsigned(152,8) ,
17924	 => std_logic_vector(to_unsigned(151,8) ,
17925	 => std_logic_vector(to_unsigned(152,8) ,
17926	 => std_logic_vector(to_unsigned(151,8) ,
17927	 => std_logic_vector(to_unsigned(151,8) ,
17928	 => std_logic_vector(to_unsigned(154,8) ,
17929	 => std_logic_vector(to_unsigned(157,8) ,
17930	 => std_logic_vector(to_unsigned(159,8) ,
17931	 => std_logic_vector(to_unsigned(154,8) ,
17932	 => std_logic_vector(to_unsigned(152,8) ,
17933	 => std_logic_vector(to_unsigned(152,8) ,
17934	 => std_logic_vector(to_unsigned(157,8) ,
17935	 => std_logic_vector(to_unsigned(156,8) ,
17936	 => std_logic_vector(to_unsigned(154,8) ,
17937	 => std_logic_vector(to_unsigned(154,8) ,
17938	 => std_logic_vector(to_unsigned(146,8) ,
17939	 => std_logic_vector(to_unsigned(147,8) ,
17940	 => std_logic_vector(to_unsigned(147,8) ,
17941	 => std_logic_vector(to_unsigned(147,8) ,
17942	 => std_logic_vector(to_unsigned(151,8) ,
17943	 => std_logic_vector(to_unsigned(154,8) ,
17944	 => std_logic_vector(to_unsigned(161,8) ,
17945	 => std_logic_vector(to_unsigned(152,8) ,
17946	 => std_logic_vector(to_unsigned(151,8) ,
17947	 => std_logic_vector(to_unsigned(170,8) ,
17948	 => std_logic_vector(to_unsigned(76,8) ,
17949	 => std_logic_vector(to_unsigned(9,8) ,
17950	 => std_logic_vector(to_unsigned(7,8) ,
17951	 => std_logic_vector(to_unsigned(8,8) ,
17952	 => std_logic_vector(to_unsigned(2,8) ,
17953	 => std_logic_vector(to_unsigned(2,8) ,
17954	 => std_logic_vector(to_unsigned(6,8) ,
17955	 => std_logic_vector(to_unsigned(54,8) ,
17956	 => std_logic_vector(to_unsigned(139,8) ,
17957	 => std_logic_vector(to_unsigned(163,8) ,
17958	 => std_logic_vector(to_unsigned(157,8) ,
17959	 => std_logic_vector(to_unsigned(159,8) ,
17960	 => std_logic_vector(to_unsigned(156,8) ,
17961	 => std_logic_vector(to_unsigned(156,8) ,
17962	 => std_logic_vector(to_unsigned(157,8) ,
17963	 => std_logic_vector(to_unsigned(159,8) ,
17964	 => std_logic_vector(to_unsigned(154,8) ,
17965	 => std_logic_vector(to_unsigned(156,8) ,
17966	 => std_logic_vector(to_unsigned(163,8) ,
17967	 => std_logic_vector(to_unsigned(164,8) ,
17968	 => std_logic_vector(to_unsigned(161,8) ,
17969	 => std_logic_vector(to_unsigned(152,8) ,
17970	 => std_logic_vector(to_unsigned(152,8) ,
17971	 => std_logic_vector(to_unsigned(157,8) ,
17972	 => std_logic_vector(to_unsigned(144,8) ,
17973	 => std_logic_vector(to_unsigned(139,8) ,
17974	 => std_logic_vector(to_unsigned(149,8) ,
17975	 => std_logic_vector(to_unsigned(91,8) ,
17976	 => std_logic_vector(to_unsigned(35,8) ,
17977	 => std_logic_vector(to_unsigned(51,8) ,
17978	 => std_logic_vector(to_unsigned(87,8) ,
17979	 => std_logic_vector(to_unsigned(70,8) ,
17980	 => std_logic_vector(to_unsigned(72,8) ,
17981	 => std_logic_vector(to_unsigned(77,8) ,
17982	 => std_logic_vector(to_unsigned(65,8) ,
17983	 => std_logic_vector(to_unsigned(62,8) ,
17984	 => std_logic_vector(to_unsigned(40,8) ,
17985	 => std_logic_vector(to_unsigned(60,8) ,
17986	 => std_logic_vector(to_unsigned(49,8) ,
17987	 => std_logic_vector(to_unsigned(30,8) ,
17988	 => std_logic_vector(to_unsigned(71,8) ,
17989	 => std_logic_vector(to_unsigned(157,8) ,
17990	 => std_logic_vector(to_unsigned(163,8) ,
17991	 => std_logic_vector(to_unsigned(163,8) ,
17992	 => std_logic_vector(to_unsigned(163,8) ,
17993	 => std_logic_vector(to_unsigned(164,8) ,
17994	 => std_logic_vector(to_unsigned(159,8) ,
17995	 => std_logic_vector(to_unsigned(144,8) ,
17996	 => std_logic_vector(to_unsigned(139,8) ,
17997	 => std_logic_vector(to_unsigned(147,8) ,
17998	 => std_logic_vector(to_unsigned(146,8) ,
17999	 => std_logic_vector(to_unsigned(147,8) ,
18000	 => std_logic_vector(to_unsigned(149,8) ,
18001	 => std_logic_vector(to_unsigned(156,8) ,
18002	 => std_logic_vector(to_unsigned(159,8) ,
18003	 => std_logic_vector(to_unsigned(164,8) ,
18004	 => std_logic_vector(to_unsigned(159,8) ,
18005	 => std_logic_vector(to_unsigned(156,8) ,
18006	 => std_logic_vector(to_unsigned(186,8) ,
18007	 => std_logic_vector(to_unsigned(68,8) ,
18008	 => std_logic_vector(to_unsigned(1,8) ,
18009	 => std_logic_vector(to_unsigned(1,8) ,
18010	 => std_logic_vector(to_unsigned(1,8) ,
18011	 => std_logic_vector(to_unsigned(1,8) ,
18012	 => std_logic_vector(to_unsigned(1,8) ,
18013	 => std_logic_vector(to_unsigned(1,8) ,
18014	 => std_logic_vector(to_unsigned(1,8) ,
18015	 => std_logic_vector(to_unsigned(1,8) ,
18016	 => std_logic_vector(to_unsigned(2,8) ,
18017	 => std_logic_vector(to_unsigned(3,8) ,
18018	 => std_logic_vector(to_unsigned(2,8) ,
18019	 => std_logic_vector(to_unsigned(2,8) ,
18020	 => std_logic_vector(to_unsigned(3,8) ,
18021	 => std_logic_vector(to_unsigned(1,8) ,
18022	 => std_logic_vector(to_unsigned(44,8) ,
18023	 => std_logic_vector(to_unsigned(186,8) ,
18024	 => std_logic_vector(to_unsigned(170,8) ,
18025	 => std_logic_vector(to_unsigned(166,8) ,
18026	 => std_logic_vector(to_unsigned(168,8) ,
18027	 => std_logic_vector(to_unsigned(170,8) ,
18028	 => std_logic_vector(to_unsigned(166,8) ,
18029	 => std_logic_vector(to_unsigned(163,8) ,
18030	 => std_logic_vector(to_unsigned(163,8) ,
18031	 => std_logic_vector(to_unsigned(163,8) ,
18032	 => std_logic_vector(to_unsigned(159,8) ,
18033	 => std_logic_vector(to_unsigned(152,8) ,
18034	 => std_logic_vector(to_unsigned(146,8) ,
18035	 => std_logic_vector(to_unsigned(154,8) ,
18036	 => std_logic_vector(to_unsigned(142,8) ,
18037	 => std_logic_vector(to_unsigned(134,8) ,
18038	 => std_logic_vector(to_unsigned(133,8) ,
18039	 => std_logic_vector(to_unsigned(133,8) ,
18040	 => std_logic_vector(to_unsigned(133,8) ,
18041	 => std_logic_vector(to_unsigned(136,8) ,
18042	 => std_logic_vector(to_unsigned(142,8) ,
18043	 => std_logic_vector(to_unsigned(139,8) ,
18044	 => std_logic_vector(to_unsigned(163,8) ,
18045	 => std_logic_vector(to_unsigned(166,8) ,
18046	 => std_logic_vector(to_unsigned(159,8) ,
18047	 => std_logic_vector(to_unsigned(144,8) ,
18048	 => std_logic_vector(to_unsigned(156,8) ,
18049	 => std_logic_vector(to_unsigned(152,8) ,
18050	 => std_logic_vector(to_unsigned(127,8) ,
18051	 => std_logic_vector(to_unsigned(127,8) ,
18052	 => std_logic_vector(to_unsigned(146,8) ,
18053	 => std_logic_vector(to_unsigned(136,8) ,
18054	 => std_logic_vector(to_unsigned(133,8) ,
18055	 => std_logic_vector(to_unsigned(139,8) ,
18056	 => std_logic_vector(to_unsigned(146,8) ,
18057	 => std_logic_vector(to_unsigned(151,8) ,
18058	 => std_logic_vector(to_unsigned(136,8) ,
18059	 => std_logic_vector(to_unsigned(139,8) ,
18060	 => std_logic_vector(to_unsigned(139,8) ,
18061	 => std_logic_vector(to_unsigned(118,8) ,
18062	 => std_logic_vector(to_unsigned(121,8) ,
18063	 => std_logic_vector(to_unsigned(121,8) ,
18064	 => std_logic_vector(to_unsigned(119,8) ,
18065	 => std_logic_vector(to_unsigned(124,8) ,
18066	 => std_logic_vector(to_unsigned(144,8) ,
18067	 => std_logic_vector(to_unsigned(124,8) ,
18068	 => std_logic_vector(to_unsigned(109,8) ,
18069	 => std_logic_vector(to_unsigned(141,8) ,
18070	 => std_logic_vector(to_unsigned(112,8) ,
18071	 => std_logic_vector(to_unsigned(96,8) ,
18072	 => std_logic_vector(to_unsigned(131,8) ,
18073	 => std_logic_vector(to_unsigned(146,8) ,
18074	 => std_logic_vector(to_unsigned(109,8) ,
18075	 => std_logic_vector(to_unsigned(101,8) ,
18076	 => std_logic_vector(to_unsigned(88,8) ,
18077	 => std_logic_vector(to_unsigned(79,8) ,
18078	 => std_logic_vector(to_unsigned(85,8) ,
18079	 => std_logic_vector(to_unsigned(81,8) ,
18080	 => std_logic_vector(to_unsigned(80,8) ,
18081	 => std_logic_vector(to_unsigned(77,8) ,
18082	 => std_logic_vector(to_unsigned(82,8) ,
18083	 => std_logic_vector(to_unsigned(103,8) ,
18084	 => std_logic_vector(to_unsigned(118,8) ,
18085	 => std_logic_vector(to_unsigned(116,8) ,
18086	 => std_logic_vector(to_unsigned(93,8) ,
18087	 => std_logic_vector(to_unsigned(87,8) ,
18088	 => std_logic_vector(to_unsigned(78,8) ,
18089	 => std_logic_vector(to_unsigned(88,8) ,
18090	 => std_logic_vector(to_unsigned(78,8) ,
18091	 => std_logic_vector(to_unsigned(87,8) ,
18092	 => std_logic_vector(to_unsigned(119,8) ,
18093	 => std_logic_vector(to_unsigned(97,8) ,
18094	 => std_logic_vector(to_unsigned(108,8) ,
18095	 => std_logic_vector(to_unsigned(112,8) ,
18096	 => std_logic_vector(to_unsigned(97,8) ,
18097	 => std_logic_vector(to_unsigned(91,8) ,
18098	 => std_logic_vector(to_unsigned(104,8) ,
18099	 => std_logic_vector(to_unsigned(118,8) ,
18100	 => std_logic_vector(to_unsigned(125,8) ,
18101	 => std_logic_vector(to_unsigned(156,8) ,
18102	 => std_logic_vector(to_unsigned(139,8) ,
18103	 => std_logic_vector(to_unsigned(118,8) ,
18104	 => std_logic_vector(to_unsigned(90,8) ,
18105	 => std_logic_vector(to_unsigned(77,8) ,
18106	 => std_logic_vector(to_unsigned(87,8) ,
18107	 => std_logic_vector(to_unsigned(93,8) ,
18108	 => std_logic_vector(to_unsigned(99,8) ,
18109	 => std_logic_vector(to_unsigned(78,8) ,
18110	 => std_logic_vector(to_unsigned(56,8) ,
18111	 => std_logic_vector(to_unsigned(54,8) ,
18112	 => std_logic_vector(to_unsigned(51,8) ,
18113	 => std_logic_vector(to_unsigned(93,8) ,
18114	 => std_logic_vector(to_unsigned(142,8) ,
18115	 => std_logic_vector(to_unsigned(108,8) ,
18116	 => std_logic_vector(to_unsigned(80,8) ,
18117	 => std_logic_vector(to_unsigned(70,8) ,
18118	 => std_logic_vector(to_unsigned(79,8) ,
18119	 => std_logic_vector(to_unsigned(72,8) ,
18120	 => std_logic_vector(to_unsigned(58,8) ,
18121	 => std_logic_vector(to_unsigned(53,8) ,
18122	 => std_logic_vector(to_unsigned(68,8) ,
18123	 => std_logic_vector(to_unsigned(72,8) ,
18124	 => std_logic_vector(to_unsigned(65,8) ,
18125	 => std_logic_vector(to_unsigned(64,8) ,
18126	 => std_logic_vector(to_unsigned(60,8) ,
18127	 => std_logic_vector(to_unsigned(53,8) ,
18128	 => std_logic_vector(to_unsigned(57,8) ,
18129	 => std_logic_vector(to_unsigned(65,8) ,
18130	 => std_logic_vector(to_unsigned(66,8) ,
18131	 => std_logic_vector(to_unsigned(60,8) ,
18132	 => std_logic_vector(to_unsigned(62,8) ,
18133	 => std_logic_vector(to_unsigned(67,8) ,
18134	 => std_logic_vector(to_unsigned(70,8) ,
18135	 => std_logic_vector(to_unsigned(66,8) ,
18136	 => std_logic_vector(to_unsigned(64,8) ,
18137	 => std_logic_vector(to_unsigned(60,8) ,
18138	 => std_logic_vector(to_unsigned(58,8) ,
18139	 => std_logic_vector(to_unsigned(65,8) ,
18140	 => std_logic_vector(to_unsigned(67,8) ,
18141	 => std_logic_vector(to_unsigned(61,8) ,
18142	 => std_logic_vector(to_unsigned(67,8) ,
18143	 => std_logic_vector(to_unsigned(67,8) ,
18144	 => std_logic_vector(to_unsigned(63,8) ,
18145	 => std_logic_vector(to_unsigned(71,8) ,
18146	 => std_logic_vector(to_unsigned(79,8) ,
18147	 => std_logic_vector(to_unsigned(71,8) ,
18148	 => std_logic_vector(to_unsigned(68,8) ,
18149	 => std_logic_vector(to_unsigned(86,8) ,
18150	 => std_logic_vector(to_unsigned(82,8) ,
18151	 => std_logic_vector(to_unsigned(72,8) ,
18152	 => std_logic_vector(to_unsigned(69,8) ,
18153	 => std_logic_vector(to_unsigned(78,8) ,
18154	 => std_logic_vector(to_unsigned(85,8) ,
18155	 => std_logic_vector(to_unsigned(74,8) ,
18156	 => std_logic_vector(to_unsigned(84,8) ,
18157	 => std_logic_vector(to_unsigned(79,8) ,
18158	 => std_logic_vector(to_unsigned(68,8) ,
18159	 => std_logic_vector(to_unsigned(87,8) ,
18160	 => std_logic_vector(to_unsigned(103,8) ,
18161	 => std_logic_vector(to_unsigned(90,8) ,
18162	 => std_logic_vector(to_unsigned(80,8) ,
18163	 => std_logic_vector(to_unsigned(100,8) ,
18164	 => std_logic_vector(to_unsigned(130,8) ,
18165	 => std_logic_vector(to_unsigned(127,8) ,
18166	 => std_logic_vector(to_unsigned(128,8) ,
18167	 => std_logic_vector(to_unsigned(121,8) ,
18168	 => std_logic_vector(to_unsigned(144,8) ,
18169	 => std_logic_vector(to_unsigned(71,8) ,
18170	 => std_logic_vector(to_unsigned(1,8) ,
18171	 => std_logic_vector(to_unsigned(0,8) ,
18172	 => std_logic_vector(to_unsigned(7,8) ,
18173	 => std_logic_vector(to_unsigned(122,8) ,
18174	 => std_logic_vector(to_unsigned(133,8) ,
18175	 => std_logic_vector(to_unsigned(108,8) ,
18176	 => std_logic_vector(to_unsigned(100,8) ,
18177	 => std_logic_vector(to_unsigned(93,8) ,
18178	 => std_logic_vector(to_unsigned(99,8) ,
18179	 => std_logic_vector(to_unsigned(108,8) ,
18180	 => std_logic_vector(to_unsigned(107,8) ,
18181	 => std_logic_vector(to_unsigned(104,8) ,
18182	 => std_logic_vector(to_unsigned(107,8) ,
18183	 => std_logic_vector(to_unsigned(105,8) ,
18184	 => std_logic_vector(to_unsigned(96,8) ,
18185	 => std_logic_vector(to_unsigned(92,8) ,
18186	 => std_logic_vector(to_unsigned(95,8) ,
18187	 => std_logic_vector(to_unsigned(88,8) ,
18188	 => std_logic_vector(to_unsigned(82,8) ,
18189	 => std_logic_vector(to_unsigned(86,8) ,
18190	 => std_logic_vector(to_unsigned(82,8) ,
18191	 => std_logic_vector(to_unsigned(80,8) ,
18192	 => std_logic_vector(to_unsigned(79,8) ,
18193	 => std_logic_vector(to_unsigned(76,8) ,
18194	 => std_logic_vector(to_unsigned(84,8) ,
18195	 => std_logic_vector(to_unsigned(81,8) ,
18196	 => std_logic_vector(to_unsigned(72,8) ,
18197	 => std_logic_vector(to_unsigned(67,8) ,
18198	 => std_logic_vector(to_unsigned(62,8) ,
18199	 => std_logic_vector(to_unsigned(71,8) ,
18200	 => std_logic_vector(to_unsigned(77,8) ,
18201	 => std_logic_vector(to_unsigned(78,8) ,
18202	 => std_logic_vector(to_unsigned(70,8) ,
18203	 => std_logic_vector(to_unsigned(68,8) ,
18204	 => std_logic_vector(to_unsigned(72,8) ,
18205	 => std_logic_vector(to_unsigned(76,8) ,
18206	 => std_logic_vector(to_unsigned(81,8) ,
18207	 => std_logic_vector(to_unsigned(84,8) ,
18208	 => std_logic_vector(to_unsigned(82,8) ,
18209	 => std_logic_vector(to_unsigned(82,8) ,
18210	 => std_logic_vector(to_unsigned(79,8) ,
18211	 => std_logic_vector(to_unsigned(85,8) ,
18212	 => std_logic_vector(to_unsigned(90,8) ,
18213	 => std_logic_vector(to_unsigned(86,8) ,
18214	 => std_logic_vector(to_unsigned(86,8) ,
18215	 => std_logic_vector(to_unsigned(84,8) ,
18216	 => std_logic_vector(to_unsigned(86,8) ,
18217	 => std_logic_vector(to_unsigned(90,8) ,
18218	 => std_logic_vector(to_unsigned(95,8) ,
18219	 => std_logic_vector(to_unsigned(95,8) ,
18220	 => std_logic_vector(to_unsigned(85,8) ,
18221	 => std_logic_vector(to_unsigned(79,8) ,
18222	 => std_logic_vector(to_unsigned(85,8) ,
18223	 => std_logic_vector(to_unsigned(93,8) ,
18224	 => std_logic_vector(to_unsigned(90,8) ,
18225	 => std_logic_vector(to_unsigned(85,8) ,
18226	 => std_logic_vector(to_unsigned(80,8) ,
18227	 => std_logic_vector(to_unsigned(80,8) ,
18228	 => std_logic_vector(to_unsigned(87,8) ,
18229	 => std_logic_vector(to_unsigned(92,8) ,
18230	 => std_logic_vector(to_unsigned(87,8) ,
18231	 => std_logic_vector(to_unsigned(90,8) ,
18232	 => std_logic_vector(to_unsigned(88,8) ,
18233	 => std_logic_vector(to_unsigned(82,8) ,
18234	 => std_logic_vector(to_unsigned(90,8) ,
18235	 => std_logic_vector(to_unsigned(82,8) ,
18236	 => std_logic_vector(to_unsigned(84,8) ,
18237	 => std_logic_vector(to_unsigned(86,8) ,
18238	 => std_logic_vector(to_unsigned(85,8) ,
18239	 => std_logic_vector(to_unsigned(86,8) ,
18240	 => std_logic_vector(to_unsigned(86,8) ,
18241	 => std_logic_vector(to_unsigned(154,8) ,
18242	 => std_logic_vector(to_unsigned(157,8) ,
18243	 => std_logic_vector(to_unsigned(156,8) ,
18244	 => std_logic_vector(to_unsigned(154,8) ,
18245	 => std_logic_vector(to_unsigned(154,8) ,
18246	 => std_logic_vector(to_unsigned(157,8) ,
18247	 => std_logic_vector(to_unsigned(156,8) ,
18248	 => std_logic_vector(to_unsigned(156,8) ,
18249	 => std_logic_vector(to_unsigned(159,8) ,
18250	 => std_logic_vector(to_unsigned(159,8) ,
18251	 => std_logic_vector(to_unsigned(157,8) ,
18252	 => std_logic_vector(to_unsigned(163,8) ,
18253	 => std_logic_vector(to_unsigned(157,8) ,
18254	 => std_logic_vector(to_unsigned(156,8) ,
18255	 => std_logic_vector(to_unsigned(156,8) ,
18256	 => std_logic_vector(to_unsigned(157,8) ,
18257	 => std_logic_vector(to_unsigned(166,8) ,
18258	 => std_logic_vector(to_unsigned(175,8) ,
18259	 => std_logic_vector(to_unsigned(166,8) ,
18260	 => std_logic_vector(to_unsigned(175,8) ,
18261	 => std_logic_vector(to_unsigned(173,8) ,
18262	 => std_logic_vector(to_unsigned(157,8) ,
18263	 => std_logic_vector(to_unsigned(152,8) ,
18264	 => std_logic_vector(to_unsigned(151,8) ,
18265	 => std_logic_vector(to_unsigned(154,8) ,
18266	 => std_logic_vector(to_unsigned(171,8) ,
18267	 => std_logic_vector(to_unsigned(108,8) ,
18268	 => std_logic_vector(to_unsigned(13,8) ,
18269	 => std_logic_vector(to_unsigned(6,8) ,
18270	 => std_logic_vector(to_unsigned(4,8) ,
18271	 => std_logic_vector(to_unsigned(2,8) ,
18272	 => std_logic_vector(to_unsigned(6,8) ,
18273	 => std_logic_vector(to_unsigned(6,8) ,
18274	 => std_logic_vector(to_unsigned(6,8) ,
18275	 => std_logic_vector(to_unsigned(2,8) ,
18276	 => std_logic_vector(to_unsigned(42,8) ,
18277	 => std_logic_vector(to_unsigned(173,8) ,
18278	 => std_logic_vector(to_unsigned(156,8) ,
18279	 => std_logic_vector(to_unsigned(157,8) ,
18280	 => std_logic_vector(to_unsigned(159,8) ,
18281	 => std_logic_vector(to_unsigned(159,8) ,
18282	 => std_logic_vector(to_unsigned(161,8) ,
18283	 => std_logic_vector(to_unsigned(161,8) ,
18284	 => std_logic_vector(to_unsigned(159,8) ,
18285	 => std_logic_vector(to_unsigned(157,8) ,
18286	 => std_logic_vector(to_unsigned(159,8) ,
18287	 => std_logic_vector(to_unsigned(166,8) ,
18288	 => std_logic_vector(to_unsigned(154,8) ,
18289	 => std_logic_vector(to_unsigned(142,8) ,
18290	 => std_logic_vector(to_unsigned(152,8) ,
18291	 => std_logic_vector(to_unsigned(161,8) ,
18292	 => std_logic_vector(to_unsigned(144,8) ,
18293	 => std_logic_vector(to_unsigned(156,8) ,
18294	 => std_logic_vector(to_unsigned(127,8) ,
18295	 => std_logic_vector(to_unsigned(20,8) ,
18296	 => std_logic_vector(to_unsigned(41,8) ,
18297	 => std_logic_vector(to_unsigned(81,8) ,
18298	 => std_logic_vector(to_unsigned(74,8) ,
18299	 => std_logic_vector(to_unsigned(71,8) ,
18300	 => std_logic_vector(to_unsigned(85,8) ,
18301	 => std_logic_vector(to_unsigned(85,8) ,
18302	 => std_logic_vector(to_unsigned(49,8) ,
18303	 => std_logic_vector(to_unsigned(51,8) ,
18304	 => std_logic_vector(to_unsigned(44,8) ,
18305	 => std_logic_vector(to_unsigned(25,8) ,
18306	 => std_logic_vector(to_unsigned(49,8) ,
18307	 => std_logic_vector(to_unsigned(55,8) ,
18308	 => std_logic_vector(to_unsigned(42,8) ,
18309	 => std_logic_vector(to_unsigned(111,8) ,
18310	 => std_logic_vector(to_unsigned(175,8) ,
18311	 => std_logic_vector(to_unsigned(166,8) ,
18312	 => std_logic_vector(to_unsigned(166,8) ,
18313	 => std_logic_vector(to_unsigned(166,8) ,
18314	 => std_logic_vector(to_unsigned(163,8) ,
18315	 => std_logic_vector(to_unsigned(163,8) ,
18316	 => std_logic_vector(to_unsigned(161,8) ,
18317	 => std_logic_vector(to_unsigned(163,8) ,
18318	 => std_logic_vector(to_unsigned(164,8) ,
18319	 => std_logic_vector(to_unsigned(164,8) ,
18320	 => std_logic_vector(to_unsigned(159,8) ,
18321	 => std_logic_vector(to_unsigned(157,8) ,
18322	 => std_logic_vector(to_unsigned(157,8) ,
18323	 => std_logic_vector(to_unsigned(157,8) ,
18324	 => std_logic_vector(to_unsigned(159,8) ,
18325	 => std_logic_vector(to_unsigned(173,8) ,
18326	 => std_logic_vector(to_unsigned(96,8) ,
18327	 => std_logic_vector(to_unsigned(4,8) ,
18328	 => std_logic_vector(to_unsigned(11,8) ,
18329	 => std_logic_vector(to_unsigned(48,8) ,
18330	 => std_logic_vector(to_unsigned(3,8) ,
18331	 => std_logic_vector(to_unsigned(0,8) ,
18332	 => std_logic_vector(to_unsigned(1,8) ,
18333	 => std_logic_vector(to_unsigned(1,8) ,
18334	 => std_logic_vector(to_unsigned(1,8) ,
18335	 => std_logic_vector(to_unsigned(1,8) ,
18336	 => std_logic_vector(to_unsigned(1,8) ,
18337	 => std_logic_vector(to_unsigned(1,8) ,
18338	 => std_logic_vector(to_unsigned(2,8) ,
18339	 => std_logic_vector(to_unsigned(1,8) ,
18340	 => std_logic_vector(to_unsigned(1,8) ,
18341	 => std_logic_vector(to_unsigned(1,8) ,
18342	 => std_logic_vector(to_unsigned(74,8) ,
18343	 => std_logic_vector(to_unsigned(196,8) ,
18344	 => std_logic_vector(to_unsigned(161,8) ,
18345	 => std_logic_vector(to_unsigned(170,8) ,
18346	 => std_logic_vector(to_unsigned(171,8) ,
18347	 => std_logic_vector(to_unsigned(170,8) ,
18348	 => std_logic_vector(to_unsigned(170,8) ,
18349	 => std_logic_vector(to_unsigned(164,8) ,
18350	 => std_logic_vector(to_unsigned(159,8) ,
18351	 => std_logic_vector(to_unsigned(159,8) ,
18352	 => std_logic_vector(to_unsigned(156,8) ,
18353	 => std_logic_vector(to_unsigned(156,8) ,
18354	 => std_logic_vector(to_unsigned(156,8) ,
18355	 => std_logic_vector(to_unsigned(154,8) ,
18356	 => std_logic_vector(to_unsigned(157,8) ,
18357	 => std_logic_vector(to_unsigned(168,8) ,
18358	 => std_logic_vector(to_unsigned(166,8) ,
18359	 => std_logic_vector(to_unsigned(152,8) ,
18360	 => std_logic_vector(to_unsigned(147,8) ,
18361	 => std_logic_vector(to_unsigned(144,8) ,
18362	 => std_logic_vector(to_unsigned(149,8) ,
18363	 => std_logic_vector(to_unsigned(149,8) ,
18364	 => std_logic_vector(to_unsigned(161,8) ,
18365	 => std_logic_vector(to_unsigned(168,8) ,
18366	 => std_logic_vector(to_unsigned(159,8) ,
18367	 => std_logic_vector(to_unsigned(141,8) ,
18368	 => std_logic_vector(to_unsigned(138,8) ,
18369	 => std_logic_vector(to_unsigned(127,8) ,
18370	 => std_logic_vector(to_unsigned(118,8) ,
18371	 => std_logic_vector(to_unsigned(118,8) ,
18372	 => std_logic_vector(to_unsigned(122,8) ,
18373	 => std_logic_vector(to_unsigned(109,8) ,
18374	 => std_logic_vector(to_unsigned(107,8) ,
18375	 => std_logic_vector(to_unsigned(134,8) ,
18376	 => std_logic_vector(to_unsigned(133,8) ,
18377	 => std_logic_vector(to_unsigned(121,8) ,
18378	 => std_logic_vector(to_unsigned(115,8) ,
18379	 => std_logic_vector(to_unsigned(111,8) ,
18380	 => std_logic_vector(to_unsigned(105,8) ,
18381	 => std_logic_vector(to_unsigned(109,8) ,
18382	 => std_logic_vector(to_unsigned(116,8) ,
18383	 => std_logic_vector(to_unsigned(119,8) ,
18384	 => std_logic_vector(to_unsigned(109,8) ,
18385	 => std_logic_vector(to_unsigned(105,8) ,
18386	 => std_logic_vector(to_unsigned(127,8) ,
18387	 => std_logic_vector(to_unsigned(115,8) ,
18388	 => std_logic_vector(to_unsigned(114,8) ,
18389	 => std_logic_vector(to_unsigned(122,8) ,
18390	 => std_logic_vector(to_unsigned(103,8) ,
18391	 => std_logic_vector(to_unsigned(97,8) ,
18392	 => std_logic_vector(to_unsigned(112,8) ,
18393	 => std_logic_vector(to_unsigned(138,8) ,
18394	 => std_logic_vector(to_unsigned(121,8) ,
18395	 => std_logic_vector(to_unsigned(121,8) ,
18396	 => std_logic_vector(to_unsigned(104,8) ,
18397	 => std_logic_vector(to_unsigned(85,8) ,
18398	 => std_logic_vector(to_unsigned(80,8) ,
18399	 => std_logic_vector(to_unsigned(73,8) ,
18400	 => std_logic_vector(to_unsigned(71,8) ,
18401	 => std_logic_vector(to_unsigned(81,8) ,
18402	 => std_logic_vector(to_unsigned(91,8) ,
18403	 => std_logic_vector(to_unsigned(108,8) ,
18404	 => std_logic_vector(to_unsigned(74,8) ,
18405	 => std_logic_vector(to_unsigned(68,8) ,
18406	 => std_logic_vector(to_unsigned(91,8) ,
18407	 => std_logic_vector(to_unsigned(77,8) ,
18408	 => std_logic_vector(to_unsigned(46,8) ,
18409	 => std_logic_vector(to_unsigned(53,8) ,
18410	 => std_logic_vector(to_unsigned(57,8) ,
18411	 => std_logic_vector(to_unsigned(78,8) ,
18412	 => std_logic_vector(to_unsigned(105,8) ,
18413	 => std_logic_vector(to_unsigned(97,8) ,
18414	 => std_logic_vector(to_unsigned(76,8) ,
18415	 => std_logic_vector(to_unsigned(77,8) ,
18416	 => std_logic_vector(to_unsigned(103,8) ,
18417	 => std_logic_vector(to_unsigned(100,8) ,
18418	 => std_logic_vector(to_unsigned(97,8) ,
18419	 => std_logic_vector(to_unsigned(111,8) ,
18420	 => std_logic_vector(to_unsigned(125,8) ,
18421	 => std_logic_vector(to_unsigned(151,8) ,
18422	 => std_logic_vector(to_unsigned(141,8) ,
18423	 => std_logic_vector(to_unsigned(121,8) ,
18424	 => std_logic_vector(to_unsigned(91,8) ,
18425	 => std_logic_vector(to_unsigned(87,8) ,
18426	 => std_logic_vector(to_unsigned(109,8) ,
18427	 => std_logic_vector(to_unsigned(111,8) ,
18428	 => std_logic_vector(to_unsigned(85,8) ,
18429	 => std_logic_vector(to_unsigned(44,8) ,
18430	 => std_logic_vector(to_unsigned(44,8) ,
18431	 => std_logic_vector(to_unsigned(53,8) ,
18432	 => std_logic_vector(to_unsigned(49,8) ,
18433	 => std_logic_vector(to_unsigned(60,8) ,
18434	 => std_logic_vector(to_unsigned(88,8) ,
18435	 => std_logic_vector(to_unsigned(84,8) ,
18436	 => std_logic_vector(to_unsigned(66,8) ,
18437	 => std_logic_vector(to_unsigned(73,8) ,
18438	 => std_logic_vector(to_unsigned(79,8) ,
18439	 => std_logic_vector(to_unsigned(70,8) ,
18440	 => std_logic_vector(to_unsigned(61,8) ,
18441	 => std_logic_vector(to_unsigned(52,8) ,
18442	 => std_logic_vector(to_unsigned(58,8) ,
18443	 => std_logic_vector(to_unsigned(71,8) ,
18444	 => std_logic_vector(to_unsigned(61,8) ,
18445	 => std_logic_vector(to_unsigned(57,8) ,
18446	 => std_logic_vector(to_unsigned(53,8) ,
18447	 => std_logic_vector(to_unsigned(49,8) ,
18448	 => std_logic_vector(to_unsigned(61,8) ,
18449	 => std_logic_vector(to_unsigned(58,8) ,
18450	 => std_logic_vector(to_unsigned(56,8) ,
18451	 => std_logic_vector(to_unsigned(59,8) ,
18452	 => std_logic_vector(to_unsigned(62,8) ,
18453	 => std_logic_vector(to_unsigned(64,8) ,
18454	 => std_logic_vector(to_unsigned(59,8) ,
18455	 => std_logic_vector(to_unsigned(61,8) ,
18456	 => std_logic_vector(to_unsigned(57,8) ,
18457	 => std_logic_vector(to_unsigned(52,8) ,
18458	 => std_logic_vector(to_unsigned(55,8) ,
18459	 => std_logic_vector(to_unsigned(58,8) ,
18460	 => std_logic_vector(to_unsigned(61,8) ,
18461	 => std_logic_vector(to_unsigned(65,8) ,
18462	 => std_logic_vector(to_unsigned(68,8) ,
18463	 => std_logic_vector(to_unsigned(68,8) ,
18464	 => std_logic_vector(to_unsigned(69,8) ,
18465	 => std_logic_vector(to_unsigned(74,8) ,
18466	 => std_logic_vector(to_unsigned(78,8) ,
18467	 => std_logic_vector(to_unsigned(72,8) ,
18468	 => std_logic_vector(to_unsigned(62,8) ,
18469	 => std_logic_vector(to_unsigned(80,8) ,
18470	 => std_logic_vector(to_unsigned(84,8) ,
18471	 => std_logic_vector(to_unsigned(81,8) ,
18472	 => std_logic_vector(to_unsigned(81,8) ,
18473	 => std_logic_vector(to_unsigned(90,8) ,
18474	 => std_logic_vector(to_unsigned(90,8) ,
18475	 => std_logic_vector(to_unsigned(85,8) ,
18476	 => std_logic_vector(to_unsigned(87,8) ,
18477	 => std_logic_vector(to_unsigned(91,8) ,
18478	 => std_logic_vector(to_unsigned(86,8) ,
18479	 => std_logic_vector(to_unsigned(97,8) ,
18480	 => std_logic_vector(to_unsigned(112,8) ,
18481	 => std_logic_vector(to_unsigned(91,8) ,
18482	 => std_logic_vector(to_unsigned(99,8) ,
18483	 => std_logic_vector(to_unsigned(124,8) ,
18484	 => std_logic_vector(to_unsigned(125,8) ,
18485	 => std_logic_vector(to_unsigned(128,8) ,
18486	 => std_logic_vector(to_unsigned(133,8) ,
18487	 => std_logic_vector(to_unsigned(131,8) ,
18488	 => std_logic_vector(to_unsigned(142,8) ,
18489	 => std_logic_vector(to_unsigned(103,8) ,
18490	 => std_logic_vector(to_unsigned(6,8) ,
18491	 => std_logic_vector(to_unsigned(0,8) ,
18492	 => std_logic_vector(to_unsigned(3,8) ,
18493	 => std_logic_vector(to_unsigned(100,8) ,
18494	 => std_logic_vector(to_unsigned(161,8) ,
18495	 => std_logic_vector(to_unsigned(136,8) ,
18496	 => std_logic_vector(to_unsigned(131,8) ,
18497	 => std_logic_vector(to_unsigned(116,8) ,
18498	 => std_logic_vector(to_unsigned(127,8) ,
18499	 => std_logic_vector(to_unsigned(134,8) ,
18500	 => std_logic_vector(to_unsigned(134,8) ,
18501	 => std_logic_vector(to_unsigned(119,8) ,
18502	 => std_logic_vector(to_unsigned(99,8) ,
18503	 => std_logic_vector(to_unsigned(93,8) ,
18504	 => std_logic_vector(to_unsigned(93,8) ,
18505	 => std_logic_vector(to_unsigned(85,8) ,
18506	 => std_logic_vector(to_unsigned(82,8) ,
18507	 => std_logic_vector(to_unsigned(86,8) ,
18508	 => std_logic_vector(to_unsigned(84,8) ,
18509	 => std_logic_vector(to_unsigned(84,8) ,
18510	 => std_logic_vector(to_unsigned(82,8) ,
18511	 => std_logic_vector(to_unsigned(86,8) ,
18512	 => std_logic_vector(to_unsigned(84,8) ,
18513	 => std_logic_vector(to_unsigned(76,8) ,
18514	 => std_logic_vector(to_unsigned(79,8) ,
18515	 => std_logic_vector(to_unsigned(82,8) ,
18516	 => std_logic_vector(to_unsigned(81,8) ,
18517	 => std_logic_vector(to_unsigned(79,8) ,
18518	 => std_logic_vector(to_unsigned(61,8) ,
18519	 => std_logic_vector(to_unsigned(58,8) ,
18520	 => std_logic_vector(to_unsigned(68,8) ,
18521	 => std_logic_vector(to_unsigned(69,8) ,
18522	 => std_logic_vector(to_unsigned(66,8) ,
18523	 => std_logic_vector(to_unsigned(74,8) ,
18524	 => std_logic_vector(to_unsigned(74,8) ,
18525	 => std_logic_vector(to_unsigned(81,8) ,
18526	 => std_logic_vector(to_unsigned(81,8) ,
18527	 => std_logic_vector(to_unsigned(82,8) ,
18528	 => std_logic_vector(to_unsigned(82,8) ,
18529	 => std_logic_vector(to_unsigned(76,8) ,
18530	 => std_logic_vector(to_unsigned(76,8) ,
18531	 => std_logic_vector(to_unsigned(82,8) ,
18532	 => std_logic_vector(to_unsigned(90,8) ,
18533	 => std_logic_vector(to_unsigned(88,8) ,
18534	 => std_logic_vector(to_unsigned(81,8) ,
18535	 => std_logic_vector(to_unsigned(88,8) ,
18536	 => std_logic_vector(to_unsigned(97,8) ,
18537	 => std_logic_vector(to_unsigned(91,8) ,
18538	 => std_logic_vector(to_unsigned(92,8) ,
18539	 => std_logic_vector(to_unsigned(100,8) ,
18540	 => std_logic_vector(to_unsigned(93,8) ,
18541	 => std_logic_vector(to_unsigned(87,8) ,
18542	 => std_logic_vector(to_unsigned(87,8) ,
18543	 => std_logic_vector(to_unsigned(87,8) ,
18544	 => std_logic_vector(to_unsigned(95,8) ,
18545	 => std_logic_vector(to_unsigned(92,8) ,
18546	 => std_logic_vector(to_unsigned(86,8) ,
18547	 => std_logic_vector(to_unsigned(90,8) ,
18548	 => std_logic_vector(to_unsigned(96,8) ,
18549	 => std_logic_vector(to_unsigned(101,8) ,
18550	 => std_logic_vector(to_unsigned(99,8) ,
18551	 => std_logic_vector(to_unsigned(91,8) ,
18552	 => std_logic_vector(to_unsigned(81,8) ,
18553	 => std_logic_vector(to_unsigned(78,8) ,
18554	 => std_logic_vector(to_unsigned(86,8) ,
18555	 => std_logic_vector(to_unsigned(85,8) ,
18556	 => std_logic_vector(to_unsigned(86,8) ,
18557	 => std_logic_vector(to_unsigned(88,8) ,
18558	 => std_logic_vector(to_unsigned(84,8) ,
18559	 => std_logic_vector(to_unsigned(80,8) ,
18560	 => std_logic_vector(to_unsigned(79,8) ,
18561	 => std_logic_vector(to_unsigned(157,8) ,
18562	 => std_logic_vector(to_unsigned(154,8) ,
18563	 => std_logic_vector(to_unsigned(154,8) ,
18564	 => std_logic_vector(to_unsigned(154,8) ,
18565	 => std_logic_vector(to_unsigned(154,8) ,
18566	 => std_logic_vector(to_unsigned(159,8) ,
18567	 => std_logic_vector(to_unsigned(156,8) ,
18568	 => std_logic_vector(to_unsigned(154,8) ,
18569	 => std_logic_vector(to_unsigned(154,8) ,
18570	 => std_logic_vector(to_unsigned(154,8) ,
18571	 => std_logic_vector(to_unsigned(152,8) ,
18572	 => std_logic_vector(to_unsigned(159,8) ,
18573	 => std_logic_vector(to_unsigned(159,8) ,
18574	 => std_logic_vector(to_unsigned(157,8) ,
18575	 => std_logic_vector(to_unsigned(171,8) ,
18576	 => std_logic_vector(to_unsigned(175,8) ,
18577	 => std_logic_vector(to_unsigned(138,8) ,
18578	 => std_logic_vector(to_unsigned(68,8) ,
18579	 => std_logic_vector(to_unsigned(45,8) ,
18580	 => std_logic_vector(to_unsigned(73,8) ,
18581	 => std_logic_vector(to_unsigned(112,8) ,
18582	 => std_logic_vector(to_unsigned(170,8) ,
18583	 => std_logic_vector(to_unsigned(164,8) ,
18584	 => std_logic_vector(to_unsigned(149,8) ,
18585	 => std_logic_vector(to_unsigned(186,8) ,
18586	 => std_logic_vector(to_unsigned(101,8) ,
18587	 => std_logic_vector(to_unsigned(11,8) ,
18588	 => std_logic_vector(to_unsigned(5,8) ,
18589	 => std_logic_vector(to_unsigned(8,8) ,
18590	 => std_logic_vector(to_unsigned(4,8) ,
18591	 => std_logic_vector(to_unsigned(5,8) ,
18592	 => std_logic_vector(to_unsigned(12,8) ,
18593	 => std_logic_vector(to_unsigned(12,8) ,
18594	 => std_logic_vector(to_unsigned(5,8) ,
18595	 => std_logic_vector(to_unsigned(1,8) ,
18596	 => std_logic_vector(to_unsigned(12,8) ,
18597	 => std_logic_vector(to_unsigned(142,8) ,
18598	 => std_logic_vector(to_unsigned(166,8) ,
18599	 => std_logic_vector(to_unsigned(154,8) ,
18600	 => std_logic_vector(to_unsigned(159,8) ,
18601	 => std_logic_vector(to_unsigned(161,8) ,
18602	 => std_logic_vector(to_unsigned(157,8) ,
18603	 => std_logic_vector(to_unsigned(159,8) ,
18604	 => std_logic_vector(to_unsigned(164,8) ,
18605	 => std_logic_vector(to_unsigned(161,8) ,
18606	 => std_logic_vector(to_unsigned(157,8) ,
18607	 => std_logic_vector(to_unsigned(163,8) ,
18608	 => std_logic_vector(to_unsigned(156,8) ,
18609	 => std_logic_vector(to_unsigned(146,8) ,
18610	 => std_logic_vector(to_unsigned(157,8) ,
18611	 => std_logic_vector(to_unsigned(157,8) ,
18612	 => std_logic_vector(to_unsigned(154,8) ,
18613	 => std_logic_vector(to_unsigned(170,8) ,
18614	 => std_logic_vector(to_unsigned(107,8) ,
18615	 => std_logic_vector(to_unsigned(28,8) ,
18616	 => std_logic_vector(to_unsigned(60,8) ,
18617	 => std_logic_vector(to_unsigned(55,8) ,
18618	 => std_logic_vector(to_unsigned(52,8) ,
18619	 => std_logic_vector(to_unsigned(65,8) ,
18620	 => std_logic_vector(to_unsigned(73,8) ,
18621	 => std_logic_vector(to_unsigned(60,8) ,
18622	 => std_logic_vector(to_unsigned(41,8) ,
18623	 => std_logic_vector(to_unsigned(43,8) ,
18624	 => std_logic_vector(to_unsigned(48,8) ,
18625	 => std_logic_vector(to_unsigned(39,8) ,
18626	 => std_logic_vector(to_unsigned(35,8) ,
18627	 => std_logic_vector(to_unsigned(54,8) ,
18628	 => std_logic_vector(to_unsigned(36,8) ,
18629	 => std_logic_vector(to_unsigned(105,8) ,
18630	 => std_logic_vector(to_unsigned(183,8) ,
18631	 => std_logic_vector(to_unsigned(164,8) ,
18632	 => std_logic_vector(to_unsigned(166,8) ,
18633	 => std_logic_vector(to_unsigned(164,8) ,
18634	 => std_logic_vector(to_unsigned(163,8) ,
18635	 => std_logic_vector(to_unsigned(164,8) ,
18636	 => std_logic_vector(to_unsigned(164,8) ,
18637	 => std_logic_vector(to_unsigned(161,8) ,
18638	 => std_logic_vector(to_unsigned(157,8) ,
18639	 => std_logic_vector(to_unsigned(161,8) ,
18640	 => std_logic_vector(to_unsigned(163,8) ,
18641	 => std_logic_vector(to_unsigned(161,8) ,
18642	 => std_logic_vector(to_unsigned(159,8) ,
18643	 => std_logic_vector(to_unsigned(161,8) ,
18644	 => std_logic_vector(to_unsigned(159,8) ,
18645	 => std_logic_vector(to_unsigned(175,8) ,
18646	 => std_logic_vector(to_unsigned(97,8) ,
18647	 => std_logic_vector(to_unsigned(7,8) ,
18648	 => std_logic_vector(to_unsigned(3,8) ,
18649	 => std_logic_vector(to_unsigned(7,8) ,
18650	 => std_logic_vector(to_unsigned(2,8) ,
18651	 => std_logic_vector(to_unsigned(1,8) ,
18652	 => std_logic_vector(to_unsigned(1,8) ,
18653	 => std_logic_vector(to_unsigned(2,8) ,
18654	 => std_logic_vector(to_unsigned(2,8) ,
18655	 => std_logic_vector(to_unsigned(1,8) ,
18656	 => std_logic_vector(to_unsigned(1,8) ,
18657	 => std_logic_vector(to_unsigned(1,8) ,
18658	 => std_logic_vector(to_unsigned(1,8) ,
18659	 => std_logic_vector(to_unsigned(1,8) ,
18660	 => std_logic_vector(to_unsigned(1,8) ,
18661	 => std_logic_vector(to_unsigned(5,8) ,
18662	 => std_logic_vector(to_unsigned(128,8) ,
18663	 => std_logic_vector(to_unsigned(192,8) ,
18664	 => std_logic_vector(to_unsigned(166,8) ,
18665	 => std_logic_vector(to_unsigned(175,8) ,
18666	 => std_logic_vector(to_unsigned(171,8) ,
18667	 => std_logic_vector(to_unsigned(171,8) ,
18668	 => std_logic_vector(to_unsigned(170,8) ,
18669	 => std_logic_vector(to_unsigned(164,8) ,
18670	 => std_logic_vector(to_unsigned(161,8) ,
18671	 => std_logic_vector(to_unsigned(159,8) ,
18672	 => std_logic_vector(to_unsigned(157,8) ,
18673	 => std_logic_vector(to_unsigned(152,8) ,
18674	 => std_logic_vector(to_unsigned(149,8) ,
18675	 => std_logic_vector(to_unsigned(159,8) ,
18676	 => std_logic_vector(to_unsigned(161,8) ,
18677	 => std_logic_vector(to_unsigned(168,8) ,
18678	 => std_logic_vector(to_unsigned(171,8) ,
18679	 => std_logic_vector(to_unsigned(161,8) ,
18680	 => std_logic_vector(to_unsigned(159,8) ,
18681	 => std_logic_vector(to_unsigned(166,8) ,
18682	 => std_logic_vector(to_unsigned(170,8) ,
18683	 => std_logic_vector(to_unsigned(168,8) ,
18684	 => std_logic_vector(to_unsigned(161,8) ,
18685	 => std_logic_vector(to_unsigned(164,8) ,
18686	 => std_logic_vector(to_unsigned(164,8) ,
18687	 => std_logic_vector(to_unsigned(146,8) ,
18688	 => std_logic_vector(to_unsigned(125,8) ,
18689	 => std_logic_vector(to_unsigned(109,8) ,
18690	 => std_logic_vector(to_unsigned(112,8) ,
18691	 => std_logic_vector(to_unsigned(107,8) ,
18692	 => std_logic_vector(to_unsigned(100,8) ,
18693	 => std_logic_vector(to_unsigned(107,8) ,
18694	 => std_logic_vector(to_unsigned(121,8) ,
18695	 => std_logic_vector(to_unsigned(119,8) ,
18696	 => std_logic_vector(to_unsigned(112,8) ,
18697	 => std_logic_vector(to_unsigned(112,8) ,
18698	 => std_logic_vector(to_unsigned(121,8) ,
18699	 => std_logic_vector(to_unsigned(115,8) ,
18700	 => std_logic_vector(to_unsigned(107,8) ,
18701	 => std_logic_vector(to_unsigned(115,8) ,
18702	 => std_logic_vector(to_unsigned(116,8) ,
18703	 => std_logic_vector(to_unsigned(127,8) ,
18704	 => std_logic_vector(to_unsigned(122,8) ,
18705	 => std_logic_vector(to_unsigned(127,8) ,
18706	 => std_logic_vector(to_unsigned(144,8) ,
18707	 => std_logic_vector(to_unsigned(122,8) ,
18708	 => std_logic_vector(to_unsigned(133,8) ,
18709	 => std_logic_vector(to_unsigned(141,8) ,
18710	 => std_logic_vector(to_unsigned(127,8) ,
18711	 => std_logic_vector(to_unsigned(122,8) ,
18712	 => std_logic_vector(to_unsigned(131,8) ,
18713	 => std_logic_vector(to_unsigned(151,8) ,
18714	 => std_logic_vector(to_unsigned(152,8) ,
18715	 => std_logic_vector(to_unsigned(151,8) ,
18716	 => std_logic_vector(to_unsigned(111,8) ,
18717	 => std_logic_vector(to_unsigned(87,8) ,
18718	 => std_logic_vector(to_unsigned(77,8) ,
18719	 => std_logic_vector(to_unsigned(78,8) ,
18720	 => std_logic_vector(to_unsigned(84,8) ,
18721	 => std_logic_vector(to_unsigned(79,8) ,
18722	 => std_logic_vector(to_unsigned(100,8) ,
18723	 => std_logic_vector(to_unsigned(72,8) ,
18724	 => std_logic_vector(to_unsigned(20,8) ,
18725	 => std_logic_vector(to_unsigned(56,8) ,
18726	 => std_logic_vector(to_unsigned(95,8) ,
18727	 => std_logic_vector(to_unsigned(49,8) ,
18728	 => std_logic_vector(to_unsigned(25,8) ,
18729	 => std_logic_vector(to_unsigned(59,8) ,
18730	 => std_logic_vector(to_unsigned(27,8) ,
18731	 => std_logic_vector(to_unsigned(31,8) ,
18732	 => std_logic_vector(to_unsigned(71,8) ,
18733	 => std_logic_vector(to_unsigned(121,8) ,
18734	 => std_logic_vector(to_unsigned(92,8) ,
18735	 => std_logic_vector(to_unsigned(63,8) ,
18736	 => std_logic_vector(to_unsigned(86,8) ,
18737	 => std_logic_vector(to_unsigned(114,8) ,
18738	 => std_logic_vector(to_unsigned(108,8) ,
18739	 => std_logic_vector(to_unsigned(122,8) ,
18740	 => std_logic_vector(to_unsigned(138,8) ,
18741	 => std_logic_vector(to_unsigned(154,8) ,
18742	 => std_logic_vector(to_unsigned(144,8) ,
18743	 => std_logic_vector(to_unsigned(133,8) ,
18744	 => std_logic_vector(to_unsigned(108,8) ,
18745	 => std_logic_vector(to_unsigned(88,8) ,
18746	 => std_logic_vector(to_unsigned(95,8) ,
18747	 => std_logic_vector(to_unsigned(103,8) ,
18748	 => std_logic_vector(to_unsigned(77,8) ,
18749	 => std_logic_vector(to_unsigned(48,8) ,
18750	 => std_logic_vector(to_unsigned(53,8) ,
18751	 => std_logic_vector(to_unsigned(56,8) ,
18752	 => std_logic_vector(to_unsigned(54,8) ,
18753	 => std_logic_vector(to_unsigned(53,8) ,
18754	 => std_logic_vector(to_unsigned(70,8) ,
18755	 => std_logic_vector(to_unsigned(84,8) ,
18756	 => std_logic_vector(to_unsigned(76,8) ,
18757	 => std_logic_vector(to_unsigned(76,8) ,
18758	 => std_logic_vector(to_unsigned(79,8) ,
18759	 => std_logic_vector(to_unsigned(70,8) ,
18760	 => std_logic_vector(to_unsigned(53,8) ,
18761	 => std_logic_vector(to_unsigned(51,8) ,
18762	 => std_logic_vector(to_unsigned(68,8) ,
18763	 => std_logic_vector(to_unsigned(76,8) ,
18764	 => std_logic_vector(to_unsigned(59,8) ,
18765	 => std_logic_vector(to_unsigned(55,8) ,
18766	 => std_logic_vector(to_unsigned(61,8) ,
18767	 => std_logic_vector(to_unsigned(53,8) ,
18768	 => std_logic_vector(to_unsigned(61,8) ,
18769	 => std_logic_vector(to_unsigned(62,8) ,
18770	 => std_logic_vector(to_unsigned(49,8) ,
18771	 => std_logic_vector(to_unsigned(47,8) ,
18772	 => std_logic_vector(to_unsigned(64,8) ,
18773	 => std_logic_vector(to_unsigned(78,8) ,
18774	 => std_logic_vector(to_unsigned(58,8) ,
18775	 => std_logic_vector(to_unsigned(57,8) ,
18776	 => std_logic_vector(to_unsigned(58,8) ,
18777	 => std_logic_vector(to_unsigned(57,8) ,
18778	 => std_logic_vector(to_unsigned(59,8) ,
18779	 => std_logic_vector(to_unsigned(62,8) ,
18780	 => std_logic_vector(to_unsigned(62,8) ,
18781	 => std_logic_vector(to_unsigned(64,8) ,
18782	 => std_logic_vector(to_unsigned(64,8) ,
18783	 => std_logic_vector(to_unsigned(65,8) ,
18784	 => std_logic_vector(to_unsigned(73,8) ,
18785	 => std_logic_vector(to_unsigned(77,8) ,
18786	 => std_logic_vector(to_unsigned(65,8) ,
18787	 => std_logic_vector(to_unsigned(55,8) ,
18788	 => std_logic_vector(to_unsigned(58,8) ,
18789	 => std_logic_vector(to_unsigned(66,8) ,
18790	 => std_logic_vector(to_unsigned(87,8) ,
18791	 => std_logic_vector(to_unsigned(107,8) ,
18792	 => std_logic_vector(to_unsigned(92,8) ,
18793	 => std_logic_vector(to_unsigned(79,8) ,
18794	 => std_logic_vector(to_unsigned(90,8) ,
18795	 => std_logic_vector(to_unsigned(92,8) ,
18796	 => std_logic_vector(to_unsigned(86,8) ,
18797	 => std_logic_vector(to_unsigned(87,8) ,
18798	 => std_logic_vector(to_unsigned(95,8) ,
18799	 => std_logic_vector(to_unsigned(111,8) ,
18800	 => std_logic_vector(to_unsigned(119,8) ,
18801	 => std_logic_vector(to_unsigned(111,8) ,
18802	 => std_logic_vector(to_unsigned(119,8) ,
18803	 => std_logic_vector(to_unsigned(134,8) ,
18804	 => std_logic_vector(to_unsigned(138,8) ,
18805	 => std_logic_vector(to_unsigned(136,8) ,
18806	 => std_logic_vector(to_unsigned(141,8) ,
18807	 => std_logic_vector(to_unsigned(131,8) ,
18808	 => std_logic_vector(to_unsigned(136,8) ,
18809	 => std_logic_vector(to_unsigned(138,8) ,
18810	 => std_logic_vector(to_unsigned(24,8) ,
18811	 => std_logic_vector(to_unsigned(0,8) ,
18812	 => std_logic_vector(to_unsigned(1,8) ,
18813	 => std_logic_vector(to_unsigned(71,8) ,
18814	 => std_logic_vector(to_unsigned(175,8) ,
18815	 => std_logic_vector(to_unsigned(149,8) ,
18816	 => std_logic_vector(to_unsigned(152,8) ,
18817	 => std_logic_vector(to_unsigned(139,8) ,
18818	 => std_logic_vector(to_unsigned(151,8) ,
18819	 => std_logic_vector(to_unsigned(159,8) ,
18820	 => std_logic_vector(to_unsigned(151,8) ,
18821	 => std_logic_vector(to_unsigned(131,8) ,
18822	 => std_logic_vector(to_unsigned(109,8) ,
18823	 => std_logic_vector(to_unsigned(99,8) ,
18824	 => std_logic_vector(to_unsigned(99,8) ,
18825	 => std_logic_vector(to_unsigned(87,8) ,
18826	 => std_logic_vector(to_unsigned(78,8) ,
18827	 => std_logic_vector(to_unsigned(82,8) ,
18828	 => std_logic_vector(to_unsigned(85,8) ,
18829	 => std_logic_vector(to_unsigned(84,8) ,
18830	 => std_logic_vector(to_unsigned(80,8) ,
18831	 => std_logic_vector(to_unsigned(81,8) ,
18832	 => std_logic_vector(to_unsigned(79,8) ,
18833	 => std_logic_vector(to_unsigned(74,8) ,
18834	 => std_logic_vector(to_unsigned(86,8) ,
18835	 => std_logic_vector(to_unsigned(103,8) ,
18836	 => std_logic_vector(to_unsigned(124,8) ,
18837	 => std_logic_vector(to_unsigned(93,8) ,
18838	 => std_logic_vector(to_unsigned(58,8) ,
18839	 => std_logic_vector(to_unsigned(55,8) ,
18840	 => std_logic_vector(to_unsigned(64,8) ,
18841	 => std_logic_vector(to_unsigned(60,8) ,
18842	 => std_logic_vector(to_unsigned(66,8) ,
18843	 => std_logic_vector(to_unsigned(79,8) ,
18844	 => std_logic_vector(to_unsigned(86,8) ,
18845	 => std_logic_vector(to_unsigned(78,8) ,
18846	 => std_logic_vector(to_unsigned(85,8) ,
18847	 => std_logic_vector(to_unsigned(82,8) ,
18848	 => std_logic_vector(to_unsigned(91,8) ,
18849	 => std_logic_vector(to_unsigned(95,8) ,
18850	 => std_logic_vector(to_unsigned(86,8) ,
18851	 => std_logic_vector(to_unsigned(85,8) ,
18852	 => std_logic_vector(to_unsigned(92,8) ,
18853	 => std_logic_vector(to_unsigned(91,8) ,
18854	 => std_logic_vector(to_unsigned(87,8) ,
18855	 => std_logic_vector(to_unsigned(92,8) ,
18856	 => std_logic_vector(to_unsigned(99,8) ,
18857	 => std_logic_vector(to_unsigned(97,8) ,
18858	 => std_logic_vector(to_unsigned(105,8) ,
18859	 => std_logic_vector(to_unsigned(108,8) ,
18860	 => std_logic_vector(to_unsigned(101,8) ,
18861	 => std_logic_vector(to_unsigned(115,8) ,
18862	 => std_logic_vector(to_unsigned(131,8) ,
18863	 => std_logic_vector(to_unsigned(96,8) ,
18864	 => std_logic_vector(to_unsigned(84,8) ,
18865	 => std_logic_vector(to_unsigned(115,8) ,
18866	 => std_logic_vector(to_unsigned(130,8) ,
18867	 => std_logic_vector(to_unsigned(118,8) ,
18868	 => std_logic_vector(to_unsigned(105,8) ,
18869	 => std_logic_vector(to_unsigned(93,8) ,
18870	 => std_logic_vector(to_unsigned(90,8) ,
18871	 => std_logic_vector(to_unsigned(87,8) ,
18872	 => std_logic_vector(to_unsigned(86,8) ,
18873	 => std_logic_vector(to_unsigned(85,8) ,
18874	 => std_logic_vector(to_unsigned(91,8) ,
18875	 => std_logic_vector(to_unsigned(90,8) ,
18876	 => std_logic_vector(to_unsigned(91,8) ,
18877	 => std_logic_vector(to_unsigned(91,8) ,
18878	 => std_logic_vector(to_unsigned(87,8) ,
18879	 => std_logic_vector(to_unsigned(81,8) ,
18880	 => std_logic_vector(to_unsigned(81,8) ,
18881	 => std_logic_vector(to_unsigned(152,8) ,
18882	 => std_logic_vector(to_unsigned(156,8) ,
18883	 => std_logic_vector(to_unsigned(154,8) ,
18884	 => std_logic_vector(to_unsigned(151,8) ,
18885	 => std_logic_vector(to_unsigned(149,8) ,
18886	 => std_logic_vector(to_unsigned(156,8) ,
18887	 => std_logic_vector(to_unsigned(154,8) ,
18888	 => std_logic_vector(to_unsigned(154,8) ,
18889	 => std_logic_vector(to_unsigned(152,8) ,
18890	 => std_logic_vector(to_unsigned(152,8) ,
18891	 => std_logic_vector(to_unsigned(154,8) ,
18892	 => std_logic_vector(to_unsigned(156,8) ,
18893	 => std_logic_vector(to_unsigned(157,8) ,
18894	 => std_logic_vector(to_unsigned(173,8) ,
18895	 => std_logic_vector(to_unsigned(144,8) ,
18896	 => std_logic_vector(to_unsigned(56,8) ,
18897	 => std_logic_vector(to_unsigned(11,8) ,
18898	 => std_logic_vector(to_unsigned(3,8) ,
18899	 => std_logic_vector(to_unsigned(3,8) ,
18900	 => std_logic_vector(to_unsigned(3,8) ,
18901	 => std_logic_vector(to_unsigned(3,8) ,
18902	 => std_logic_vector(to_unsigned(41,8) ,
18903	 => std_logic_vector(to_unsigned(157,8) ,
18904	 => std_logic_vector(to_unsigned(146,8) ,
18905	 => std_logic_vector(to_unsigned(91,8) ,
18906	 => std_logic_vector(to_unsigned(13,8) ,
18907	 => std_logic_vector(to_unsigned(1,8) ,
18908	 => std_logic_vector(to_unsigned(4,8) ,
18909	 => std_logic_vector(to_unsigned(4,8) ,
18910	 => std_logic_vector(to_unsigned(6,8) ,
18911	 => std_logic_vector(to_unsigned(7,8) ,
18912	 => std_logic_vector(to_unsigned(13,8) ,
18913	 => std_logic_vector(to_unsigned(10,8) ,
18914	 => std_logic_vector(to_unsigned(4,8) ,
18915	 => std_logic_vector(to_unsigned(2,8) ,
18916	 => std_logic_vector(to_unsigned(6,8) ,
18917	 => std_logic_vector(to_unsigned(100,8) ,
18918	 => std_logic_vector(to_unsigned(183,8) ,
18919	 => std_logic_vector(to_unsigned(156,8) ,
18920	 => std_logic_vector(to_unsigned(164,8) ,
18921	 => std_logic_vector(to_unsigned(159,8) ,
18922	 => std_logic_vector(to_unsigned(157,8) ,
18923	 => std_logic_vector(to_unsigned(159,8) ,
18924	 => std_logic_vector(to_unsigned(163,8) ,
18925	 => std_logic_vector(to_unsigned(159,8) ,
18926	 => std_logic_vector(to_unsigned(156,8) ,
18927	 => std_logic_vector(to_unsigned(157,8) ,
18928	 => std_logic_vector(to_unsigned(163,8) ,
18929	 => std_logic_vector(to_unsigned(157,8) ,
18930	 => std_logic_vector(to_unsigned(154,8) ,
18931	 => std_logic_vector(to_unsigned(152,8) ,
18932	 => std_logic_vector(to_unsigned(147,8) ,
18933	 => std_logic_vector(to_unsigned(161,8) ,
18934	 => std_logic_vector(to_unsigned(142,8) ,
18935	 => std_logic_vector(to_unsigned(50,8) ,
18936	 => std_logic_vector(to_unsigned(26,8) ,
18937	 => std_logic_vector(to_unsigned(31,8) ,
18938	 => std_logic_vector(to_unsigned(76,8) ,
18939	 => std_logic_vector(to_unsigned(74,8) ,
18940	 => std_logic_vector(to_unsigned(52,8) ,
18941	 => std_logic_vector(to_unsigned(37,8) ,
18942	 => std_logic_vector(to_unsigned(35,8) ,
18943	 => std_logic_vector(to_unsigned(32,8) ,
18944	 => std_logic_vector(to_unsigned(40,8) ,
18945	 => std_logic_vector(to_unsigned(48,8) ,
18946	 => std_logic_vector(to_unsigned(15,8) ,
18947	 => std_logic_vector(to_unsigned(15,8) ,
18948	 => std_logic_vector(to_unsigned(41,8) ,
18949	 => std_logic_vector(to_unsigned(127,8) ,
18950	 => std_logic_vector(to_unsigned(173,8) ,
18951	 => std_logic_vector(to_unsigned(171,8) ,
18952	 => std_logic_vector(to_unsigned(171,8) ,
18953	 => std_logic_vector(to_unsigned(164,8) ,
18954	 => std_logic_vector(to_unsigned(163,8) ,
18955	 => std_logic_vector(to_unsigned(164,8) ,
18956	 => std_logic_vector(to_unsigned(164,8) ,
18957	 => std_logic_vector(to_unsigned(159,8) ,
18958	 => std_logic_vector(to_unsigned(161,8) ,
18959	 => std_logic_vector(to_unsigned(161,8) ,
18960	 => std_logic_vector(to_unsigned(164,8) ,
18961	 => std_logic_vector(to_unsigned(164,8) ,
18962	 => std_logic_vector(to_unsigned(157,8) ,
18963	 => std_logic_vector(to_unsigned(163,8) ,
18964	 => std_logic_vector(to_unsigned(163,8) ,
18965	 => std_logic_vector(to_unsigned(164,8) ,
18966	 => std_logic_vector(to_unsigned(170,8) ,
18967	 => std_logic_vector(to_unsigned(142,8) ,
18968	 => std_logic_vector(to_unsigned(74,8) ,
18969	 => std_logic_vector(to_unsigned(52,8) ,
18970	 => std_logic_vector(to_unsigned(9,8) ,
18971	 => std_logic_vector(to_unsigned(1,8) ,
18972	 => std_logic_vector(to_unsigned(4,8) ,
18973	 => std_logic_vector(to_unsigned(7,8) ,
18974	 => std_logic_vector(to_unsigned(6,8) ,
18975	 => std_logic_vector(to_unsigned(3,8) ,
18976	 => std_logic_vector(to_unsigned(5,8) ,
18977	 => std_logic_vector(to_unsigned(10,8) ,
18978	 => std_logic_vector(to_unsigned(5,8) ,
18979	 => std_logic_vector(to_unsigned(2,8) ,
18980	 => std_logic_vector(to_unsigned(1,8) ,
18981	 => std_logic_vector(to_unsigned(37,8) ,
18982	 => std_logic_vector(to_unsigned(181,8) ,
18983	 => std_logic_vector(to_unsigned(170,8) ,
18984	 => std_logic_vector(to_unsigned(171,8) ,
18985	 => std_logic_vector(to_unsigned(173,8) ,
18986	 => std_logic_vector(to_unsigned(173,8) ,
18987	 => std_logic_vector(to_unsigned(173,8) ,
18988	 => std_logic_vector(to_unsigned(168,8) ,
18989	 => std_logic_vector(to_unsigned(161,8) ,
18990	 => std_logic_vector(to_unsigned(161,8) ,
18991	 => std_logic_vector(to_unsigned(161,8) ,
18992	 => std_logic_vector(to_unsigned(161,8) ,
18993	 => std_logic_vector(to_unsigned(146,8) ,
18994	 => std_logic_vector(to_unsigned(133,8) ,
18995	 => std_logic_vector(to_unsigned(164,8) ,
18996	 => std_logic_vector(to_unsigned(164,8) ,
18997	 => std_logic_vector(to_unsigned(166,8) ,
18998	 => std_logic_vector(to_unsigned(171,8) ,
18999	 => std_logic_vector(to_unsigned(168,8) ,
19000	 => std_logic_vector(to_unsigned(171,8) ,
19001	 => std_logic_vector(to_unsigned(173,8) ,
19002	 => std_logic_vector(to_unsigned(164,8) ,
19003	 => std_logic_vector(to_unsigned(164,8) ,
19004	 => std_logic_vector(to_unsigned(159,8) ,
19005	 => std_logic_vector(to_unsigned(163,8) ,
19006	 => std_logic_vector(to_unsigned(163,8) ,
19007	 => std_logic_vector(to_unsigned(154,8) ,
19008	 => std_logic_vector(to_unsigned(133,8) ,
19009	 => std_logic_vector(to_unsigned(124,8) ,
19010	 => std_logic_vector(to_unsigned(128,8) ,
19011	 => std_logic_vector(to_unsigned(107,8) ,
19012	 => std_logic_vector(to_unsigned(116,8) ,
19013	 => std_logic_vector(to_unsigned(130,8) ,
19014	 => std_logic_vector(to_unsigned(134,8) ,
19015	 => std_logic_vector(to_unsigned(127,8) ,
19016	 => std_logic_vector(to_unsigned(116,8) ,
19017	 => std_logic_vector(to_unsigned(127,8) ,
19018	 => std_logic_vector(to_unsigned(121,8) ,
19019	 => std_logic_vector(to_unsigned(122,8) ,
19020	 => std_logic_vector(to_unsigned(124,8) ,
19021	 => std_logic_vector(to_unsigned(118,8) ,
19022	 => std_logic_vector(to_unsigned(124,8) ,
19023	 => std_logic_vector(to_unsigned(133,8) ,
19024	 => std_logic_vector(to_unsigned(136,8) ,
19025	 => std_logic_vector(to_unsigned(151,8) ,
19026	 => std_logic_vector(to_unsigned(164,8) ,
19027	 => std_logic_vector(to_unsigned(156,8) ,
19028	 => std_logic_vector(to_unsigned(161,8) ,
19029	 => std_logic_vector(to_unsigned(159,8) ,
19030	 => std_logic_vector(to_unsigned(154,8) ,
19031	 => std_logic_vector(to_unsigned(157,8) ,
19032	 => std_logic_vector(to_unsigned(159,8) ,
19033	 => std_logic_vector(to_unsigned(157,8) ,
19034	 => std_logic_vector(to_unsigned(156,8) ,
19035	 => std_logic_vector(to_unsigned(151,8) ,
19036	 => std_logic_vector(to_unsigned(112,8) ,
19037	 => std_logic_vector(to_unsigned(92,8) ,
19038	 => std_logic_vector(to_unsigned(87,8) ,
19039	 => std_logic_vector(to_unsigned(97,8) ,
19040	 => std_logic_vector(to_unsigned(92,8) ,
19041	 => std_logic_vector(to_unsigned(85,8) ,
19042	 => std_logic_vector(to_unsigned(91,8) ,
19043	 => std_logic_vector(to_unsigned(15,8) ,
19044	 => std_logic_vector(to_unsigned(11,8) ,
19045	 => std_logic_vector(to_unsigned(59,8) ,
19046	 => std_logic_vector(to_unsigned(48,8) ,
19047	 => std_logic_vector(to_unsigned(27,8) ,
19048	 => std_logic_vector(to_unsigned(47,8) ,
19049	 => std_logic_vector(to_unsigned(64,8) ,
19050	 => std_logic_vector(to_unsigned(45,8) ,
19051	 => std_logic_vector(to_unsigned(17,8) ,
19052	 => std_logic_vector(to_unsigned(18,8) ,
19053	 => std_logic_vector(to_unsigned(63,8) ,
19054	 => std_logic_vector(to_unsigned(119,8) ,
19055	 => std_logic_vector(to_unsigned(87,8) ,
19056	 => std_logic_vector(to_unsigned(59,8) ,
19057	 => std_logic_vector(to_unsigned(77,8) ,
19058	 => std_logic_vector(to_unsigned(85,8) ,
19059	 => std_logic_vector(to_unsigned(96,8) ,
19060	 => std_logic_vector(to_unsigned(112,8) ,
19061	 => std_logic_vector(to_unsigned(147,8) ,
19062	 => std_logic_vector(to_unsigned(139,8) ,
19063	 => std_logic_vector(to_unsigned(133,8) ,
19064	 => std_logic_vector(to_unsigned(125,8) ,
19065	 => std_logic_vector(to_unsigned(103,8) ,
19066	 => std_logic_vector(to_unsigned(95,8) ,
19067	 => std_logic_vector(to_unsigned(81,8) ,
19068	 => std_logic_vector(to_unsigned(70,8) ,
19069	 => std_logic_vector(to_unsigned(61,8) ,
19070	 => std_logic_vector(to_unsigned(65,8) ,
19071	 => std_logic_vector(to_unsigned(64,8) ,
19072	 => std_logic_vector(to_unsigned(63,8) ,
19073	 => std_logic_vector(to_unsigned(57,8) ,
19074	 => std_logic_vector(to_unsigned(68,8) ,
19075	 => std_logic_vector(to_unsigned(79,8) ,
19076	 => std_logic_vector(to_unsigned(82,8) ,
19077	 => std_logic_vector(to_unsigned(73,8) ,
19078	 => std_logic_vector(to_unsigned(71,8) ,
19079	 => std_logic_vector(to_unsigned(85,8) ,
19080	 => std_logic_vector(to_unsigned(78,8) ,
19081	 => std_logic_vector(to_unsigned(73,8) ,
19082	 => std_logic_vector(to_unsigned(86,8) ,
19083	 => std_logic_vector(to_unsigned(69,8) ,
19084	 => std_logic_vector(to_unsigned(53,8) ,
19085	 => std_logic_vector(to_unsigned(62,8) ,
19086	 => std_logic_vector(to_unsigned(69,8) ,
19087	 => std_logic_vector(to_unsigned(59,8) ,
19088	 => std_logic_vector(to_unsigned(78,8) ,
19089	 => std_logic_vector(to_unsigned(77,8) ,
19090	 => std_logic_vector(to_unsigned(55,8) ,
19091	 => std_logic_vector(to_unsigned(50,8) ,
19092	 => std_logic_vector(to_unsigned(63,8) ,
19093	 => std_logic_vector(to_unsigned(78,8) ,
19094	 => std_logic_vector(to_unsigned(66,8) ,
19095	 => std_logic_vector(to_unsigned(58,8) ,
19096	 => std_logic_vector(to_unsigned(61,8) ,
19097	 => std_logic_vector(to_unsigned(59,8) ,
19098	 => std_logic_vector(to_unsigned(61,8) ,
19099	 => std_logic_vector(to_unsigned(57,8) ,
19100	 => std_logic_vector(to_unsigned(61,8) ,
19101	 => std_logic_vector(to_unsigned(64,8) ,
19102	 => std_logic_vector(to_unsigned(67,8) ,
19103	 => std_logic_vector(to_unsigned(73,8) ,
19104	 => std_logic_vector(to_unsigned(70,8) ,
19105	 => std_logic_vector(to_unsigned(81,8) ,
19106	 => std_logic_vector(to_unsigned(80,8) ,
19107	 => std_logic_vector(to_unsigned(64,8) ,
19108	 => std_logic_vector(to_unsigned(70,8) ,
19109	 => std_logic_vector(to_unsigned(74,8) ,
19110	 => std_logic_vector(to_unsigned(79,8) ,
19111	 => std_logic_vector(to_unsigned(97,8) ,
19112	 => std_logic_vector(to_unsigned(92,8) ,
19113	 => std_logic_vector(to_unsigned(87,8) ,
19114	 => std_logic_vector(to_unsigned(90,8) ,
19115	 => std_logic_vector(to_unsigned(95,8) ,
19116	 => std_logic_vector(to_unsigned(114,8) ,
19117	 => std_logic_vector(to_unsigned(122,8) ,
19118	 => std_logic_vector(to_unsigned(124,8) ,
19119	 => std_logic_vector(to_unsigned(136,8) ,
19120	 => std_logic_vector(to_unsigned(136,8) ,
19121	 => std_logic_vector(to_unsigned(139,8) ,
19122	 => std_logic_vector(to_unsigned(141,8) ,
19123	 => std_logic_vector(to_unsigned(141,8) ,
19124	 => std_logic_vector(to_unsigned(142,8) ,
19125	 => std_logic_vector(to_unsigned(138,8) ,
19126	 => std_logic_vector(to_unsigned(141,8) ,
19127	 => std_logic_vector(to_unsigned(142,8) ,
19128	 => std_logic_vector(to_unsigned(144,8) ,
19129	 => std_logic_vector(to_unsigned(149,8) ,
19130	 => std_logic_vector(to_unsigned(45,8) ,
19131	 => std_logic_vector(to_unsigned(0,8) ,
19132	 => std_logic_vector(to_unsigned(0,8) ,
19133	 => std_logic_vector(to_unsigned(28,8) ,
19134	 => std_logic_vector(to_unsigned(175,8) ,
19135	 => std_logic_vector(to_unsigned(152,8) ,
19136	 => std_logic_vector(to_unsigned(151,8) ,
19137	 => std_logic_vector(to_unsigned(152,8) ,
19138	 => std_logic_vector(to_unsigned(139,8) ,
19139	 => std_logic_vector(to_unsigned(151,8) ,
19140	 => std_logic_vector(to_unsigned(159,8) ,
19141	 => std_logic_vector(to_unsigned(125,8) ,
19142	 => std_logic_vector(to_unsigned(107,8) ,
19143	 => std_logic_vector(to_unsigned(103,8) ,
19144	 => std_logic_vector(to_unsigned(93,8) ,
19145	 => std_logic_vector(to_unsigned(93,8) ,
19146	 => std_logic_vector(to_unsigned(86,8) ,
19147	 => std_logic_vector(to_unsigned(82,8) ,
19148	 => std_logic_vector(to_unsigned(80,8) ,
19149	 => std_logic_vector(to_unsigned(79,8) ,
19150	 => std_logic_vector(to_unsigned(79,8) ,
19151	 => std_logic_vector(to_unsigned(84,8) ,
19152	 => std_logic_vector(to_unsigned(84,8) ,
19153	 => std_logic_vector(to_unsigned(73,8) ,
19154	 => std_logic_vector(to_unsigned(81,8) ,
19155	 => std_logic_vector(to_unsigned(90,8) ,
19156	 => std_logic_vector(to_unsigned(104,8) ,
19157	 => std_logic_vector(to_unsigned(80,8) ,
19158	 => std_logic_vector(to_unsigned(57,8) ,
19159	 => std_logic_vector(to_unsigned(68,8) ,
19160	 => std_logic_vector(to_unsigned(82,8) ,
19161	 => std_logic_vector(to_unsigned(96,8) ,
19162	 => std_logic_vector(to_unsigned(97,8) ,
19163	 => std_logic_vector(to_unsigned(100,8) ,
19164	 => std_logic_vector(to_unsigned(105,8) ,
19165	 => std_logic_vector(to_unsigned(97,8) ,
19166	 => std_logic_vector(to_unsigned(84,8) ,
19167	 => std_logic_vector(to_unsigned(78,8) ,
19168	 => std_logic_vector(to_unsigned(93,8) ,
19169	 => std_logic_vector(to_unsigned(97,8) ,
19170	 => std_logic_vector(to_unsigned(87,8) ,
19171	 => std_logic_vector(to_unsigned(91,8) ,
19172	 => std_logic_vector(to_unsigned(95,8) ,
19173	 => std_logic_vector(to_unsigned(91,8) ,
19174	 => std_logic_vector(to_unsigned(93,8) ,
19175	 => std_logic_vector(to_unsigned(92,8) ,
19176	 => std_logic_vector(to_unsigned(86,8) ,
19177	 => std_logic_vector(to_unsigned(101,8) ,
19178	 => std_logic_vector(to_unsigned(124,8) ,
19179	 => std_logic_vector(to_unsigned(134,8) ,
19180	 => std_logic_vector(to_unsigned(133,8) ,
19181	 => std_logic_vector(to_unsigned(151,8) ,
19182	 => std_logic_vector(to_unsigned(154,8) ,
19183	 => std_logic_vector(to_unsigned(124,8) ,
19184	 => std_logic_vector(to_unsigned(105,8) ,
19185	 => std_logic_vector(to_unsigned(131,8) ,
19186	 => std_logic_vector(to_unsigned(147,8) ,
19187	 => std_logic_vector(to_unsigned(121,8) ,
19188	 => std_logic_vector(to_unsigned(107,8) ,
19189	 => std_logic_vector(to_unsigned(99,8) ,
19190	 => std_logic_vector(to_unsigned(88,8) ,
19191	 => std_logic_vector(to_unsigned(85,8) ,
19192	 => std_logic_vector(to_unsigned(91,8) ,
19193	 => std_logic_vector(to_unsigned(91,8) ,
19194	 => std_logic_vector(to_unsigned(96,8) ,
19195	 => std_logic_vector(to_unsigned(96,8) ,
19196	 => std_logic_vector(to_unsigned(95,8) ,
19197	 => std_logic_vector(to_unsigned(93,8) ,
19198	 => std_logic_vector(to_unsigned(87,8) ,
19199	 => std_logic_vector(to_unsigned(86,8) ,
19200	 => std_logic_vector(to_unsigned(90,8) ,
19201	 => std_logic_vector(to_unsigned(156,8) ,
19202	 => std_logic_vector(to_unsigned(154,8) ,
19203	 => std_logic_vector(to_unsigned(154,8) ,
19204	 => std_logic_vector(to_unsigned(151,8) ,
19205	 => std_logic_vector(to_unsigned(146,8) ,
19206	 => std_logic_vector(to_unsigned(154,8) ,
19207	 => std_logic_vector(to_unsigned(157,8) ,
19208	 => std_logic_vector(to_unsigned(156,8) ,
19209	 => std_logic_vector(to_unsigned(156,8) ,
19210	 => std_logic_vector(to_unsigned(156,8) ,
19211	 => std_logic_vector(to_unsigned(157,8) ,
19212	 => std_logic_vector(to_unsigned(156,8) ,
19213	 => std_logic_vector(to_unsigned(173,8) ,
19214	 => std_logic_vector(to_unsigned(118,8) ,
19215	 => std_logic_vector(to_unsigned(13,8) ,
19216	 => std_logic_vector(to_unsigned(1,8) ,
19217	 => std_logic_vector(to_unsigned(2,8) ,
19218	 => std_logic_vector(to_unsigned(5,8) ,
19219	 => std_logic_vector(to_unsigned(3,8) ,
19220	 => std_logic_vector(to_unsigned(2,8) ,
19221	 => std_logic_vector(to_unsigned(1,8) ,
19222	 => std_logic_vector(to_unsigned(1,8) ,
19223	 => std_logic_vector(to_unsigned(42,8) ,
19224	 => std_logic_vector(to_unsigned(78,8) ,
19225	 => std_logic_vector(to_unsigned(6,8) ,
19226	 => std_logic_vector(to_unsigned(1,8) ,
19227	 => std_logic_vector(to_unsigned(2,8) ,
19228	 => std_logic_vector(to_unsigned(4,8) ,
19229	 => std_logic_vector(to_unsigned(7,8) ,
19230	 => std_logic_vector(to_unsigned(5,8) ,
19231	 => std_logic_vector(to_unsigned(8,8) ,
19232	 => std_logic_vector(to_unsigned(6,8) ,
19233	 => std_logic_vector(to_unsigned(2,8) ,
19234	 => std_logic_vector(to_unsigned(2,8) ,
19235	 => std_logic_vector(to_unsigned(2,8) ,
19236	 => std_logic_vector(to_unsigned(3,8) ,
19237	 => std_logic_vector(to_unsigned(70,8) ,
19238	 => std_logic_vector(to_unsigned(183,8) ,
19239	 => std_logic_vector(to_unsigned(161,8) ,
19240	 => std_logic_vector(to_unsigned(163,8) ,
19241	 => std_logic_vector(to_unsigned(157,8) ,
19242	 => std_logic_vector(to_unsigned(157,8) ,
19243	 => std_logic_vector(to_unsigned(159,8) ,
19244	 => std_logic_vector(to_unsigned(159,8) ,
19245	 => std_logic_vector(to_unsigned(164,8) ,
19246	 => std_logic_vector(to_unsigned(161,8) ,
19247	 => std_logic_vector(to_unsigned(159,8) ,
19248	 => std_logic_vector(to_unsigned(161,8) ,
19249	 => std_logic_vector(to_unsigned(154,8) ,
19250	 => std_logic_vector(to_unsigned(154,8) ,
19251	 => std_logic_vector(to_unsigned(159,8) ,
19252	 => std_logic_vector(to_unsigned(157,8) ,
19253	 => std_logic_vector(to_unsigned(156,8) ,
19254	 => std_logic_vector(to_unsigned(171,8) ,
19255	 => std_logic_vector(to_unsigned(88,8) ,
19256	 => std_logic_vector(to_unsigned(10,8) ,
19257	 => std_logic_vector(to_unsigned(21,8) ,
19258	 => std_logic_vector(to_unsigned(63,8) ,
19259	 => std_logic_vector(to_unsigned(68,8) ,
19260	 => std_logic_vector(to_unsigned(55,8) ,
19261	 => std_logic_vector(to_unsigned(32,8) ,
19262	 => std_logic_vector(to_unsigned(25,8) ,
19263	 => std_logic_vector(to_unsigned(17,8) ,
19264	 => std_logic_vector(to_unsigned(17,8) ,
19265	 => std_logic_vector(to_unsigned(19,8) ,
19266	 => std_logic_vector(to_unsigned(24,8) ,
19267	 => std_logic_vector(to_unsigned(60,8) ,
19268	 => std_logic_vector(to_unsigned(147,8) ,
19269	 => std_logic_vector(to_unsigned(177,8) ,
19270	 => std_logic_vector(to_unsigned(166,8) ,
19271	 => std_logic_vector(to_unsigned(166,8) ,
19272	 => std_logic_vector(to_unsigned(170,8) ,
19273	 => std_logic_vector(to_unsigned(170,8) ,
19274	 => std_logic_vector(to_unsigned(170,8) ,
19275	 => std_logic_vector(to_unsigned(164,8) ,
19276	 => std_logic_vector(to_unsigned(166,8) ,
19277	 => std_logic_vector(to_unsigned(164,8) ,
19278	 => std_logic_vector(to_unsigned(170,8) ,
19279	 => std_logic_vector(to_unsigned(164,8) ,
19280	 => std_logic_vector(to_unsigned(163,8) ,
19281	 => std_logic_vector(to_unsigned(163,8) ,
19282	 => std_logic_vector(to_unsigned(161,8) ,
19283	 => std_logic_vector(to_unsigned(161,8) ,
19284	 => std_logic_vector(to_unsigned(163,8) ,
19285	 => std_logic_vector(to_unsigned(161,8) ,
19286	 => std_logic_vector(to_unsigned(168,8) ,
19287	 => std_logic_vector(to_unsigned(175,8) ,
19288	 => std_logic_vector(to_unsigned(192,8) ,
19289	 => std_logic_vector(to_unsigned(204,8) ,
19290	 => std_logic_vector(to_unsigned(27,8) ,
19291	 => std_logic_vector(to_unsigned(1,8) ,
19292	 => std_logic_vector(to_unsigned(6,8) ,
19293	 => std_logic_vector(to_unsigned(10,8) ,
19294	 => std_logic_vector(to_unsigned(8,8) ,
19295	 => std_logic_vector(to_unsigned(4,8) ,
19296	 => std_logic_vector(to_unsigned(6,8) ,
19297	 => std_logic_vector(to_unsigned(6,8) ,
19298	 => std_logic_vector(to_unsigned(8,8) ,
19299	 => std_logic_vector(to_unsigned(8,8) ,
19300	 => std_logic_vector(to_unsigned(6,8) ,
19301	 => std_logic_vector(to_unsigned(107,8) ,
19302	 => std_logic_vector(to_unsigned(194,8) ,
19303	 => std_logic_vector(to_unsigned(168,8) ,
19304	 => std_logic_vector(to_unsigned(166,8) ,
19305	 => std_logic_vector(to_unsigned(171,8) ,
19306	 => std_logic_vector(to_unsigned(175,8) ,
19307	 => std_logic_vector(to_unsigned(171,8) ,
19308	 => std_logic_vector(to_unsigned(164,8) ,
19309	 => std_logic_vector(to_unsigned(166,8) ,
19310	 => std_logic_vector(to_unsigned(163,8) ,
19311	 => std_logic_vector(to_unsigned(159,8) ,
19312	 => std_logic_vector(to_unsigned(161,8) ,
19313	 => std_logic_vector(to_unsigned(141,8) ,
19314	 => std_logic_vector(to_unsigned(133,8) ,
19315	 => std_logic_vector(to_unsigned(161,8) ,
19316	 => std_logic_vector(to_unsigned(168,8) ,
19317	 => std_logic_vector(to_unsigned(168,8) ,
19318	 => std_logic_vector(to_unsigned(166,8) ,
19319	 => std_logic_vector(to_unsigned(168,8) ,
19320	 => std_logic_vector(to_unsigned(168,8) ,
19321	 => std_logic_vector(to_unsigned(166,8) ,
19322	 => std_logic_vector(to_unsigned(161,8) ,
19323	 => std_logic_vector(to_unsigned(163,8) ,
19324	 => std_logic_vector(to_unsigned(166,8) ,
19325	 => std_logic_vector(to_unsigned(164,8) ,
19326	 => std_logic_vector(to_unsigned(151,8) ,
19327	 => std_logic_vector(to_unsigned(147,8) ,
19328	 => std_logic_vector(to_unsigned(147,8) ,
19329	 => std_logic_vector(to_unsigned(125,8) ,
19330	 => std_logic_vector(to_unsigned(121,8) ,
19331	 => std_logic_vector(to_unsigned(124,8) ,
19332	 => std_logic_vector(to_unsigned(128,8) ,
19333	 => std_logic_vector(to_unsigned(125,8) ,
19334	 => std_logic_vector(to_unsigned(114,8) ,
19335	 => std_logic_vector(to_unsigned(115,8) ,
19336	 => std_logic_vector(to_unsigned(114,8) ,
19337	 => std_logic_vector(to_unsigned(127,8) ,
19338	 => std_logic_vector(to_unsigned(119,8) ,
19339	 => std_logic_vector(to_unsigned(105,8) ,
19340	 => std_logic_vector(to_unsigned(118,8) ,
19341	 => std_logic_vector(to_unsigned(119,8) ,
19342	 => std_logic_vector(to_unsigned(124,8) ,
19343	 => std_logic_vector(to_unsigned(139,8) ,
19344	 => std_logic_vector(to_unsigned(134,8) ,
19345	 => std_logic_vector(to_unsigned(139,8) ,
19346	 => std_logic_vector(to_unsigned(151,8) ,
19347	 => std_logic_vector(to_unsigned(144,8) ,
19348	 => std_logic_vector(to_unsigned(142,8) ,
19349	 => std_logic_vector(to_unsigned(151,8) ,
19350	 => std_logic_vector(to_unsigned(154,8) ,
19351	 => std_logic_vector(to_unsigned(157,8) ,
19352	 => std_logic_vector(to_unsigned(159,8) ,
19353	 => std_logic_vector(to_unsigned(154,8) ,
19354	 => std_logic_vector(to_unsigned(156,8) ,
19355	 => std_logic_vector(to_unsigned(152,8) ,
19356	 => std_logic_vector(to_unsigned(122,8) ,
19357	 => std_logic_vector(to_unsigned(99,8) ,
19358	 => std_logic_vector(to_unsigned(88,8) ,
19359	 => std_logic_vector(to_unsigned(96,8) ,
19360	 => std_logic_vector(to_unsigned(93,8) ,
19361	 => std_logic_vector(to_unsigned(109,8) ,
19362	 => std_logic_vector(to_unsigned(60,8) ,
19363	 => std_logic_vector(to_unsigned(2,8) ,
19364	 => std_logic_vector(to_unsigned(3,8) ,
19365	 => std_logic_vector(to_unsigned(8,8) ,
19366	 => std_logic_vector(to_unsigned(12,8) ,
19367	 => std_logic_vector(to_unsigned(12,8) ,
19368	 => std_logic_vector(to_unsigned(30,8) ,
19369	 => std_logic_vector(to_unsigned(72,8) ,
19370	 => std_logic_vector(to_unsigned(81,8) ,
19371	 => std_logic_vector(to_unsigned(32,8) ,
19372	 => std_logic_vector(to_unsigned(7,8) ,
19373	 => std_logic_vector(to_unsigned(20,8) ,
19374	 => std_logic_vector(to_unsigned(78,8) ,
19375	 => std_logic_vector(to_unsigned(90,8) ,
19376	 => std_logic_vector(to_unsigned(56,8) ,
19377	 => std_logic_vector(to_unsigned(51,8) ,
19378	 => std_logic_vector(to_unsigned(69,8) ,
19379	 => std_logic_vector(to_unsigned(91,8) ,
19380	 => std_logic_vector(to_unsigned(95,8) ,
19381	 => std_logic_vector(to_unsigned(134,8) ,
19382	 => std_logic_vector(to_unsigned(115,8) ,
19383	 => std_logic_vector(to_unsigned(100,8) ,
19384	 => std_logic_vector(to_unsigned(90,8) ,
19385	 => std_logic_vector(to_unsigned(80,8) ,
19386	 => std_logic_vector(to_unsigned(73,8) ,
19387	 => std_logic_vector(to_unsigned(57,8) ,
19388	 => std_logic_vector(to_unsigned(64,8) ,
19389	 => std_logic_vector(to_unsigned(64,8) ,
19390	 => std_logic_vector(to_unsigned(67,8) ,
19391	 => std_logic_vector(to_unsigned(76,8) ,
19392	 => std_logic_vector(to_unsigned(73,8) ,
19393	 => std_logic_vector(to_unsigned(67,8) ,
19394	 => std_logic_vector(to_unsigned(68,8) ,
19395	 => std_logic_vector(to_unsigned(70,8) ,
19396	 => std_logic_vector(to_unsigned(81,8) ,
19397	 => std_logic_vector(to_unsigned(72,8) ,
19398	 => std_logic_vector(to_unsigned(81,8) ,
19399	 => std_logic_vector(to_unsigned(105,8) ,
19400	 => std_logic_vector(to_unsigned(114,8) ,
19401	 => std_logic_vector(to_unsigned(97,8) ,
19402	 => std_logic_vector(to_unsigned(90,8) ,
19403	 => std_logic_vector(to_unsigned(77,8) ,
19404	 => std_logic_vector(to_unsigned(60,8) ,
19405	 => std_logic_vector(to_unsigned(62,8) ,
19406	 => std_logic_vector(to_unsigned(61,8) ,
19407	 => std_logic_vector(to_unsigned(54,8) ,
19408	 => std_logic_vector(to_unsigned(65,8) ,
19409	 => std_logic_vector(to_unsigned(66,8) ,
19410	 => std_logic_vector(to_unsigned(67,8) ,
19411	 => std_logic_vector(to_unsigned(70,8) ,
19412	 => std_logic_vector(to_unsigned(67,8) ,
19413	 => std_logic_vector(to_unsigned(55,8) ,
19414	 => std_logic_vector(to_unsigned(59,8) ,
19415	 => std_logic_vector(to_unsigned(61,8) ,
19416	 => std_logic_vector(to_unsigned(61,8) ,
19417	 => std_logic_vector(to_unsigned(59,8) ,
19418	 => std_logic_vector(to_unsigned(56,8) ,
19419	 => std_logic_vector(to_unsigned(52,8) ,
19420	 => std_logic_vector(to_unsigned(51,8) ,
19421	 => std_logic_vector(to_unsigned(62,8) ,
19422	 => std_logic_vector(to_unsigned(73,8) ,
19423	 => std_logic_vector(to_unsigned(77,8) ,
19424	 => std_logic_vector(to_unsigned(87,8) ,
19425	 => std_logic_vector(to_unsigned(97,8) ,
19426	 => std_logic_vector(to_unsigned(76,8) ,
19427	 => std_logic_vector(to_unsigned(67,8) ,
19428	 => std_logic_vector(to_unsigned(80,8) ,
19429	 => std_logic_vector(to_unsigned(84,8) ,
19430	 => std_logic_vector(to_unsigned(81,8) ,
19431	 => std_logic_vector(to_unsigned(85,8) ,
19432	 => std_logic_vector(to_unsigned(86,8) ,
19433	 => std_logic_vector(to_unsigned(95,8) ,
19434	 => std_logic_vector(to_unsigned(92,8) ,
19435	 => std_logic_vector(to_unsigned(86,8) ,
19436	 => std_logic_vector(to_unsigned(111,8) ,
19437	 => std_logic_vector(to_unsigned(142,8) ,
19438	 => std_logic_vector(to_unsigned(142,8) ,
19439	 => std_logic_vector(to_unsigned(142,8) ,
19440	 => std_logic_vector(to_unsigned(144,8) ,
19441	 => std_logic_vector(to_unsigned(141,8) ,
19442	 => std_logic_vector(to_unsigned(146,8) ,
19443	 => std_logic_vector(to_unsigned(144,8) ,
19444	 => std_logic_vector(to_unsigned(139,8) ,
19445	 => std_logic_vector(to_unsigned(147,8) ,
19446	 => std_logic_vector(to_unsigned(127,8) ,
19447	 => std_logic_vector(to_unsigned(109,8) ,
19448	 => std_logic_vector(to_unsigned(107,8) ,
19449	 => std_logic_vector(to_unsigned(97,8) ,
19450	 => std_logic_vector(to_unsigned(40,8) ,
19451	 => std_logic_vector(to_unsigned(1,8) ,
19452	 => std_logic_vector(to_unsigned(0,8) ,
19453	 => std_logic_vector(to_unsigned(10,8) ,
19454	 => std_logic_vector(to_unsigned(146,8) ,
19455	 => std_logic_vector(to_unsigned(164,8) ,
19456	 => std_logic_vector(to_unsigned(154,8) ,
19457	 => std_logic_vector(to_unsigned(157,8) ,
19458	 => std_logic_vector(to_unsigned(121,8) ,
19459	 => std_logic_vector(to_unsigned(131,8) ,
19460	 => std_logic_vector(to_unsigned(164,8) ,
19461	 => std_logic_vector(to_unsigned(146,8) ,
19462	 => std_logic_vector(to_unsigned(118,8) ,
19463	 => std_logic_vector(to_unsigned(101,8) ,
19464	 => std_logic_vector(to_unsigned(103,8) ,
19465	 => std_logic_vector(to_unsigned(116,8) ,
19466	 => std_logic_vector(to_unsigned(91,8) ,
19467	 => std_logic_vector(to_unsigned(79,8) ,
19468	 => std_logic_vector(to_unsigned(90,8) ,
19469	 => std_logic_vector(to_unsigned(81,8) ,
19470	 => std_logic_vector(to_unsigned(73,8) ,
19471	 => std_logic_vector(to_unsigned(85,8) ,
19472	 => std_logic_vector(to_unsigned(95,8) ,
19473	 => std_logic_vector(to_unsigned(82,8) ,
19474	 => std_logic_vector(to_unsigned(80,8) ,
19475	 => std_logic_vector(to_unsigned(78,8) ,
19476	 => std_logic_vector(to_unsigned(76,8) ,
19477	 => std_logic_vector(to_unsigned(37,8) ,
19478	 => std_logic_vector(to_unsigned(8,8) ,
19479	 => std_logic_vector(to_unsigned(7,8) ,
19480	 => std_logic_vector(to_unsigned(10,8) ,
19481	 => std_logic_vector(to_unsigned(18,8) ,
19482	 => std_logic_vector(to_unsigned(22,8) ,
19483	 => std_logic_vector(to_unsigned(20,8) ,
19484	 => std_logic_vector(to_unsigned(29,8) ,
19485	 => std_logic_vector(to_unsigned(79,8) ,
19486	 => std_logic_vector(to_unsigned(122,8) ,
19487	 => std_logic_vector(to_unsigned(101,8) ,
19488	 => std_logic_vector(to_unsigned(96,8) ,
19489	 => std_logic_vector(to_unsigned(95,8) ,
19490	 => std_logic_vector(to_unsigned(90,8) ,
19491	 => std_logic_vector(to_unsigned(97,8) ,
19492	 => std_logic_vector(to_unsigned(105,8) ,
19493	 => std_logic_vector(to_unsigned(101,8) ,
19494	 => std_logic_vector(to_unsigned(100,8) ,
19495	 => std_logic_vector(to_unsigned(105,8) ,
19496	 => std_logic_vector(to_unsigned(97,8) ,
19497	 => std_logic_vector(to_unsigned(97,8) ,
19498	 => std_logic_vector(to_unsigned(115,8) ,
19499	 => std_logic_vector(to_unsigned(146,8) ,
19500	 => std_logic_vector(to_unsigned(157,8) ,
19501	 => std_logic_vector(to_unsigned(151,8) ,
19502	 => std_logic_vector(to_unsigned(138,8) ,
19503	 => std_logic_vector(to_unsigned(115,8) ,
19504	 => std_logic_vector(to_unsigned(100,8) ,
19505	 => std_logic_vector(to_unsigned(107,8) ,
19506	 => std_logic_vector(to_unsigned(105,8) ,
19507	 => std_logic_vector(to_unsigned(95,8) ,
19508	 => std_logic_vector(to_unsigned(97,8) ,
19509	 => std_logic_vector(to_unsigned(109,8) ,
19510	 => std_logic_vector(to_unsigned(103,8) ,
19511	 => std_logic_vector(to_unsigned(92,8) ,
19512	 => std_logic_vector(to_unsigned(96,8) ,
19513	 => std_logic_vector(to_unsigned(95,8) ,
19514	 => std_logic_vector(to_unsigned(91,8) ,
19515	 => std_logic_vector(to_unsigned(92,8) ,
19516	 => std_logic_vector(to_unsigned(95,8) ,
19517	 => std_logic_vector(to_unsigned(96,8) ,
19518	 => std_logic_vector(to_unsigned(88,8) ,
19519	 => std_logic_vector(to_unsigned(85,8) ,
19520	 => std_logic_vector(to_unsigned(88,8) ,
19521	 => std_logic_vector(to_unsigned(154,8) ,
19522	 => std_logic_vector(to_unsigned(149,8) ,
19523	 => std_logic_vector(to_unsigned(146,8) ,
19524	 => std_logic_vector(to_unsigned(146,8) ,
19525	 => std_logic_vector(to_unsigned(144,8) ,
19526	 => std_logic_vector(to_unsigned(151,8) ,
19527	 => std_logic_vector(to_unsigned(157,8) ,
19528	 => std_logic_vector(to_unsigned(159,8) ,
19529	 => std_logic_vector(to_unsigned(157,8) ,
19530	 => std_logic_vector(to_unsigned(157,8) ,
19531	 => std_logic_vector(to_unsigned(159,8) ,
19532	 => std_logic_vector(to_unsigned(159,8) ,
19533	 => std_logic_vector(to_unsigned(175,8) ,
19534	 => std_logic_vector(to_unsigned(29,8) ,
19535	 => std_logic_vector(to_unsigned(0,8) ,
19536	 => std_logic_vector(to_unsigned(3,8) ,
19537	 => std_logic_vector(to_unsigned(5,8) ,
19538	 => std_logic_vector(to_unsigned(5,8) ,
19539	 => std_logic_vector(to_unsigned(4,8) ,
19540	 => std_logic_vector(to_unsigned(2,8) ,
19541	 => std_logic_vector(to_unsigned(4,8) ,
19542	 => std_logic_vector(to_unsigned(2,8) ,
19543	 => std_logic_vector(to_unsigned(9,8) ,
19544	 => std_logic_vector(to_unsigned(27,8) ,
19545	 => std_logic_vector(to_unsigned(2,8) ,
19546	 => std_logic_vector(to_unsigned(1,8) ,
19547	 => std_logic_vector(to_unsigned(1,8) ,
19548	 => std_logic_vector(to_unsigned(4,8) ,
19549	 => std_logic_vector(to_unsigned(7,8) ,
19550	 => std_logic_vector(to_unsigned(3,8) ,
19551	 => std_logic_vector(to_unsigned(2,8) ,
19552	 => std_logic_vector(to_unsigned(1,8) ,
19553	 => std_logic_vector(to_unsigned(1,8) ,
19554	 => std_logic_vector(to_unsigned(1,8) ,
19555	 => std_logic_vector(to_unsigned(2,8) ,
19556	 => std_logic_vector(to_unsigned(4,8) ,
19557	 => std_logic_vector(to_unsigned(63,8) ,
19558	 => std_logic_vector(to_unsigned(179,8) ,
19559	 => std_logic_vector(to_unsigned(159,8) ,
19560	 => std_logic_vector(to_unsigned(157,8) ,
19561	 => std_logic_vector(to_unsigned(157,8) ,
19562	 => std_logic_vector(to_unsigned(156,8) ,
19563	 => std_logic_vector(to_unsigned(154,8) ,
19564	 => std_logic_vector(to_unsigned(161,8) ,
19565	 => std_logic_vector(to_unsigned(163,8) ,
19566	 => std_logic_vector(to_unsigned(159,8) ,
19567	 => std_logic_vector(to_unsigned(156,8) ,
19568	 => std_logic_vector(to_unsigned(159,8) ,
19569	 => std_logic_vector(to_unsigned(156,8) ,
19570	 => std_logic_vector(to_unsigned(159,8) ,
19571	 => std_logic_vector(to_unsigned(163,8) ,
19572	 => std_logic_vector(to_unsigned(166,8) ,
19573	 => std_logic_vector(to_unsigned(163,8) ,
19574	 => std_logic_vector(to_unsigned(156,8) ,
19575	 => std_logic_vector(to_unsigned(181,8) ,
19576	 => std_logic_vector(to_unsigned(47,8) ,
19577	 => std_logic_vector(to_unsigned(2,8) ,
19578	 => std_logic_vector(to_unsigned(5,8) ,
19579	 => std_logic_vector(to_unsigned(11,8) ,
19580	 => std_logic_vector(to_unsigned(9,8) ,
19581	 => std_logic_vector(to_unsigned(7,8) ,
19582	 => std_logic_vector(to_unsigned(18,8) ,
19583	 => std_logic_vector(to_unsigned(27,8) ,
19584	 => std_logic_vector(to_unsigned(24,8) ,
19585	 => std_logic_vector(to_unsigned(22,8) ,
19586	 => std_logic_vector(to_unsigned(9,8) ,
19587	 => std_logic_vector(to_unsigned(46,8) ,
19588	 => std_logic_vector(to_unsigned(134,8) ,
19589	 => std_logic_vector(to_unsigned(130,8) ,
19590	 => std_logic_vector(to_unsigned(173,8) ,
19591	 => std_logic_vector(to_unsigned(171,8) ,
19592	 => std_logic_vector(to_unsigned(168,8) ,
19593	 => std_logic_vector(to_unsigned(168,8) ,
19594	 => std_logic_vector(to_unsigned(170,8) ,
19595	 => std_logic_vector(to_unsigned(164,8) ,
19596	 => std_logic_vector(to_unsigned(168,8) ,
19597	 => std_logic_vector(to_unsigned(166,8) ,
19598	 => std_logic_vector(to_unsigned(166,8) ,
19599	 => std_logic_vector(to_unsigned(168,8) ,
19600	 => std_logic_vector(to_unsigned(164,8) ,
19601	 => std_logic_vector(to_unsigned(163,8) ,
19602	 => std_logic_vector(to_unsigned(164,8) ,
19603	 => std_logic_vector(to_unsigned(166,8) ,
19604	 => std_logic_vector(to_unsigned(164,8) ,
19605	 => std_logic_vector(to_unsigned(163,8) ,
19606	 => std_logic_vector(to_unsigned(168,8) ,
19607	 => std_logic_vector(to_unsigned(154,8) ,
19608	 => std_logic_vector(to_unsigned(163,8) ,
19609	 => std_logic_vector(to_unsigned(108,8) ,
19610	 => std_logic_vector(to_unsigned(7,8) ,
19611	 => std_logic_vector(to_unsigned(1,8) ,
19612	 => std_logic_vector(to_unsigned(5,8) ,
19613	 => std_logic_vector(to_unsigned(12,8) ,
19614	 => std_logic_vector(to_unsigned(9,8) ,
19615	 => std_logic_vector(to_unsigned(8,8) ,
19616	 => std_logic_vector(to_unsigned(9,8) ,
19617	 => std_logic_vector(to_unsigned(15,8) ,
19618	 => std_logic_vector(to_unsigned(16,8) ,
19619	 => std_logic_vector(to_unsigned(5,8) ,
19620	 => std_logic_vector(to_unsigned(5,8) ,
19621	 => std_logic_vector(to_unsigned(76,8) ,
19622	 => std_logic_vector(to_unsigned(202,8) ,
19623	 => std_logic_vector(to_unsigned(166,8) ,
19624	 => std_logic_vector(to_unsigned(166,8) ,
19625	 => std_logic_vector(to_unsigned(170,8) ,
19626	 => std_logic_vector(to_unsigned(170,8) ,
19627	 => std_logic_vector(to_unsigned(170,8) ,
19628	 => std_logic_vector(to_unsigned(168,8) ,
19629	 => std_logic_vector(to_unsigned(171,8) ,
19630	 => std_logic_vector(to_unsigned(166,8) ,
19631	 => std_logic_vector(to_unsigned(157,8) ,
19632	 => std_logic_vector(to_unsigned(157,8) ,
19633	 => std_logic_vector(to_unsigned(141,8) ,
19634	 => std_logic_vector(to_unsigned(144,8) ,
19635	 => std_logic_vector(to_unsigned(166,8) ,
19636	 => std_logic_vector(to_unsigned(168,8) ,
19637	 => std_logic_vector(to_unsigned(168,8) ,
19638	 => std_logic_vector(to_unsigned(163,8) ,
19639	 => std_logic_vector(to_unsigned(170,8) ,
19640	 => std_logic_vector(to_unsigned(164,8) ,
19641	 => std_logic_vector(to_unsigned(164,8) ,
19642	 => std_logic_vector(to_unsigned(163,8) ,
19643	 => std_logic_vector(to_unsigned(164,8) ,
19644	 => std_logic_vector(to_unsigned(164,8) ,
19645	 => std_logic_vector(to_unsigned(157,8) ,
19646	 => std_logic_vector(to_unsigned(152,8) ,
19647	 => std_logic_vector(to_unsigned(154,8) ,
19648	 => std_logic_vector(to_unsigned(151,8) ,
19649	 => std_logic_vector(to_unsigned(125,8) ,
19650	 => std_logic_vector(to_unsigned(114,8) ,
19651	 => std_logic_vector(to_unsigned(121,8) ,
19652	 => std_logic_vector(to_unsigned(124,8) ,
19653	 => std_logic_vector(to_unsigned(124,8) ,
19654	 => std_logic_vector(to_unsigned(125,8) ,
19655	 => std_logic_vector(to_unsigned(125,8) ,
19656	 => std_logic_vector(to_unsigned(128,8) ,
19657	 => std_logic_vector(to_unsigned(130,8) ,
19658	 => std_logic_vector(to_unsigned(130,8) ,
19659	 => std_logic_vector(to_unsigned(107,8) ,
19660	 => std_logic_vector(to_unsigned(104,8) ,
19661	 => std_logic_vector(to_unsigned(116,8) ,
19662	 => std_logic_vector(to_unsigned(124,8) ,
19663	 => std_logic_vector(to_unsigned(138,8) ,
19664	 => std_logic_vector(to_unsigned(128,8) ,
19665	 => std_logic_vector(to_unsigned(105,8) ,
19666	 => std_logic_vector(to_unsigned(109,8) ,
19667	 => std_logic_vector(to_unsigned(122,8) ,
19668	 => std_logic_vector(to_unsigned(122,8) ,
19669	 => std_logic_vector(to_unsigned(133,8) ,
19670	 => std_logic_vector(to_unsigned(146,8) ,
19671	 => std_logic_vector(to_unsigned(144,8) ,
19672	 => std_logic_vector(to_unsigned(151,8) ,
19673	 => std_logic_vector(to_unsigned(157,8) ,
19674	 => std_logic_vector(to_unsigned(154,8) ,
19675	 => std_logic_vector(to_unsigned(152,8) ,
19676	 => std_logic_vector(to_unsigned(149,8) ,
19677	 => std_logic_vector(to_unsigned(127,8) ,
19678	 => std_logic_vector(to_unsigned(96,8) ,
19679	 => std_logic_vector(to_unsigned(91,8) ,
19680	 => std_logic_vector(to_unsigned(104,8) ,
19681	 => std_logic_vector(to_unsigned(62,8) ,
19682	 => std_logic_vector(to_unsigned(8,8) ,
19683	 => std_logic_vector(to_unsigned(3,8) ,
19684	 => std_logic_vector(to_unsigned(16,8) ,
19685	 => std_logic_vector(to_unsigned(23,8) ,
19686	 => std_logic_vector(to_unsigned(20,8) ,
19687	 => std_logic_vector(to_unsigned(8,8) ,
19688	 => std_logic_vector(to_unsigned(7,8) ,
19689	 => std_logic_vector(to_unsigned(37,8) ,
19690	 => std_logic_vector(to_unsigned(44,8) ,
19691	 => std_logic_vector(to_unsigned(25,8) ,
19692	 => std_logic_vector(to_unsigned(4,8) ,
19693	 => std_logic_vector(to_unsigned(4,8) ,
19694	 => std_logic_vector(to_unsigned(25,8) ,
19695	 => std_logic_vector(to_unsigned(52,8) ,
19696	 => std_logic_vector(to_unsigned(35,8) ,
19697	 => std_logic_vector(to_unsigned(52,8) ,
19698	 => std_logic_vector(to_unsigned(62,8) ,
19699	 => std_logic_vector(to_unsigned(103,8) ,
19700	 => std_logic_vector(to_unsigned(147,8) ,
19701	 => std_logic_vector(to_unsigned(144,8) ,
19702	 => std_logic_vector(to_unsigned(101,8) ,
19703	 => std_logic_vector(to_unsigned(79,8) ,
19704	 => std_logic_vector(to_unsigned(74,8) ,
19705	 => std_logic_vector(to_unsigned(74,8) ,
19706	 => std_logic_vector(to_unsigned(71,8) ,
19707	 => std_logic_vector(to_unsigned(65,8) ,
19708	 => std_logic_vector(to_unsigned(59,8) ,
19709	 => std_logic_vector(to_unsigned(65,8) ,
19710	 => std_logic_vector(to_unsigned(69,8) ,
19711	 => std_logic_vector(to_unsigned(73,8) ,
19712	 => std_logic_vector(to_unsigned(71,8) ,
19713	 => std_logic_vector(to_unsigned(65,8) ,
19714	 => std_logic_vector(to_unsigned(73,8) ,
19715	 => std_logic_vector(to_unsigned(78,8) ,
19716	 => std_logic_vector(to_unsigned(73,8) ,
19717	 => std_logic_vector(to_unsigned(71,8) ,
19718	 => std_logic_vector(to_unsigned(96,8) ,
19719	 => std_logic_vector(to_unsigned(104,8) ,
19720	 => std_logic_vector(to_unsigned(99,8) ,
19721	 => std_logic_vector(to_unsigned(77,8) ,
19722	 => std_logic_vector(to_unsigned(80,8) ,
19723	 => std_logic_vector(to_unsigned(86,8) ,
19724	 => std_logic_vector(to_unsigned(61,8) ,
19725	 => std_logic_vector(to_unsigned(61,8) ,
19726	 => std_logic_vector(to_unsigned(68,8) ,
19727	 => std_logic_vector(to_unsigned(63,8) ,
19728	 => std_logic_vector(to_unsigned(64,8) ,
19729	 => std_logic_vector(to_unsigned(62,8) ,
19730	 => std_logic_vector(to_unsigned(62,8) ,
19731	 => std_logic_vector(to_unsigned(65,8) ,
19732	 => std_logic_vector(to_unsigned(60,8) ,
19733	 => std_logic_vector(to_unsigned(51,8) ,
19734	 => std_logic_vector(to_unsigned(56,8) ,
19735	 => std_logic_vector(to_unsigned(58,8) ,
19736	 => std_logic_vector(to_unsigned(56,8) ,
19737	 => std_logic_vector(to_unsigned(61,8) ,
19738	 => std_logic_vector(to_unsigned(59,8) ,
19739	 => std_logic_vector(to_unsigned(64,8) ,
19740	 => std_logic_vector(to_unsigned(63,8) ,
19741	 => std_logic_vector(to_unsigned(70,8) ,
19742	 => std_logic_vector(to_unsigned(71,8) ,
19743	 => std_logic_vector(to_unsigned(79,8) ,
19744	 => std_logic_vector(to_unsigned(73,8) ,
19745	 => std_logic_vector(to_unsigned(35,8) ,
19746	 => std_logic_vector(to_unsigned(35,8) ,
19747	 => std_logic_vector(to_unsigned(55,8) ,
19748	 => std_logic_vector(to_unsigned(71,8) ,
19749	 => std_logic_vector(to_unsigned(87,8) ,
19750	 => std_logic_vector(to_unsigned(107,8) ,
19751	 => std_logic_vector(to_unsigned(100,8) ,
19752	 => std_logic_vector(to_unsigned(96,8) ,
19753	 => std_logic_vector(to_unsigned(97,8) ,
19754	 => std_logic_vector(to_unsigned(92,8) ,
19755	 => std_logic_vector(to_unsigned(87,8) ,
19756	 => std_logic_vector(to_unsigned(104,8) ,
19757	 => std_logic_vector(to_unsigned(136,8) ,
19758	 => std_logic_vector(to_unsigned(138,8) ,
19759	 => std_logic_vector(to_unsigned(141,8) ,
19760	 => std_logic_vector(to_unsigned(146,8) ,
19761	 => std_logic_vector(to_unsigned(139,8) ,
19762	 => std_logic_vector(to_unsigned(142,8) ,
19763	 => std_logic_vector(to_unsigned(144,8) ,
19764	 => std_logic_vector(to_unsigned(146,8) ,
19765	 => std_logic_vector(to_unsigned(121,8) ,
19766	 => std_logic_vector(to_unsigned(79,8) ,
19767	 => std_logic_vector(to_unsigned(67,8) ,
19768	 => std_logic_vector(to_unsigned(64,8) ,
19769	 => std_logic_vector(to_unsigned(66,8) ,
19770	 => std_logic_vector(to_unsigned(51,8) ,
19771	 => std_logic_vector(to_unsigned(5,8) ,
19772	 => std_logic_vector(to_unsigned(0,8) ,
19773	 => std_logic_vector(to_unsigned(2,8) ,
19774	 => std_logic_vector(to_unsigned(82,8) ,
19775	 => std_logic_vector(to_unsigned(179,8) ,
19776	 => std_logic_vector(to_unsigned(157,8) ,
19777	 => std_logic_vector(to_unsigned(147,8) ,
19778	 => std_logic_vector(to_unsigned(130,8) ,
19779	 => std_logic_vector(to_unsigned(127,8) ,
19780	 => std_logic_vector(to_unsigned(136,8) ,
19781	 => std_logic_vector(to_unsigned(130,8) ,
19782	 => std_logic_vector(to_unsigned(116,8) ,
19783	 => std_logic_vector(to_unsigned(100,8) ,
19784	 => std_logic_vector(to_unsigned(118,8) ,
19785	 => std_logic_vector(to_unsigned(138,8) ,
19786	 => std_logic_vector(to_unsigned(103,8) ,
19787	 => std_logic_vector(to_unsigned(87,8) ,
19788	 => std_logic_vector(to_unsigned(103,8) ,
19789	 => std_logic_vector(to_unsigned(92,8) ,
19790	 => std_logic_vector(to_unsigned(80,8) ,
19791	 => std_logic_vector(to_unsigned(82,8) ,
19792	 => std_logic_vector(to_unsigned(84,8) ,
19793	 => std_logic_vector(to_unsigned(71,8) ,
19794	 => std_logic_vector(to_unsigned(87,8) ,
19795	 => std_logic_vector(to_unsigned(77,8) ,
19796	 => std_logic_vector(to_unsigned(25,8) ,
19797	 => std_logic_vector(to_unsigned(2,8) ,
19798	 => std_logic_vector(to_unsigned(0,8) ,
19799	 => std_logic_vector(to_unsigned(1,8) ,
19800	 => std_logic_vector(to_unsigned(0,8) ,
19801	 => std_logic_vector(to_unsigned(0,8) ,
19802	 => std_logic_vector(to_unsigned(0,8) ,
19803	 => std_logic_vector(to_unsigned(1,8) ,
19804	 => std_logic_vector(to_unsigned(2,8) ,
19805	 => std_logic_vector(to_unsigned(9,8) ,
19806	 => std_logic_vector(to_unsigned(61,8) ,
19807	 => std_logic_vector(to_unsigned(118,8) ,
19808	 => std_logic_vector(to_unsigned(96,8) ,
19809	 => std_logic_vector(to_unsigned(92,8) ,
19810	 => std_logic_vector(to_unsigned(99,8) ,
19811	 => std_logic_vector(to_unsigned(95,8) ,
19812	 => std_logic_vector(to_unsigned(105,8) ,
19813	 => std_logic_vector(to_unsigned(100,8) ,
19814	 => std_logic_vector(to_unsigned(101,8) ,
19815	 => std_logic_vector(to_unsigned(118,8) ,
19816	 => std_logic_vector(to_unsigned(118,8) ,
19817	 => std_logic_vector(to_unsigned(124,8) ,
19818	 => std_logic_vector(to_unsigned(136,8) ,
19819	 => std_logic_vector(to_unsigned(138,8) ,
19820	 => std_logic_vector(to_unsigned(136,8) ,
19821	 => std_logic_vector(to_unsigned(133,8) ,
19822	 => std_logic_vector(to_unsigned(130,8) ,
19823	 => std_logic_vector(to_unsigned(111,8) ,
19824	 => std_logic_vector(to_unsigned(100,8) ,
19825	 => std_logic_vector(to_unsigned(100,8) ,
19826	 => std_logic_vector(to_unsigned(101,8) ,
19827	 => std_logic_vector(to_unsigned(99,8) ,
19828	 => std_logic_vector(to_unsigned(100,8) ,
19829	 => std_logic_vector(to_unsigned(109,8) ,
19830	 => std_logic_vector(to_unsigned(115,8) ,
19831	 => std_logic_vector(to_unsigned(108,8) ,
19832	 => std_logic_vector(to_unsigned(104,8) ,
19833	 => std_logic_vector(to_unsigned(99,8) ,
19834	 => std_logic_vector(to_unsigned(107,8) ,
19835	 => std_logic_vector(to_unsigned(105,8) ,
19836	 => std_logic_vector(to_unsigned(95,8) ,
19837	 => std_logic_vector(to_unsigned(100,8) ,
19838	 => std_logic_vector(to_unsigned(104,8) ,
19839	 => std_logic_vector(to_unsigned(96,8) ,
19840	 => std_logic_vector(to_unsigned(97,8) ,
19841	 => std_logic_vector(to_unsigned(149,8) ,
19842	 => std_logic_vector(to_unsigned(152,8) ,
19843	 => std_logic_vector(to_unsigned(151,8) ,
19844	 => std_logic_vector(to_unsigned(149,8) ,
19845	 => std_logic_vector(to_unsigned(151,8) ,
19846	 => std_logic_vector(to_unsigned(151,8) ,
19847	 => std_logic_vector(to_unsigned(152,8) ,
19848	 => std_logic_vector(to_unsigned(156,8) ,
19849	 => std_logic_vector(to_unsigned(154,8) ,
19850	 => std_logic_vector(to_unsigned(157,8) ,
19851	 => std_logic_vector(to_unsigned(152,8) ,
19852	 => std_logic_vector(to_unsigned(159,8) ,
19853	 => std_logic_vector(to_unsigned(147,8) ,
19854	 => std_logic_vector(to_unsigned(12,8) ,
19855	 => std_logic_vector(to_unsigned(0,8) ,
19856	 => std_logic_vector(to_unsigned(3,8) ,
19857	 => std_logic_vector(to_unsigned(3,8) ,
19858	 => std_logic_vector(to_unsigned(3,8) ,
19859	 => std_logic_vector(to_unsigned(3,8) ,
19860	 => std_logic_vector(to_unsigned(2,8) ,
19861	 => std_logic_vector(to_unsigned(4,8) ,
19862	 => std_logic_vector(to_unsigned(1,8) ,
19863	 => std_logic_vector(to_unsigned(3,8) ,
19864	 => std_logic_vector(to_unsigned(27,8) ,
19865	 => std_logic_vector(to_unsigned(4,8) ,
19866	 => std_logic_vector(to_unsigned(1,8) ,
19867	 => std_logic_vector(to_unsigned(13,8) ,
19868	 => std_logic_vector(to_unsigned(23,8) ,
19869	 => std_logic_vector(to_unsigned(1,8) ,
19870	 => std_logic_vector(to_unsigned(4,8) ,
19871	 => std_logic_vector(to_unsigned(4,8) ,
19872	 => std_logic_vector(to_unsigned(4,8) ,
19873	 => std_logic_vector(to_unsigned(13,8) ,
19874	 => std_logic_vector(to_unsigned(17,8) ,
19875	 => std_logic_vector(to_unsigned(6,8) ,
19876	 => std_logic_vector(to_unsigned(8,8) ,
19877	 => std_logic_vector(to_unsigned(43,8) ,
19878	 => std_logic_vector(to_unsigned(171,8) ,
19879	 => std_logic_vector(to_unsigned(175,8) ,
19880	 => std_logic_vector(to_unsigned(152,8) ,
19881	 => std_logic_vector(to_unsigned(156,8) ,
19882	 => std_logic_vector(to_unsigned(152,8) ,
19883	 => std_logic_vector(to_unsigned(152,8) ,
19884	 => std_logic_vector(to_unsigned(156,8) ,
19885	 => std_logic_vector(to_unsigned(154,8) ,
19886	 => std_logic_vector(to_unsigned(157,8) ,
19887	 => std_logic_vector(to_unsigned(157,8) ,
19888	 => std_logic_vector(to_unsigned(163,8) ,
19889	 => std_logic_vector(to_unsigned(161,8) ,
19890	 => std_logic_vector(to_unsigned(157,8) ,
19891	 => std_logic_vector(to_unsigned(159,8) ,
19892	 => std_logic_vector(to_unsigned(164,8) ,
19893	 => std_logic_vector(to_unsigned(163,8) ,
19894	 => std_logic_vector(to_unsigned(156,8) ,
19895	 => std_logic_vector(to_unsigned(190,8) ,
19896	 => std_logic_vector(to_unsigned(86,8) ,
19897	 => std_logic_vector(to_unsigned(1,8) ,
19898	 => std_logic_vector(to_unsigned(1,8) ,
19899	 => std_logic_vector(to_unsigned(2,8) ,
19900	 => std_logic_vector(to_unsigned(1,8) ,
19901	 => std_logic_vector(to_unsigned(3,8) ,
19902	 => std_logic_vector(to_unsigned(8,8) ,
19903	 => std_logic_vector(to_unsigned(5,8) ,
19904	 => std_logic_vector(to_unsigned(2,8) ,
19905	 => std_logic_vector(to_unsigned(5,8) ,
19906	 => std_logic_vector(to_unsigned(8,8) ,
19907	 => std_logic_vector(to_unsigned(18,8) ,
19908	 => std_logic_vector(to_unsigned(10,8) ,
19909	 => std_logic_vector(to_unsigned(16,8) ,
19910	 => std_logic_vector(to_unsigned(136,8) ,
19911	 => std_logic_vector(to_unsigned(184,8) ,
19912	 => std_logic_vector(to_unsigned(164,8) ,
19913	 => std_logic_vector(to_unsigned(170,8) ,
19914	 => std_logic_vector(to_unsigned(171,8) ,
19915	 => std_logic_vector(to_unsigned(170,8) ,
19916	 => std_logic_vector(to_unsigned(166,8) ,
19917	 => std_logic_vector(to_unsigned(170,8) ,
19918	 => std_logic_vector(to_unsigned(170,8) ,
19919	 => std_logic_vector(to_unsigned(163,8) ,
19920	 => std_logic_vector(to_unsigned(163,8) ,
19921	 => std_logic_vector(to_unsigned(166,8) ,
19922	 => std_logic_vector(to_unsigned(164,8) ,
19923	 => std_logic_vector(to_unsigned(166,8) ,
19924	 => std_logic_vector(to_unsigned(166,8) ,
19925	 => std_logic_vector(to_unsigned(164,8) ,
19926	 => std_logic_vector(to_unsigned(170,8) ,
19927	 => std_logic_vector(to_unsigned(157,8) ,
19928	 => std_logic_vector(to_unsigned(166,8) ,
19929	 => std_logic_vector(to_unsigned(92,8) ,
19930	 => std_logic_vector(to_unsigned(5,8) ,
19931	 => std_logic_vector(to_unsigned(3,8) ,
19932	 => std_logic_vector(to_unsigned(7,8) ,
19933	 => std_logic_vector(to_unsigned(8,8) ,
19934	 => std_logic_vector(to_unsigned(7,8) ,
19935	 => std_logic_vector(to_unsigned(6,8) ,
19936	 => std_logic_vector(to_unsigned(7,8) ,
19937	 => std_logic_vector(to_unsigned(22,8) ,
19938	 => std_logic_vector(to_unsigned(20,8) ,
19939	 => std_logic_vector(to_unsigned(5,8) ,
19940	 => std_logic_vector(to_unsigned(7,8) ,
19941	 => std_logic_vector(to_unsigned(26,8) ,
19942	 => std_logic_vector(to_unsigned(101,8) ,
19943	 => std_logic_vector(to_unsigned(173,8) ,
19944	 => std_logic_vector(to_unsigned(171,8) ,
19945	 => std_logic_vector(to_unsigned(166,8) ,
19946	 => std_logic_vector(to_unsigned(173,8) ,
19947	 => std_logic_vector(to_unsigned(173,8) ,
19948	 => std_logic_vector(to_unsigned(168,8) ,
19949	 => std_logic_vector(to_unsigned(170,8) ,
19950	 => std_logic_vector(to_unsigned(166,8) ,
19951	 => std_logic_vector(to_unsigned(159,8) ,
19952	 => std_logic_vector(to_unsigned(157,8) ,
19953	 => std_logic_vector(to_unsigned(152,8) ,
19954	 => std_logic_vector(to_unsigned(151,8) ,
19955	 => std_logic_vector(to_unsigned(168,8) ,
19956	 => std_logic_vector(to_unsigned(166,8) ,
19957	 => std_logic_vector(to_unsigned(166,8) ,
19958	 => std_logic_vector(to_unsigned(170,8) ,
19959	 => std_logic_vector(to_unsigned(171,8) ,
19960	 => std_logic_vector(to_unsigned(168,8) ,
19961	 => std_logic_vector(to_unsigned(166,8) ,
19962	 => std_logic_vector(to_unsigned(161,8) ,
19963	 => std_logic_vector(to_unsigned(159,8) ,
19964	 => std_logic_vector(to_unsigned(156,8) ,
19965	 => std_logic_vector(to_unsigned(157,8) ,
19966	 => std_logic_vector(to_unsigned(159,8) ,
19967	 => std_logic_vector(to_unsigned(157,8) ,
19968	 => std_logic_vector(to_unsigned(149,8) ,
19969	 => std_logic_vector(to_unsigned(142,8) ,
19970	 => std_logic_vector(to_unsigned(122,8) ,
19971	 => std_logic_vector(to_unsigned(114,8) ,
19972	 => std_logic_vector(to_unsigned(125,8) ,
19973	 => std_logic_vector(to_unsigned(138,8) ,
19974	 => std_logic_vector(to_unsigned(146,8) ,
19975	 => std_logic_vector(to_unsigned(146,8) ,
19976	 => std_logic_vector(to_unsigned(131,8) ,
19977	 => std_logic_vector(to_unsigned(130,8) ,
19978	 => std_logic_vector(to_unsigned(142,8) ,
19979	 => std_logic_vector(to_unsigned(122,8) ,
19980	 => std_logic_vector(to_unsigned(109,8) ,
19981	 => std_logic_vector(to_unsigned(119,8) ,
19982	 => std_logic_vector(to_unsigned(121,8) ,
19983	 => std_logic_vector(to_unsigned(121,8) ,
19984	 => std_logic_vector(to_unsigned(121,8) ,
19985	 => std_logic_vector(to_unsigned(99,8) ,
19986	 => std_logic_vector(to_unsigned(90,8) ,
19987	 => std_logic_vector(to_unsigned(95,8) ,
19988	 => std_logic_vector(to_unsigned(112,8) ,
19989	 => std_logic_vector(to_unsigned(128,8) ,
19990	 => std_logic_vector(to_unsigned(131,8) ,
19991	 => std_logic_vector(to_unsigned(115,8) ,
19992	 => std_logic_vector(to_unsigned(124,8) ,
19993	 => std_logic_vector(to_unsigned(152,8) ,
19994	 => std_logic_vector(to_unsigned(157,8) ,
19995	 => std_logic_vector(to_unsigned(154,8) ,
19996	 => std_logic_vector(to_unsigned(154,8) ,
19997	 => std_logic_vector(to_unsigned(152,8) ,
19998	 => std_logic_vector(to_unsigned(134,8) ,
19999	 => std_logic_vector(to_unsigned(108,8) ,
20000	 => std_logic_vector(to_unsigned(114,8) ,
20001	 => std_logic_vector(to_unsigned(31,8) ,
20002	 => std_logic_vector(to_unsigned(0,8) ,
20003	 => std_logic_vector(to_unsigned(0,8) ,
20004	 => std_logic_vector(to_unsigned(6,8) ,
20005	 => std_logic_vector(to_unsigned(57,8) ,
20006	 => std_logic_vector(to_unsigned(104,8) ,
20007	 => std_logic_vector(to_unsigned(84,8) ,
20008	 => std_logic_vector(to_unsigned(46,8) ,
20009	 => std_logic_vector(to_unsigned(12,8) ,
20010	 => std_logic_vector(to_unsigned(2,8) ,
20011	 => std_logic_vector(to_unsigned(1,8) ,
20012	 => std_logic_vector(to_unsigned(0,8) ,
20013	 => std_logic_vector(to_unsigned(0,8) ,
20014	 => std_logic_vector(to_unsigned(2,8) ,
20015	 => std_logic_vector(to_unsigned(4,8) ,
20016	 => std_logic_vector(to_unsigned(3,8) ,
20017	 => std_logic_vector(to_unsigned(59,8) ,
20018	 => std_logic_vector(to_unsigned(96,8) ,
20019	 => std_logic_vector(to_unsigned(108,8) ,
20020	 => std_logic_vector(to_unsigned(141,8) ,
20021	 => std_logic_vector(to_unsigned(108,8) ,
20022	 => std_logic_vector(to_unsigned(96,8) ,
20023	 => std_logic_vector(to_unsigned(92,8) ,
20024	 => std_logic_vector(to_unsigned(74,8) ,
20025	 => std_logic_vector(to_unsigned(76,8) ,
20026	 => std_logic_vector(to_unsigned(76,8) ,
20027	 => std_logic_vector(to_unsigned(79,8) ,
20028	 => std_logic_vector(to_unsigned(69,8) ,
20029	 => std_logic_vector(to_unsigned(69,8) ,
20030	 => std_logic_vector(to_unsigned(72,8) ,
20031	 => std_logic_vector(to_unsigned(73,8) ,
20032	 => std_logic_vector(to_unsigned(72,8) ,
20033	 => std_logic_vector(to_unsigned(65,8) ,
20034	 => std_logic_vector(to_unsigned(76,8) ,
20035	 => std_logic_vector(to_unsigned(74,8) ,
20036	 => std_logic_vector(to_unsigned(65,8) ,
20037	 => std_logic_vector(to_unsigned(77,8) ,
20038	 => std_logic_vector(to_unsigned(104,8) ,
20039	 => std_logic_vector(to_unsigned(107,8) ,
20040	 => std_logic_vector(to_unsigned(99,8) ,
20041	 => std_logic_vector(to_unsigned(88,8) ,
20042	 => std_logic_vector(to_unsigned(77,8) ,
20043	 => std_logic_vector(to_unsigned(72,8) ,
20044	 => std_logic_vector(to_unsigned(63,8) ,
20045	 => std_logic_vector(to_unsigned(69,8) ,
20046	 => std_logic_vector(to_unsigned(76,8) ,
20047	 => std_logic_vector(to_unsigned(71,8) ,
20048	 => std_logic_vector(to_unsigned(72,8) ,
20049	 => std_logic_vector(to_unsigned(74,8) ,
20050	 => std_logic_vector(to_unsigned(70,8) ,
20051	 => std_logic_vector(to_unsigned(65,8) ,
20052	 => std_logic_vector(to_unsigned(64,8) ,
20053	 => std_logic_vector(to_unsigned(61,8) ,
20054	 => std_logic_vector(to_unsigned(70,8) ,
20055	 => std_logic_vector(to_unsigned(66,8) ,
20056	 => std_logic_vector(to_unsigned(60,8) ,
20057	 => std_logic_vector(to_unsigned(76,8) ,
20058	 => std_logic_vector(to_unsigned(80,8) ,
20059	 => std_logic_vector(to_unsigned(71,8) ,
20060	 => std_logic_vector(to_unsigned(82,8) ,
20061	 => std_logic_vector(to_unsigned(86,8) ,
20062	 => std_logic_vector(to_unsigned(77,8) ,
20063	 => std_logic_vector(to_unsigned(91,8) ,
20064	 => std_logic_vector(to_unsigned(29,8) ,
20065	 => std_logic_vector(to_unsigned(8,8) ,
20066	 => std_logic_vector(to_unsigned(24,8) ,
20067	 => std_logic_vector(to_unsigned(30,8) ,
20068	 => std_logic_vector(to_unsigned(22,8) ,
20069	 => std_logic_vector(to_unsigned(34,8) ,
20070	 => std_logic_vector(to_unsigned(62,8) ,
20071	 => std_logic_vector(to_unsigned(78,8) ,
20072	 => std_logic_vector(to_unsigned(88,8) ,
20073	 => std_logic_vector(to_unsigned(93,8) ,
20074	 => std_logic_vector(to_unsigned(101,8) ,
20075	 => std_logic_vector(to_unsigned(100,8) ,
20076	 => std_logic_vector(to_unsigned(100,8) ,
20077	 => std_logic_vector(to_unsigned(122,8) ,
20078	 => std_logic_vector(to_unsigned(136,8) ,
20079	 => std_logic_vector(to_unsigned(147,8) ,
20080	 => std_logic_vector(to_unsigned(142,8) ,
20081	 => std_logic_vector(to_unsigned(141,8) ,
20082	 => std_logic_vector(to_unsigned(142,8) ,
20083	 => std_logic_vector(to_unsigned(146,8) ,
20084	 => std_logic_vector(to_unsigned(152,8) ,
20085	 => std_logic_vector(to_unsigned(103,8) ,
20086	 => std_logic_vector(to_unsigned(70,8) ,
20087	 => std_logic_vector(to_unsigned(72,8) ,
20088	 => std_logic_vector(to_unsigned(67,8) ,
20089	 => std_logic_vector(to_unsigned(72,8) ,
20090	 => std_logic_vector(to_unsigned(79,8) ,
20091	 => std_logic_vector(to_unsigned(9,8) ,
20092	 => std_logic_vector(to_unsigned(0,8) ,
20093	 => std_logic_vector(to_unsigned(0,8) ,
20094	 => std_logic_vector(to_unsigned(35,8) ,
20095	 => std_logic_vector(to_unsigned(147,8) ,
20096	 => std_logic_vector(to_unsigned(133,8) ,
20097	 => std_logic_vector(to_unsigned(116,8) ,
20098	 => std_logic_vector(to_unsigned(138,8) ,
20099	 => std_logic_vector(to_unsigned(128,8) ,
20100	 => std_logic_vector(to_unsigned(100,8) ,
20101	 => std_logic_vector(to_unsigned(101,8) ,
20102	 => std_logic_vector(to_unsigned(108,8) ,
20103	 => std_logic_vector(to_unsigned(99,8) ,
20104	 => std_logic_vector(to_unsigned(100,8) ,
20105	 => std_logic_vector(to_unsigned(109,8) ,
20106	 => std_logic_vector(to_unsigned(108,8) ,
20107	 => std_logic_vector(to_unsigned(108,8) ,
20108	 => std_logic_vector(to_unsigned(99,8) ,
20109	 => std_logic_vector(to_unsigned(92,8) ,
20110	 => std_logic_vector(to_unsigned(86,8) ,
20111	 => std_logic_vector(to_unsigned(85,8) ,
20112	 => std_logic_vector(to_unsigned(76,8) ,
20113	 => std_logic_vector(to_unsigned(78,8) ,
20114	 => std_logic_vector(to_unsigned(69,8) ,
20115	 => std_logic_vector(to_unsigned(15,8) ,
20116	 => std_logic_vector(to_unsigned(0,8) ,
20117	 => std_logic_vector(to_unsigned(0,8) ,
20118	 => std_logic_vector(to_unsigned(1,8) ,
20119	 => std_logic_vector(to_unsigned(1,8) ,
20120	 => std_logic_vector(to_unsigned(1,8) ,
20121	 => std_logic_vector(to_unsigned(1,8) ,
20122	 => std_logic_vector(to_unsigned(0,8) ,
20123	 => std_logic_vector(to_unsigned(1,8) ,
20124	 => std_logic_vector(to_unsigned(3,8) ,
20125	 => std_logic_vector(to_unsigned(1,8) ,
20126	 => std_logic_vector(to_unsigned(3,8) ,
20127	 => std_logic_vector(to_unsigned(29,8) ,
20128	 => std_logic_vector(to_unsigned(45,8) ,
20129	 => std_logic_vector(to_unsigned(71,8) ,
20130	 => std_logic_vector(to_unsigned(105,8) ,
20131	 => std_logic_vector(to_unsigned(108,8) ,
20132	 => std_logic_vector(to_unsigned(101,8) ,
20133	 => std_logic_vector(to_unsigned(95,8) ,
20134	 => std_logic_vector(to_unsigned(108,8) ,
20135	 => std_logic_vector(to_unsigned(130,8) ,
20136	 => std_logic_vector(to_unsigned(136,8) ,
20137	 => std_logic_vector(to_unsigned(139,8) ,
20138	 => std_logic_vector(to_unsigned(134,8) ,
20139	 => std_logic_vector(to_unsigned(144,8) ,
20140	 => std_logic_vector(to_unsigned(157,8) ,
20141	 => std_logic_vector(to_unsigned(156,8) ,
20142	 => std_logic_vector(to_unsigned(154,8) ,
20143	 => std_logic_vector(to_unsigned(142,8) ,
20144	 => std_logic_vector(to_unsigned(116,8) ,
20145	 => std_logic_vector(to_unsigned(100,8) ,
20146	 => std_logic_vector(to_unsigned(109,8) ,
20147	 => std_logic_vector(to_unsigned(122,8) ,
20148	 => std_logic_vector(to_unsigned(119,8) ,
20149	 => std_logic_vector(to_unsigned(116,8) ,
20150	 => std_logic_vector(to_unsigned(118,8) ,
20151	 => std_logic_vector(to_unsigned(108,8) ,
20152	 => std_logic_vector(to_unsigned(112,8) ,
20153	 => std_logic_vector(to_unsigned(112,8) ,
20154	 => std_logic_vector(to_unsigned(109,8) ,
20155	 => std_logic_vector(to_unsigned(108,8) ,
20156	 => std_logic_vector(to_unsigned(95,8) ,
20157	 => std_logic_vector(to_unsigned(101,8) ,
20158	 => std_logic_vector(to_unsigned(109,8) ,
20159	 => std_logic_vector(to_unsigned(97,8) ,
20160	 => std_logic_vector(to_unsigned(93,8) ,
20161	 => std_logic_vector(to_unsigned(152,8) ,
20162	 => std_logic_vector(to_unsigned(156,8) ,
20163	 => std_logic_vector(to_unsigned(156,8) ,
20164	 => std_logic_vector(to_unsigned(157,8) ,
20165	 => std_logic_vector(to_unsigned(164,8) ,
20166	 => std_logic_vector(to_unsigned(159,8) ,
20167	 => std_logic_vector(to_unsigned(159,8) ,
20168	 => std_logic_vector(to_unsigned(161,8) ,
20169	 => std_logic_vector(to_unsigned(163,8) ,
20170	 => std_logic_vector(to_unsigned(161,8) ,
20171	 => std_logic_vector(to_unsigned(154,8) ,
20172	 => std_logic_vector(to_unsigned(159,8) ,
20173	 => std_logic_vector(to_unsigned(146,8) ,
20174	 => std_logic_vector(to_unsigned(13,8) ,
20175	 => std_logic_vector(to_unsigned(0,8) ,
20176	 => std_logic_vector(to_unsigned(8,8) ,
20177	 => std_logic_vector(to_unsigned(12,8) ,
20178	 => std_logic_vector(to_unsigned(1,8) ,
20179	 => std_logic_vector(to_unsigned(0,8) ,
20180	 => std_logic_vector(to_unsigned(1,8) ,
20181	 => std_logic_vector(to_unsigned(2,8) ,
20182	 => std_logic_vector(to_unsigned(5,8) ,
20183	 => std_logic_vector(to_unsigned(3,8) ,
20184	 => std_logic_vector(to_unsigned(27,8) ,
20185	 => std_logic_vector(to_unsigned(44,8) ,
20186	 => std_logic_vector(to_unsigned(37,8) ,
20187	 => std_logic_vector(to_unsigned(30,8) ,
20188	 => std_logic_vector(to_unsigned(46,8) ,
20189	 => std_logic_vector(to_unsigned(18,8) ,
20190	 => std_logic_vector(to_unsigned(9,8) ,
20191	 => std_logic_vector(to_unsigned(5,8) ,
20192	 => std_logic_vector(to_unsigned(4,8) ,
20193	 => std_logic_vector(to_unsigned(10,8) ,
20194	 => std_logic_vector(to_unsigned(27,8) ,
20195	 => std_logic_vector(to_unsigned(23,8) ,
20196	 => std_logic_vector(to_unsigned(10,8) ,
20197	 => std_logic_vector(to_unsigned(19,8) ,
20198	 => std_logic_vector(to_unsigned(48,8) ,
20199	 => std_logic_vector(to_unsigned(118,8) ,
20200	 => std_logic_vector(to_unsigned(177,8) ,
20201	 => std_logic_vector(to_unsigned(159,8) ,
20202	 => std_logic_vector(to_unsigned(157,8) ,
20203	 => std_logic_vector(to_unsigned(156,8) ,
20204	 => std_logic_vector(to_unsigned(157,8) ,
20205	 => std_logic_vector(to_unsigned(159,8) ,
20206	 => std_logic_vector(to_unsigned(163,8) ,
20207	 => std_logic_vector(to_unsigned(159,8) ,
20208	 => std_logic_vector(to_unsigned(161,8) ,
20209	 => std_logic_vector(to_unsigned(163,8) ,
20210	 => std_logic_vector(to_unsigned(159,8) ,
20211	 => std_logic_vector(to_unsigned(159,8) ,
20212	 => std_logic_vector(to_unsigned(164,8) ,
20213	 => std_logic_vector(to_unsigned(166,8) ,
20214	 => std_logic_vector(to_unsigned(163,8) ,
20215	 => std_logic_vector(to_unsigned(166,8) ,
20216	 => std_logic_vector(to_unsigned(156,8) ,
20217	 => std_logic_vector(to_unsigned(18,8) ,
20218	 => std_logic_vector(to_unsigned(1,8) ,
20219	 => std_logic_vector(to_unsigned(5,8) ,
20220	 => std_logic_vector(to_unsigned(6,8) ,
20221	 => std_logic_vector(to_unsigned(7,8) ,
20222	 => std_logic_vector(to_unsigned(4,8) ,
20223	 => std_logic_vector(to_unsigned(5,8) ,
20224	 => std_logic_vector(to_unsigned(5,8) ,
20225	 => std_logic_vector(to_unsigned(15,8) ,
20226	 => std_logic_vector(to_unsigned(25,8) ,
20227	 => std_logic_vector(to_unsigned(17,8) ,
20228	 => std_logic_vector(to_unsigned(8,8) ,
20229	 => std_logic_vector(to_unsigned(4,8) ,
20230	 => std_logic_vector(to_unsigned(73,8) ,
20231	 => std_logic_vector(to_unsigned(181,8) ,
20232	 => std_logic_vector(to_unsigned(163,8) ,
20233	 => std_logic_vector(to_unsigned(170,8) ,
20234	 => std_logic_vector(to_unsigned(173,8) ,
20235	 => std_logic_vector(to_unsigned(173,8) ,
20236	 => std_logic_vector(to_unsigned(171,8) ,
20237	 => std_logic_vector(to_unsigned(170,8) ,
20238	 => std_logic_vector(to_unsigned(170,8) ,
20239	 => std_logic_vector(to_unsigned(166,8) ,
20240	 => std_logic_vector(to_unsigned(163,8) ,
20241	 => std_logic_vector(to_unsigned(168,8) ,
20242	 => std_logic_vector(to_unsigned(163,8) ,
20243	 => std_logic_vector(to_unsigned(163,8) ,
20244	 => std_logic_vector(to_unsigned(166,8) ,
20245	 => std_logic_vector(to_unsigned(164,8) ,
20246	 => std_logic_vector(to_unsigned(168,8) ,
20247	 => std_logic_vector(to_unsigned(161,8) ,
20248	 => std_logic_vector(to_unsigned(149,8) ,
20249	 => std_logic_vector(to_unsigned(138,8) ,
20250	 => std_logic_vector(to_unsigned(57,8) ,
20251	 => std_logic_vector(to_unsigned(4,8) ,
20252	 => std_logic_vector(to_unsigned(3,8) ,
20253	 => std_logic_vector(to_unsigned(6,8) ,
20254	 => std_logic_vector(to_unsigned(7,8) ,
20255	 => std_logic_vector(to_unsigned(6,8) ,
20256	 => std_logic_vector(to_unsigned(6,8) ,
20257	 => std_logic_vector(to_unsigned(5,8) ,
20258	 => std_logic_vector(to_unsigned(4,8) ,
20259	 => std_logic_vector(to_unsigned(8,8) ,
20260	 => std_logic_vector(to_unsigned(14,8) ,
20261	 => std_logic_vector(to_unsigned(16,8) ,
20262	 => std_logic_vector(to_unsigned(33,8) ,
20263	 => std_logic_vector(to_unsigned(166,8) ,
20264	 => std_logic_vector(to_unsigned(181,8) ,
20265	 => std_logic_vector(to_unsigned(166,8) ,
20266	 => std_logic_vector(to_unsigned(173,8) ,
20267	 => std_logic_vector(to_unsigned(171,8) ,
20268	 => std_logic_vector(to_unsigned(170,8) ,
20269	 => std_logic_vector(to_unsigned(173,8) ,
20270	 => std_logic_vector(to_unsigned(170,8) ,
20271	 => std_logic_vector(to_unsigned(171,8) ,
20272	 => std_logic_vector(to_unsigned(170,8) ,
20273	 => std_logic_vector(to_unsigned(166,8) ,
20274	 => std_logic_vector(to_unsigned(161,8) ,
20275	 => std_logic_vector(to_unsigned(166,8) ,
20276	 => std_logic_vector(to_unsigned(166,8) ,
20277	 => std_logic_vector(to_unsigned(166,8) ,
20278	 => std_logic_vector(to_unsigned(163,8) ,
20279	 => std_logic_vector(to_unsigned(138,8) ,
20280	 => std_logic_vector(to_unsigned(144,8) ,
20281	 => std_logic_vector(to_unsigned(159,8) ,
20282	 => std_logic_vector(to_unsigned(170,8) ,
20283	 => std_logic_vector(to_unsigned(163,8) ,
20284	 => std_logic_vector(to_unsigned(159,8) ,
20285	 => std_logic_vector(to_unsigned(164,8) ,
20286	 => std_logic_vector(to_unsigned(156,8) ,
20287	 => std_logic_vector(to_unsigned(157,8) ,
20288	 => std_logic_vector(to_unsigned(157,8) ,
20289	 => std_logic_vector(to_unsigned(154,8) ,
20290	 => std_logic_vector(to_unsigned(134,8) ,
20291	 => std_logic_vector(to_unsigned(121,8) ,
20292	 => std_logic_vector(to_unsigned(131,8) ,
20293	 => std_logic_vector(to_unsigned(142,8) ,
20294	 => std_logic_vector(to_unsigned(144,8) ,
20295	 => std_logic_vector(to_unsigned(146,8) ,
20296	 => std_logic_vector(to_unsigned(142,8) ,
20297	 => std_logic_vector(to_unsigned(139,8) ,
20298	 => std_logic_vector(to_unsigned(142,8) ,
20299	 => std_logic_vector(to_unsigned(125,8) ,
20300	 => std_logic_vector(to_unsigned(122,8) ,
20301	 => std_logic_vector(to_unsigned(119,8) ,
20302	 => std_logic_vector(to_unsigned(115,8) ,
20303	 => std_logic_vector(to_unsigned(121,8) ,
20304	 => std_logic_vector(to_unsigned(108,8) ,
20305	 => std_logic_vector(to_unsigned(99,8) ,
20306	 => std_logic_vector(to_unsigned(93,8) ,
20307	 => std_logic_vector(to_unsigned(84,8) ,
20308	 => std_logic_vector(to_unsigned(87,8) ,
20309	 => std_logic_vector(to_unsigned(119,8) ,
20310	 => std_logic_vector(to_unsigned(119,8) ,
20311	 => std_logic_vector(to_unsigned(111,8) ,
20312	 => std_logic_vector(to_unsigned(103,8) ,
20313	 => std_logic_vector(to_unsigned(136,8) ,
20314	 => std_logic_vector(to_unsigned(168,8) ,
20315	 => std_logic_vector(to_unsigned(157,8) ,
20316	 => std_logic_vector(to_unsigned(152,8) ,
20317	 => std_logic_vector(to_unsigned(154,8) ,
20318	 => std_logic_vector(to_unsigned(151,8) ,
20319	 => std_logic_vector(to_unsigned(118,8) ,
20320	 => std_logic_vector(to_unsigned(111,8) ,
20321	 => std_logic_vector(to_unsigned(87,8) ,
20322	 => std_logic_vector(to_unsigned(37,8) ,
20323	 => std_logic_vector(to_unsigned(36,8) ,
20324	 => std_logic_vector(to_unsigned(22,8) ,
20325	 => std_logic_vector(to_unsigned(2,8) ,
20326	 => std_logic_vector(to_unsigned(9,8) ,
20327	 => std_logic_vector(to_unsigned(16,8) ,
20328	 => std_logic_vector(to_unsigned(11,8) ,
20329	 => std_logic_vector(to_unsigned(2,8) ,
20330	 => std_logic_vector(to_unsigned(0,8) ,
20331	 => std_logic_vector(to_unsigned(1,8) ,
20332	 => std_logic_vector(to_unsigned(2,8) ,
20333	 => std_logic_vector(to_unsigned(2,8) ,
20334	 => std_logic_vector(to_unsigned(2,8) ,
20335	 => std_logic_vector(to_unsigned(3,8) ,
20336	 => std_logic_vector(to_unsigned(8,8) ,
20337	 => std_logic_vector(to_unsigned(107,8) ,
20338	 => std_logic_vector(to_unsigned(152,8) ,
20339	 => std_logic_vector(to_unsigned(147,8) ,
20340	 => std_logic_vector(to_unsigned(134,8) ,
20341	 => std_logic_vector(to_unsigned(114,8) ,
20342	 => std_logic_vector(to_unsigned(99,8) ,
20343	 => std_logic_vector(to_unsigned(107,8) ,
20344	 => std_logic_vector(to_unsigned(88,8) ,
20345	 => std_logic_vector(to_unsigned(79,8) ,
20346	 => std_logic_vector(to_unsigned(80,8) ,
20347	 => std_logic_vector(to_unsigned(79,8) ,
20348	 => std_logic_vector(to_unsigned(72,8) ,
20349	 => std_logic_vector(to_unsigned(77,8) ,
20350	 => std_logic_vector(to_unsigned(79,8) ,
20351	 => std_logic_vector(to_unsigned(77,8) ,
20352	 => std_logic_vector(to_unsigned(78,8) ,
20353	 => std_logic_vector(to_unsigned(76,8) ,
20354	 => std_logic_vector(to_unsigned(72,8) ,
20355	 => std_logic_vector(to_unsigned(77,8) ,
20356	 => std_logic_vector(to_unsigned(85,8) ,
20357	 => std_logic_vector(to_unsigned(64,8) ,
20358	 => std_logic_vector(to_unsigned(69,8) ,
20359	 => std_logic_vector(to_unsigned(56,8) ,
20360	 => std_logic_vector(to_unsigned(47,8) ,
20361	 => std_logic_vector(to_unsigned(70,8) ,
20362	 => std_logic_vector(to_unsigned(80,8) ,
20363	 => std_logic_vector(to_unsigned(72,8) ,
20364	 => std_logic_vector(to_unsigned(77,8) ,
20365	 => std_logic_vector(to_unsigned(81,8) ,
20366	 => std_logic_vector(to_unsigned(79,8) ,
20367	 => std_logic_vector(to_unsigned(78,8) ,
20368	 => std_logic_vector(to_unsigned(86,8) ,
20369	 => std_logic_vector(to_unsigned(91,8) ,
20370	 => std_logic_vector(to_unsigned(81,8) ,
20371	 => std_logic_vector(to_unsigned(78,8) ,
20372	 => std_logic_vector(to_unsigned(81,8) ,
20373	 => std_logic_vector(to_unsigned(73,8) ,
20374	 => std_logic_vector(to_unsigned(74,8) ,
20375	 => std_logic_vector(to_unsigned(79,8) ,
20376	 => std_logic_vector(to_unsigned(77,8) ,
20377	 => std_logic_vector(to_unsigned(82,8) ,
20378	 => std_logic_vector(to_unsigned(84,8) ,
20379	 => std_logic_vector(to_unsigned(80,8) ,
20380	 => std_logic_vector(to_unsigned(90,8) ,
20381	 => std_logic_vector(to_unsigned(88,8) ,
20382	 => std_logic_vector(to_unsigned(103,8) ,
20383	 => std_logic_vector(to_unsigned(78,8) ,
20384	 => std_logic_vector(to_unsigned(19,8) ,
20385	 => std_logic_vector(to_unsigned(12,8) ,
20386	 => std_logic_vector(to_unsigned(7,8) ,
20387	 => std_logic_vector(to_unsigned(8,8) ,
20388	 => std_logic_vector(to_unsigned(16,8) ,
20389	 => std_logic_vector(to_unsigned(27,8) ,
20390	 => std_logic_vector(to_unsigned(37,8) ,
20391	 => std_logic_vector(to_unsigned(47,8) ,
20392	 => std_logic_vector(to_unsigned(67,8) ,
20393	 => std_logic_vector(to_unsigned(53,8) ,
20394	 => std_logic_vector(to_unsigned(49,8) ,
20395	 => std_logic_vector(to_unsigned(96,8) ,
20396	 => std_logic_vector(to_unsigned(99,8) ,
20397	 => std_logic_vector(to_unsigned(100,8) ,
20398	 => std_logic_vector(to_unsigned(115,8) ,
20399	 => std_logic_vector(to_unsigned(131,8) ,
20400	 => std_logic_vector(to_unsigned(114,8) ,
20401	 => std_logic_vector(to_unsigned(116,8) ,
20402	 => std_logic_vector(to_unsigned(144,8) ,
20403	 => std_logic_vector(to_unsigned(138,8) ,
20404	 => std_logic_vector(to_unsigned(131,8) ,
20405	 => std_logic_vector(to_unsigned(121,8) ,
20406	 => std_logic_vector(to_unsigned(82,8) ,
20407	 => std_logic_vector(to_unsigned(78,8) ,
20408	 => std_logic_vector(to_unsigned(76,8) ,
20409	 => std_logic_vector(to_unsigned(79,8) ,
20410	 => std_logic_vector(to_unsigned(90,8) ,
20411	 => std_logic_vector(to_unsigned(23,8) ,
20412	 => std_logic_vector(to_unsigned(0,8) ,
20413	 => std_logic_vector(to_unsigned(0,8) ,
20414	 => std_logic_vector(to_unsigned(18,8) ,
20415	 => std_logic_vector(to_unsigned(108,8) ,
20416	 => std_logic_vector(to_unsigned(91,8) ,
20417	 => std_logic_vector(to_unsigned(99,8) ,
20418	 => std_logic_vector(to_unsigned(125,8) ,
20419	 => std_logic_vector(to_unsigned(112,8) ,
20420	 => std_logic_vector(to_unsigned(99,8) ,
20421	 => std_logic_vector(to_unsigned(114,8) ,
20422	 => std_logic_vector(to_unsigned(112,8) ,
20423	 => std_logic_vector(to_unsigned(104,8) ,
20424	 => std_logic_vector(to_unsigned(104,8) ,
20425	 => std_logic_vector(to_unsigned(114,8) ,
20426	 => std_logic_vector(to_unsigned(111,8) ,
20427	 => std_logic_vector(to_unsigned(103,8) ,
20428	 => std_logic_vector(to_unsigned(99,8) ,
20429	 => std_logic_vector(to_unsigned(93,8) ,
20430	 => std_logic_vector(to_unsigned(87,8) ,
20431	 => std_logic_vector(to_unsigned(87,8) ,
20432	 => std_logic_vector(to_unsigned(90,8) ,
20433	 => std_logic_vector(to_unsigned(67,8) ,
20434	 => std_logic_vector(to_unsigned(8,8) ,
20435	 => std_logic_vector(to_unsigned(0,8) ,
20436	 => std_logic_vector(to_unsigned(1,8) ,
20437	 => std_logic_vector(to_unsigned(1,8) ,
20438	 => std_logic_vector(to_unsigned(0,8) ,
20439	 => std_logic_vector(to_unsigned(0,8) ,
20440	 => std_logic_vector(to_unsigned(0,8) ,
20441	 => std_logic_vector(to_unsigned(0,8) ,
20442	 => std_logic_vector(to_unsigned(0,8) ,
20443	 => std_logic_vector(to_unsigned(0,8) ,
20444	 => std_logic_vector(to_unsigned(1,8) ,
20445	 => std_logic_vector(to_unsigned(2,8) ,
20446	 => std_logic_vector(to_unsigned(1,8) ,
20447	 => std_logic_vector(to_unsigned(1,8) ,
20448	 => std_logic_vector(to_unsigned(11,8) ,
20449	 => std_logic_vector(to_unsigned(76,8) ,
20450	 => std_logic_vector(to_unsigned(108,8) ,
20451	 => std_logic_vector(to_unsigned(97,8) ,
20452	 => std_logic_vector(to_unsigned(97,8) ,
20453	 => std_logic_vector(to_unsigned(95,8) ,
20454	 => std_logic_vector(to_unsigned(100,8) ,
20455	 => std_logic_vector(to_unsigned(112,8) ,
20456	 => std_logic_vector(to_unsigned(115,8) ,
20457	 => std_logic_vector(to_unsigned(108,8) ,
20458	 => std_logic_vector(to_unsigned(96,8) ,
20459	 => std_logic_vector(to_unsigned(109,8) ,
20460	 => std_logic_vector(to_unsigned(154,8) ,
20461	 => std_logic_vector(to_unsigned(168,8) ,
20462	 => std_logic_vector(to_unsigned(164,8) ,
20463	 => std_logic_vector(to_unsigned(164,8) ,
20464	 => std_logic_vector(to_unsigned(142,8) ,
20465	 => std_logic_vector(to_unsigned(112,8) ,
20466	 => std_logic_vector(to_unsigned(128,8) ,
20467	 => std_logic_vector(to_unsigned(141,8) ,
20468	 => std_logic_vector(to_unsigned(128,8) ,
20469	 => std_logic_vector(to_unsigned(121,8) ,
20470	 => std_logic_vector(to_unsigned(108,8) ,
20471	 => std_logic_vector(to_unsigned(101,8) ,
20472	 => std_logic_vector(to_unsigned(101,8) ,
20473	 => std_logic_vector(to_unsigned(108,8) ,
20474	 => std_logic_vector(to_unsigned(99,8) ,
20475	 => std_logic_vector(to_unsigned(88,8) ,
20476	 => std_logic_vector(to_unsigned(88,8) ,
20477	 => std_logic_vector(to_unsigned(87,8) ,
20478	 => std_logic_vector(to_unsigned(90,8) ,
20479	 => std_logic_vector(to_unsigned(91,8) ,
20480	 => std_logic_vector(to_unsigned(85,8) ,
20481	 => std_logic_vector(to_unsigned(146,8) ,
20482	 => std_logic_vector(to_unsigned(141,8) ,
20483	 => std_logic_vector(to_unsigned(142,8) ,
20484	 => std_logic_vector(to_unsigned(152,8) ,
20485	 => std_logic_vector(to_unsigned(164,8) ,
20486	 => std_logic_vector(to_unsigned(161,8) ,
20487	 => std_logic_vector(to_unsigned(163,8) ,
20488	 => std_logic_vector(to_unsigned(161,8) ,
20489	 => std_logic_vector(to_unsigned(159,8) ,
20490	 => std_logic_vector(to_unsigned(164,8) ,
20491	 => std_logic_vector(to_unsigned(163,8) ,
20492	 => std_logic_vector(to_unsigned(163,8) ,
20493	 => std_logic_vector(to_unsigned(198,8) ,
20494	 => std_logic_vector(to_unsigned(35,8) ,
20495	 => std_logic_vector(to_unsigned(0,8) ,
20496	 => std_logic_vector(to_unsigned(23,8) ,
20497	 => std_logic_vector(to_unsigned(42,8) ,
20498	 => std_logic_vector(to_unsigned(15,8) ,
20499	 => std_logic_vector(to_unsigned(5,8) ,
20500	 => std_logic_vector(to_unsigned(3,8) ,
20501	 => std_logic_vector(to_unsigned(5,8) ,
20502	 => std_logic_vector(to_unsigned(11,8) ,
20503	 => std_logic_vector(to_unsigned(5,8) ,
20504	 => std_logic_vector(to_unsigned(2,8) ,
20505	 => std_logic_vector(to_unsigned(60,8) ,
20506	 => std_logic_vector(to_unsigned(114,8) ,
20507	 => std_logic_vector(to_unsigned(21,8) ,
20508	 => std_logic_vector(to_unsigned(45,8) ,
20509	 => std_logic_vector(to_unsigned(72,8) ,
20510	 => std_logic_vector(to_unsigned(28,8) ,
20511	 => std_logic_vector(to_unsigned(20,8) ,
20512	 => std_logic_vector(to_unsigned(23,8) ,
20513	 => std_logic_vector(to_unsigned(15,8) ,
20514	 => std_logic_vector(to_unsigned(13,8) ,
20515	 => std_logic_vector(to_unsigned(16,8) ,
20516	 => std_logic_vector(to_unsigned(17,8) ,
20517	 => std_logic_vector(to_unsigned(23,8) ,
20518	 => std_logic_vector(to_unsigned(15,8) ,
20519	 => std_logic_vector(to_unsigned(28,8) ,
20520	 => std_logic_vector(to_unsigned(149,8) ,
20521	 => std_logic_vector(to_unsigned(184,8) ,
20522	 => std_logic_vector(to_unsigned(186,8) ,
20523	 => std_logic_vector(to_unsigned(183,8) ,
20524	 => std_logic_vector(to_unsigned(171,8) ,
20525	 => std_logic_vector(to_unsigned(170,8) ,
20526	 => std_logic_vector(to_unsigned(170,8) ,
20527	 => std_logic_vector(to_unsigned(164,8) ,
20528	 => std_logic_vector(to_unsigned(161,8) ,
20529	 => std_logic_vector(to_unsigned(159,8) ,
20530	 => std_logic_vector(to_unsigned(161,8) ,
20531	 => std_logic_vector(to_unsigned(157,8) ,
20532	 => std_logic_vector(to_unsigned(164,8) ,
20533	 => std_logic_vector(to_unsigned(163,8) ,
20534	 => std_logic_vector(to_unsigned(161,8) ,
20535	 => std_logic_vector(to_unsigned(156,8) ,
20536	 => std_logic_vector(to_unsigned(175,8) ,
20537	 => std_logic_vector(to_unsigned(105,8) ,
20538	 => std_logic_vector(to_unsigned(11,8) ,
20539	 => std_logic_vector(to_unsigned(3,8) ,
20540	 => std_logic_vector(to_unsigned(4,8) ,
20541	 => std_logic_vector(to_unsigned(7,8) ,
20542	 => std_logic_vector(to_unsigned(10,8) ,
20543	 => std_logic_vector(to_unsigned(14,8) ,
20544	 => std_logic_vector(to_unsigned(7,8) ,
20545	 => std_logic_vector(to_unsigned(13,8) ,
20546	 => std_logic_vector(to_unsigned(11,8) ,
20547	 => std_logic_vector(to_unsigned(26,8) ,
20548	 => std_logic_vector(to_unsigned(72,8) ,
20549	 => std_logic_vector(to_unsigned(3,8) ,
20550	 => std_logic_vector(to_unsigned(36,8) ,
20551	 => std_logic_vector(to_unsigned(175,8) ,
20552	 => std_logic_vector(to_unsigned(161,8) ,
20553	 => std_logic_vector(to_unsigned(164,8) ,
20554	 => std_logic_vector(to_unsigned(168,8) ,
20555	 => std_logic_vector(to_unsigned(157,8) ,
20556	 => std_logic_vector(to_unsigned(142,8) ,
20557	 => std_logic_vector(to_unsigned(170,8) ,
20558	 => std_logic_vector(to_unsigned(171,8) ,
20559	 => std_logic_vector(to_unsigned(166,8) ,
20560	 => std_logic_vector(to_unsigned(166,8) ,
20561	 => std_logic_vector(to_unsigned(166,8) ,
20562	 => std_logic_vector(to_unsigned(163,8) ,
20563	 => std_logic_vector(to_unsigned(164,8) ,
20564	 => std_logic_vector(to_unsigned(168,8) ,
20565	 => std_logic_vector(to_unsigned(164,8) ,
20566	 => std_logic_vector(to_unsigned(163,8) ,
20567	 => std_logic_vector(to_unsigned(163,8) ,
20568	 => std_logic_vector(to_unsigned(152,8) ,
20569	 => std_logic_vector(to_unsigned(161,8) ,
20570	 => std_logic_vector(to_unsigned(170,8) ,
20571	 => std_logic_vector(to_unsigned(19,8) ,
20572	 => std_logic_vector(to_unsigned(2,8) ,
20573	 => std_logic_vector(to_unsigned(8,8) ,
20574	 => std_logic_vector(to_unsigned(8,8) ,
20575	 => std_logic_vector(to_unsigned(6,8) ,
20576	 => std_logic_vector(to_unsigned(5,8) ,
20577	 => std_logic_vector(to_unsigned(3,8) ,
20578	 => std_logic_vector(to_unsigned(5,8) ,
20579	 => std_logic_vector(to_unsigned(9,8) ,
20580	 => std_logic_vector(to_unsigned(19,8) ,
20581	 => std_logic_vector(to_unsigned(27,8) ,
20582	 => std_logic_vector(to_unsigned(86,8) ,
20583	 => std_logic_vector(to_unsigned(183,8) ,
20584	 => std_logic_vector(to_unsigned(170,8) ,
20585	 => std_logic_vector(to_unsigned(170,8) ,
20586	 => std_logic_vector(to_unsigned(173,8) ,
20587	 => std_logic_vector(to_unsigned(170,8) ,
20588	 => std_logic_vector(to_unsigned(173,8) ,
20589	 => std_logic_vector(to_unsigned(175,8) ,
20590	 => std_logic_vector(to_unsigned(173,8) ,
20591	 => std_logic_vector(to_unsigned(175,8) ,
20592	 => std_logic_vector(to_unsigned(173,8) ,
20593	 => std_logic_vector(to_unsigned(170,8) ,
20594	 => std_logic_vector(to_unsigned(168,8) ,
20595	 => std_logic_vector(to_unsigned(171,8) ,
20596	 => std_logic_vector(to_unsigned(170,8) ,
20597	 => std_logic_vector(to_unsigned(164,8) ,
20598	 => std_logic_vector(to_unsigned(151,8) ,
20599	 => std_logic_vector(to_unsigned(127,8) ,
20600	 => std_logic_vector(to_unsigned(139,8) ,
20601	 => std_logic_vector(to_unsigned(109,8) ,
20602	 => std_logic_vector(to_unsigned(109,8) ,
20603	 => std_logic_vector(to_unsigned(133,8) ,
20604	 => std_logic_vector(to_unsigned(146,8) ,
20605	 => std_logic_vector(to_unsigned(154,8) ,
20606	 => std_logic_vector(to_unsigned(151,8) ,
20607	 => std_logic_vector(to_unsigned(142,8) ,
20608	 => std_logic_vector(to_unsigned(157,8) ,
20609	 => std_logic_vector(to_unsigned(156,8) ,
20610	 => std_logic_vector(to_unsigned(130,8) ,
20611	 => std_logic_vector(to_unsigned(125,8) ,
20612	 => std_logic_vector(to_unsigned(134,8) ,
20613	 => std_logic_vector(to_unsigned(142,8) ,
20614	 => std_logic_vector(to_unsigned(147,8) ,
20615	 => std_logic_vector(to_unsigned(144,8) ,
20616	 => std_logic_vector(to_unsigned(144,8) ,
20617	 => std_logic_vector(to_unsigned(138,8) ,
20618	 => std_logic_vector(to_unsigned(134,8) ,
20619	 => std_logic_vector(to_unsigned(125,8) ,
20620	 => std_logic_vector(to_unsigned(121,8) ,
20621	 => std_logic_vector(to_unsigned(112,8) ,
20622	 => std_logic_vector(to_unsigned(124,8) ,
20623	 => std_logic_vector(to_unsigned(128,8) ,
20624	 => std_logic_vector(to_unsigned(104,8) ,
20625	 => std_logic_vector(to_unsigned(104,8) ,
20626	 => std_logic_vector(to_unsigned(99,8) ,
20627	 => std_logic_vector(to_unsigned(90,8) ,
20628	 => std_logic_vector(to_unsigned(77,8) ,
20629	 => std_logic_vector(to_unsigned(91,8) ,
20630	 => std_logic_vector(to_unsigned(103,8) ,
20631	 => std_logic_vector(to_unsigned(100,8) ,
20632	 => std_logic_vector(to_unsigned(71,8) ,
20633	 => std_logic_vector(to_unsigned(74,8) ,
20634	 => std_logic_vector(to_unsigned(156,8) ,
20635	 => std_logic_vector(to_unsigned(157,8) ,
20636	 => std_logic_vector(to_unsigned(154,8) ,
20637	 => std_logic_vector(to_unsigned(156,8) ,
20638	 => std_logic_vector(to_unsigned(151,8) ,
20639	 => std_logic_vector(to_unsigned(118,8) ,
20640	 => std_logic_vector(to_unsigned(112,8) ,
20641	 => std_logic_vector(to_unsigned(115,8) ,
20642	 => std_logic_vector(to_unsigned(124,8) ,
20643	 => std_logic_vector(to_unsigned(156,8) ,
20644	 => std_logic_vector(to_unsigned(57,8) ,
20645	 => std_logic_vector(to_unsigned(1,8) ,
20646	 => std_logic_vector(to_unsigned(2,8) ,
20647	 => std_logic_vector(to_unsigned(6,8) ,
20648	 => std_logic_vector(to_unsigned(16,8) ,
20649	 => std_logic_vector(to_unsigned(8,8) ,
20650	 => std_logic_vector(to_unsigned(2,8) ,
20651	 => std_logic_vector(to_unsigned(2,8) ,
20652	 => std_logic_vector(to_unsigned(3,8) ,
20653	 => std_logic_vector(to_unsigned(5,8) ,
20654	 => std_logic_vector(to_unsigned(5,8) ,
20655	 => std_logic_vector(to_unsigned(1,8) ,
20656	 => std_logic_vector(to_unsigned(45,8) ,
20657	 => std_logic_vector(to_unsigned(170,8) ,
20658	 => std_logic_vector(to_unsigned(154,8) ,
20659	 => std_logic_vector(to_unsigned(147,8) ,
20660	 => std_logic_vector(to_unsigned(142,8) ,
20661	 => std_logic_vector(to_unsigned(146,8) ,
20662	 => std_logic_vector(to_unsigned(108,8) ,
20663	 => std_logic_vector(to_unsigned(96,8) ,
20664	 => std_logic_vector(to_unsigned(96,8) ,
20665	 => std_logic_vector(to_unsigned(86,8) ,
20666	 => std_logic_vector(to_unsigned(87,8) ,
20667	 => std_logic_vector(to_unsigned(90,8) ,
20668	 => std_logic_vector(to_unsigned(80,8) ,
20669	 => std_logic_vector(to_unsigned(77,8) ,
20670	 => std_logic_vector(to_unsigned(82,8) ,
20671	 => std_logic_vector(to_unsigned(87,8) ,
20672	 => std_logic_vector(to_unsigned(85,8) ,
20673	 => std_logic_vector(to_unsigned(78,8) ,
20674	 => std_logic_vector(to_unsigned(86,8) ,
20675	 => std_logic_vector(to_unsigned(88,8) ,
20676	 => std_logic_vector(to_unsigned(32,8) ,
20677	 => std_logic_vector(to_unsigned(5,8) ,
20678	 => std_logic_vector(to_unsigned(3,8) ,
20679	 => std_logic_vector(to_unsigned(2,8) ,
20680	 => std_logic_vector(to_unsigned(2,8) ,
20681	 => std_logic_vector(to_unsigned(4,8) ,
20682	 => std_logic_vector(to_unsigned(31,8) ,
20683	 => std_logic_vector(to_unsigned(99,8) ,
20684	 => std_logic_vector(to_unsigned(91,8) ,
20685	 => std_logic_vector(to_unsigned(93,8) ,
20686	 => std_logic_vector(to_unsigned(97,8) ,
20687	 => std_logic_vector(to_unsigned(95,8) ,
20688	 => std_logic_vector(to_unsigned(92,8) ,
20689	 => std_logic_vector(to_unsigned(90,8) ,
20690	 => std_logic_vector(to_unsigned(84,8) ,
20691	 => std_logic_vector(to_unsigned(84,8) ,
20692	 => std_logic_vector(to_unsigned(85,8) ,
20693	 => std_logic_vector(to_unsigned(79,8) ,
20694	 => std_logic_vector(to_unsigned(70,8) ,
20695	 => std_logic_vector(to_unsigned(79,8) ,
20696	 => std_logic_vector(to_unsigned(82,8) ,
20697	 => std_logic_vector(to_unsigned(86,8) ,
20698	 => std_logic_vector(to_unsigned(82,8) ,
20699	 => std_logic_vector(to_unsigned(84,8) ,
20700	 => std_logic_vector(to_unsigned(92,8) ,
20701	 => std_logic_vector(to_unsigned(99,8) ,
20702	 => std_logic_vector(to_unsigned(114,8) ,
20703	 => std_logic_vector(to_unsigned(77,8) ,
20704	 => std_logic_vector(to_unsigned(7,8) ,
20705	 => std_logic_vector(to_unsigned(3,8) ,
20706	 => std_logic_vector(to_unsigned(8,8) ,
20707	 => std_logic_vector(to_unsigned(19,8) ,
20708	 => std_logic_vector(to_unsigned(33,8) ,
20709	 => std_logic_vector(to_unsigned(34,8) ,
20710	 => std_logic_vector(to_unsigned(27,8) ,
20711	 => std_logic_vector(to_unsigned(35,8) ,
20712	 => std_logic_vector(to_unsigned(55,8) ,
20713	 => std_logic_vector(to_unsigned(43,8) ,
20714	 => std_logic_vector(to_unsigned(24,8) ,
20715	 => std_logic_vector(to_unsigned(65,8) ,
20716	 => std_logic_vector(to_unsigned(109,8) ,
20717	 => std_logic_vector(to_unsigned(99,8) ,
20718	 => std_logic_vector(to_unsigned(101,8) ,
20719	 => std_logic_vector(to_unsigned(111,8) ,
20720	 => std_logic_vector(to_unsigned(95,8) ,
20721	 => std_logic_vector(to_unsigned(97,8) ,
20722	 => std_logic_vector(to_unsigned(116,8) ,
20723	 => std_logic_vector(to_unsigned(103,8) ,
20724	 => std_logic_vector(to_unsigned(88,8) ,
20725	 => std_logic_vector(to_unsigned(111,8) ,
20726	 => std_logic_vector(to_unsigned(107,8) ,
20727	 => std_logic_vector(to_unsigned(86,8) ,
20728	 => std_logic_vector(to_unsigned(90,8) ,
20729	 => std_logic_vector(to_unsigned(81,8) ,
20730	 => std_logic_vector(to_unsigned(91,8) ,
20731	 => std_logic_vector(to_unsigned(54,8) ,
20732	 => std_logic_vector(to_unsigned(1,8) ,
20733	 => std_logic_vector(to_unsigned(0,8) ,
20734	 => std_logic_vector(to_unsigned(4,8) ,
20735	 => std_logic_vector(to_unsigned(78,8) ,
20736	 => std_logic_vector(to_unsigned(93,8) ,
20737	 => std_logic_vector(to_unsigned(105,8) ,
20738	 => std_logic_vector(to_unsigned(121,8) ,
20739	 => std_logic_vector(to_unsigned(108,8) ,
20740	 => std_logic_vector(to_unsigned(99,8) ,
20741	 => std_logic_vector(to_unsigned(105,8) ,
20742	 => std_logic_vector(to_unsigned(108,8) ,
20743	 => std_logic_vector(to_unsigned(111,8) ,
20744	 => std_logic_vector(to_unsigned(119,8) ,
20745	 => std_logic_vector(to_unsigned(125,8) ,
20746	 => std_logic_vector(to_unsigned(111,8) ,
20747	 => std_logic_vector(to_unsigned(97,8) ,
20748	 => std_logic_vector(to_unsigned(97,8) ,
20749	 => std_logic_vector(to_unsigned(95,8) ,
20750	 => std_logic_vector(to_unsigned(92,8) ,
20751	 => std_logic_vector(to_unsigned(97,8) ,
20752	 => std_logic_vector(to_unsigned(103,8) ,
20753	 => std_logic_vector(to_unsigned(22,8) ,
20754	 => std_logic_vector(to_unsigned(0,8) ,
20755	 => std_logic_vector(to_unsigned(1,8) ,
20756	 => std_logic_vector(to_unsigned(1,8) ,
20757	 => std_logic_vector(to_unsigned(0,8) ,
20758	 => std_logic_vector(to_unsigned(0,8) ,
20759	 => std_logic_vector(to_unsigned(1,8) ,
20760	 => std_logic_vector(to_unsigned(3,8) ,
20761	 => std_logic_vector(to_unsigned(6,8) ,
20762	 => std_logic_vector(to_unsigned(3,8) ,
20763	 => std_logic_vector(to_unsigned(2,8) ,
20764	 => std_logic_vector(to_unsigned(1,8) ,
20765	 => std_logic_vector(to_unsigned(1,8) ,
20766	 => std_logic_vector(to_unsigned(1,8) ,
20767	 => std_logic_vector(to_unsigned(0,8) ,
20768	 => std_logic_vector(to_unsigned(3,8) ,
20769	 => std_logic_vector(to_unsigned(84,8) ,
20770	 => std_logic_vector(to_unsigned(108,8) ,
20771	 => std_logic_vector(to_unsigned(90,8) ,
20772	 => std_logic_vector(to_unsigned(95,8) ,
20773	 => std_logic_vector(to_unsigned(95,8) ,
20774	 => std_logic_vector(to_unsigned(95,8) ,
20775	 => std_logic_vector(to_unsigned(99,8) ,
20776	 => std_logic_vector(to_unsigned(90,8) ,
20777	 => std_logic_vector(to_unsigned(87,8) ,
20778	 => std_logic_vector(to_unsigned(93,8) ,
20779	 => std_logic_vector(to_unsigned(93,8) ,
20780	 => std_logic_vector(to_unsigned(112,8) ,
20781	 => std_logic_vector(to_unsigned(156,8) ,
20782	 => std_logic_vector(to_unsigned(166,8) ,
20783	 => std_logic_vector(to_unsigned(168,8) ,
20784	 => std_logic_vector(to_unsigned(161,8) ,
20785	 => std_logic_vector(to_unsigned(138,8) ,
20786	 => std_logic_vector(to_unsigned(136,8) ,
20787	 => std_logic_vector(to_unsigned(131,8) ,
20788	 => std_logic_vector(to_unsigned(112,8) ,
20789	 => std_logic_vector(to_unsigned(111,8) ,
20790	 => std_logic_vector(to_unsigned(97,8) ,
20791	 => std_logic_vector(to_unsigned(92,8) ,
20792	 => std_logic_vector(to_unsigned(99,8) ,
20793	 => std_logic_vector(to_unsigned(103,8) ,
20794	 => std_logic_vector(to_unsigned(86,8) ,
20795	 => std_logic_vector(to_unsigned(78,8) ,
20796	 => std_logic_vector(to_unsigned(95,8) ,
20797	 => std_logic_vector(to_unsigned(105,8) ,
20798	 => std_logic_vector(to_unsigned(105,8) ,
20799	 => std_logic_vector(to_unsigned(92,8) ,
20800	 => std_logic_vector(to_unsigned(81,8) ,
20801	 => std_logic_vector(to_unsigned(141,8) ,
20802	 => std_logic_vector(to_unsigned(134,8) ,
20803	 => std_logic_vector(to_unsigned(138,8) ,
20804	 => std_logic_vector(to_unsigned(152,8) ,
20805	 => std_logic_vector(to_unsigned(163,8) ,
20806	 => std_logic_vector(to_unsigned(157,8) ,
20807	 => std_logic_vector(to_unsigned(159,8) ,
20808	 => std_logic_vector(to_unsigned(161,8) ,
20809	 => std_logic_vector(to_unsigned(163,8) ,
20810	 => std_logic_vector(to_unsigned(164,8) ,
20811	 => std_logic_vector(to_unsigned(166,8) ,
20812	 => std_logic_vector(to_unsigned(146,8) ,
20813	 => std_logic_vector(to_unsigned(78,8) ,
20814	 => std_logic_vector(to_unsigned(24,8) ,
20815	 => std_logic_vector(to_unsigned(2,8) ,
20816	 => std_logic_vector(to_unsigned(11,8) ,
20817	 => std_logic_vector(to_unsigned(26,8) ,
20818	 => std_logic_vector(to_unsigned(27,8) ,
20819	 => std_logic_vector(to_unsigned(18,8) ,
20820	 => std_logic_vector(to_unsigned(19,8) ,
20821	 => std_logic_vector(to_unsigned(15,8) ,
20822	 => std_logic_vector(to_unsigned(5,8) ,
20823	 => std_logic_vector(to_unsigned(6,8) ,
20824	 => std_logic_vector(to_unsigned(1,8) ,
20825	 => std_logic_vector(to_unsigned(37,8) ,
20826	 => std_logic_vector(to_unsigned(116,8) ,
20827	 => std_logic_vector(to_unsigned(25,8) ,
20828	 => std_logic_vector(to_unsigned(8,8) ,
20829	 => std_logic_vector(to_unsigned(20,8) ,
20830	 => std_logic_vector(to_unsigned(44,8) ,
20831	 => std_logic_vector(to_unsigned(52,8) ,
20832	 => std_logic_vector(to_unsigned(19,8) ,
20833	 => std_logic_vector(to_unsigned(15,8) ,
20834	 => std_logic_vector(to_unsigned(22,8) ,
20835	 => std_logic_vector(to_unsigned(11,8) ,
20836	 => std_logic_vector(to_unsigned(20,8) ,
20837	 => std_logic_vector(to_unsigned(41,8) ,
20838	 => std_logic_vector(to_unsigned(37,8) ,
20839	 => std_logic_vector(to_unsigned(27,8) ,
20840	 => std_logic_vector(to_unsigned(67,8) ,
20841	 => std_logic_vector(to_unsigned(51,8) ,
20842	 => std_logic_vector(to_unsigned(59,8) ,
20843	 => std_logic_vector(to_unsigned(124,8) ,
20844	 => std_logic_vector(to_unsigned(154,8) ,
20845	 => std_logic_vector(to_unsigned(164,8) ,
20846	 => std_logic_vector(to_unsigned(171,8) ,
20847	 => std_logic_vector(to_unsigned(168,8) ,
20848	 => std_logic_vector(to_unsigned(164,8) ,
20849	 => std_logic_vector(to_unsigned(161,8) ,
20850	 => std_logic_vector(to_unsigned(159,8) ,
20851	 => std_logic_vector(to_unsigned(168,8) ,
20852	 => std_logic_vector(to_unsigned(166,8) ,
20853	 => std_logic_vector(to_unsigned(164,8) ,
20854	 => std_logic_vector(to_unsigned(164,8) ,
20855	 => std_logic_vector(to_unsigned(154,8) ,
20856	 => std_logic_vector(to_unsigned(166,8) ,
20857	 => std_logic_vector(to_unsigned(147,8) ,
20858	 => std_logic_vector(to_unsigned(12,8) ,
20859	 => std_logic_vector(to_unsigned(2,8) ,
20860	 => std_logic_vector(to_unsigned(6,8) ,
20861	 => std_logic_vector(to_unsigned(6,8) ,
20862	 => std_logic_vector(to_unsigned(7,8) ,
20863	 => std_logic_vector(to_unsigned(6,8) ,
20864	 => std_logic_vector(to_unsigned(3,8) ,
20865	 => std_logic_vector(to_unsigned(5,8) ,
20866	 => std_logic_vector(to_unsigned(5,8) ,
20867	 => std_logic_vector(to_unsigned(47,8) ,
20868	 => std_logic_vector(to_unsigned(214,8) ,
20869	 => std_logic_vector(to_unsigned(22,8) ,
20870	 => std_logic_vector(to_unsigned(14,8) ,
20871	 => std_logic_vector(to_unsigned(154,8) ,
20872	 => std_logic_vector(to_unsigned(166,8) ,
20873	 => std_logic_vector(to_unsigned(159,8) ,
20874	 => std_logic_vector(to_unsigned(168,8) ,
20875	 => std_logic_vector(to_unsigned(157,8) ,
20876	 => std_logic_vector(to_unsigned(147,8) ,
20877	 => std_logic_vector(to_unsigned(171,8) ,
20878	 => std_logic_vector(to_unsigned(170,8) ,
20879	 => std_logic_vector(to_unsigned(166,8) ,
20880	 => std_logic_vector(to_unsigned(166,8) ,
20881	 => std_logic_vector(to_unsigned(164,8) ,
20882	 => std_logic_vector(to_unsigned(164,8) ,
20883	 => std_logic_vector(to_unsigned(164,8) ,
20884	 => std_logic_vector(to_unsigned(166,8) ,
20885	 => std_logic_vector(to_unsigned(166,8) ,
20886	 => std_logic_vector(to_unsigned(164,8) ,
20887	 => std_logic_vector(to_unsigned(163,8) ,
20888	 => std_logic_vector(to_unsigned(161,8) ,
20889	 => std_logic_vector(to_unsigned(156,8) ,
20890	 => std_logic_vector(to_unsigned(173,8) ,
20891	 => std_logic_vector(to_unsigned(87,8) ,
20892	 => std_logic_vector(to_unsigned(3,8) ,
20893	 => std_logic_vector(to_unsigned(3,8) ,
20894	 => std_logic_vector(to_unsigned(4,8) ,
20895	 => std_logic_vector(to_unsigned(3,8) ,
20896	 => std_logic_vector(to_unsigned(2,8) ,
20897	 => std_logic_vector(to_unsigned(3,8) ,
20898	 => std_logic_vector(to_unsigned(7,8) ,
20899	 => std_logic_vector(to_unsigned(10,8) ,
20900	 => std_logic_vector(to_unsigned(17,8) ,
20901	 => std_logic_vector(to_unsigned(62,8) ,
20902	 => std_logic_vector(to_unsigned(159,8) ,
20903	 => std_logic_vector(to_unsigned(179,8) ,
20904	 => std_logic_vector(to_unsigned(170,8) ,
20905	 => std_logic_vector(to_unsigned(168,8) ,
20906	 => std_logic_vector(to_unsigned(171,8) ,
20907	 => std_logic_vector(to_unsigned(171,8) ,
20908	 => std_logic_vector(to_unsigned(171,8) ,
20909	 => std_logic_vector(to_unsigned(173,8) ,
20910	 => std_logic_vector(to_unsigned(171,8) ,
20911	 => std_logic_vector(to_unsigned(168,8) ,
20912	 => std_logic_vector(to_unsigned(168,8) ,
20913	 => std_logic_vector(to_unsigned(168,8) ,
20914	 => std_logic_vector(to_unsigned(168,8) ,
20915	 => std_logic_vector(to_unsigned(168,8) ,
20916	 => std_logic_vector(to_unsigned(164,8) ,
20917	 => std_logic_vector(to_unsigned(157,8) ,
20918	 => std_logic_vector(to_unsigned(161,8) ,
20919	 => std_logic_vector(to_unsigned(161,8) ,
20920	 => std_logic_vector(to_unsigned(152,8) ,
20921	 => std_logic_vector(to_unsigned(119,8) ,
20922	 => std_logic_vector(to_unsigned(73,8) ,
20923	 => std_logic_vector(to_unsigned(46,8) ,
20924	 => std_logic_vector(to_unsigned(103,8) ,
20925	 => std_logic_vector(to_unsigned(131,8) ,
20926	 => std_logic_vector(to_unsigned(96,8) ,
20927	 => std_logic_vector(to_unsigned(80,8) ,
20928	 => std_logic_vector(to_unsigned(131,8) ,
20929	 => std_logic_vector(to_unsigned(166,8) ,
20930	 => std_logic_vector(to_unsigned(136,8) ,
20931	 => std_logic_vector(to_unsigned(125,8) ,
20932	 => std_logic_vector(to_unsigned(131,8) ,
20933	 => std_logic_vector(to_unsigned(142,8) ,
20934	 => std_logic_vector(to_unsigned(151,8) ,
20935	 => std_logic_vector(to_unsigned(142,8) ,
20936	 => std_logic_vector(to_unsigned(136,8) ,
20937	 => std_logic_vector(to_unsigned(139,8) ,
20938	 => std_logic_vector(to_unsigned(138,8) ,
20939	 => std_logic_vector(to_unsigned(128,8) ,
20940	 => std_logic_vector(to_unsigned(114,8) ,
20941	 => std_logic_vector(to_unsigned(119,8) ,
20942	 => std_logic_vector(to_unsigned(131,8) ,
20943	 => std_logic_vector(to_unsigned(118,8) ,
20944	 => std_logic_vector(to_unsigned(91,8) ,
20945	 => std_logic_vector(to_unsigned(90,8) ,
20946	 => std_logic_vector(to_unsigned(90,8) ,
20947	 => std_logic_vector(to_unsigned(90,8) ,
20948	 => std_logic_vector(to_unsigned(85,8) ,
20949	 => std_logic_vector(to_unsigned(70,8) ,
20950	 => std_logic_vector(to_unsigned(80,8) ,
20951	 => std_logic_vector(to_unsigned(77,8) ,
20952	 => std_logic_vector(to_unsigned(36,8) ,
20953	 => std_logic_vector(to_unsigned(45,8) ,
20954	 => std_logic_vector(to_unsigned(146,8) ,
20955	 => std_logic_vector(to_unsigned(157,8) ,
20956	 => std_logic_vector(to_unsigned(156,8) ,
20957	 => std_logic_vector(to_unsigned(157,8) ,
20958	 => std_logic_vector(to_unsigned(152,8) ,
20959	 => std_logic_vector(to_unsigned(125,8) ,
20960	 => std_logic_vector(to_unsigned(124,8) ,
20961	 => std_logic_vector(to_unsigned(127,8) ,
20962	 => std_logic_vector(to_unsigned(115,8) ,
20963	 => std_logic_vector(to_unsigned(138,8) ,
20964	 => std_logic_vector(to_unsigned(52,8) ,
20965	 => std_logic_vector(to_unsigned(2,8) ,
20966	 => std_logic_vector(to_unsigned(3,8) ,
20967	 => std_logic_vector(to_unsigned(11,8) ,
20968	 => std_logic_vector(to_unsigned(29,8) ,
20969	 => std_logic_vector(to_unsigned(26,8) ,
20970	 => std_logic_vector(to_unsigned(13,8) ,
20971	 => std_logic_vector(to_unsigned(5,8) ,
20972	 => std_logic_vector(to_unsigned(3,8) ,
20973	 => std_logic_vector(to_unsigned(3,8) ,
20974	 => std_logic_vector(to_unsigned(2,8) ,
20975	 => std_logic_vector(to_unsigned(3,8) ,
20976	 => std_logic_vector(to_unsigned(76,8) ,
20977	 => std_logic_vector(to_unsigned(173,8) ,
20978	 => std_logic_vector(to_unsigned(151,8) ,
20979	 => std_logic_vector(to_unsigned(152,8) ,
20980	 => std_logic_vector(to_unsigned(151,8) ,
20981	 => std_logic_vector(to_unsigned(141,8) ,
20982	 => std_logic_vector(to_unsigned(104,8) ,
20983	 => std_logic_vector(to_unsigned(90,8) ,
20984	 => std_logic_vector(to_unsigned(103,8) ,
20985	 => std_logic_vector(to_unsigned(88,8) ,
20986	 => std_logic_vector(to_unsigned(86,8) ,
20987	 => std_logic_vector(to_unsigned(92,8) ,
20988	 => std_logic_vector(to_unsigned(85,8) ,
20989	 => std_logic_vector(to_unsigned(78,8) ,
20990	 => std_logic_vector(to_unsigned(84,8) ,
20991	 => std_logic_vector(to_unsigned(86,8) ,
20992	 => std_logic_vector(to_unsigned(77,8) ,
20993	 => std_logic_vector(to_unsigned(86,8) ,
20994	 => std_logic_vector(to_unsigned(73,8) ,
20995	 => std_logic_vector(to_unsigned(14,8) ,
20996	 => std_logic_vector(to_unsigned(1,8) ,
20997	 => std_logic_vector(to_unsigned(0,8) ,
20998	 => std_logic_vector(to_unsigned(0,8) ,
20999	 => std_logic_vector(to_unsigned(0,8) ,
21000	 => std_logic_vector(to_unsigned(1,8) ,
21001	 => std_logic_vector(to_unsigned(0,8) ,
21002	 => std_logic_vector(to_unsigned(2,8) ,
21003	 => std_logic_vector(to_unsigned(60,8) ,
21004	 => std_logic_vector(to_unsigned(109,8) ,
21005	 => std_logic_vector(to_unsigned(96,8) ,
21006	 => std_logic_vector(to_unsigned(111,8) ,
21007	 => std_logic_vector(to_unsigned(105,8) ,
21008	 => std_logic_vector(to_unsigned(88,8) ,
21009	 => std_logic_vector(to_unsigned(77,8) ,
21010	 => std_logic_vector(to_unsigned(82,8) ,
21011	 => std_logic_vector(to_unsigned(80,8) ,
21012	 => std_logic_vector(to_unsigned(81,8) ,
21013	 => std_logic_vector(to_unsigned(84,8) ,
21014	 => std_logic_vector(to_unsigned(81,8) ,
21015	 => std_logic_vector(to_unsigned(90,8) ,
21016	 => std_logic_vector(to_unsigned(85,8) ,
21017	 => std_logic_vector(to_unsigned(91,8) ,
21018	 => std_logic_vector(to_unsigned(95,8) ,
21019	 => std_logic_vector(to_unsigned(88,8) ,
21020	 => std_logic_vector(to_unsigned(105,8) ,
21021	 => std_logic_vector(to_unsigned(79,8) ,
21022	 => std_logic_vector(to_unsigned(23,8) ,
21023	 => std_logic_vector(to_unsigned(17,8) ,
21024	 => std_logic_vector(to_unsigned(5,8) ,
21025	 => std_logic_vector(to_unsigned(2,8) ,
21026	 => std_logic_vector(to_unsigned(9,8) ,
21027	 => std_logic_vector(to_unsigned(20,8) ,
21028	 => std_logic_vector(to_unsigned(23,8) ,
21029	 => std_logic_vector(to_unsigned(23,8) ,
21030	 => std_logic_vector(to_unsigned(17,8) ,
21031	 => std_logic_vector(to_unsigned(20,8) ,
21032	 => std_logic_vector(to_unsigned(41,8) ,
21033	 => std_logic_vector(to_unsigned(49,8) ,
21034	 => std_logic_vector(to_unsigned(45,8) ,
21035	 => std_logic_vector(to_unsigned(69,8) ,
21036	 => std_logic_vector(to_unsigned(109,8) ,
21037	 => std_logic_vector(to_unsigned(109,8) ,
21038	 => std_logic_vector(to_unsigned(107,8) ,
21039	 => std_logic_vector(to_unsigned(114,8) ,
21040	 => std_logic_vector(to_unsigned(109,8) ,
21041	 => std_logic_vector(to_unsigned(105,8) ,
21042	 => std_logic_vector(to_unsigned(104,8) ,
21043	 => std_logic_vector(to_unsigned(99,8) ,
21044	 => std_logic_vector(to_unsigned(95,8) ,
21045	 => std_logic_vector(to_unsigned(96,8) ,
21046	 => std_logic_vector(to_unsigned(105,8) ,
21047	 => std_logic_vector(to_unsigned(99,8) ,
21048	 => std_logic_vector(to_unsigned(100,8) ,
21049	 => std_logic_vector(to_unsigned(95,8) ,
21050	 => std_logic_vector(to_unsigned(107,8) ,
21051	 => std_logic_vector(to_unsigned(91,8) ,
21052	 => std_logic_vector(to_unsigned(5,8) ,
21053	 => std_logic_vector(to_unsigned(0,8) ,
21054	 => std_logic_vector(to_unsigned(1,8) ,
21055	 => std_logic_vector(to_unsigned(57,8) ,
21056	 => std_logic_vector(to_unsigned(112,8) ,
21057	 => std_logic_vector(to_unsigned(104,8) ,
21058	 => std_logic_vector(to_unsigned(112,8) ,
21059	 => std_logic_vector(to_unsigned(111,8) ,
21060	 => std_logic_vector(to_unsigned(109,8) ,
21061	 => std_logic_vector(to_unsigned(116,8) ,
21062	 => std_logic_vector(to_unsigned(122,8) ,
21063	 => std_logic_vector(to_unsigned(119,8) ,
21064	 => std_logic_vector(to_unsigned(122,8) ,
21065	 => std_logic_vector(to_unsigned(122,8) ,
21066	 => std_logic_vector(to_unsigned(118,8) ,
21067	 => std_logic_vector(to_unsigned(112,8) ,
21068	 => std_logic_vector(to_unsigned(101,8) ,
21069	 => std_logic_vector(to_unsigned(99,8) ,
21070	 => std_logic_vector(to_unsigned(101,8) ,
21071	 => std_logic_vector(to_unsigned(103,8) ,
21072	 => std_logic_vector(to_unsigned(86,8) ,
21073	 => std_logic_vector(to_unsigned(7,8) ,
21074	 => std_logic_vector(to_unsigned(0,8) ,
21075	 => std_logic_vector(to_unsigned(1,8) ,
21076	 => std_logic_vector(to_unsigned(0,8) ,
21077	 => std_logic_vector(to_unsigned(1,8) ,
21078	 => std_logic_vector(to_unsigned(2,8) ,
21079	 => std_logic_vector(to_unsigned(8,8) ,
21080	 => std_logic_vector(to_unsigned(13,8) ,
21081	 => std_logic_vector(to_unsigned(13,8) ,
21082	 => std_logic_vector(to_unsigned(6,8) ,
21083	 => std_logic_vector(to_unsigned(7,8) ,
21084	 => std_logic_vector(to_unsigned(8,8) ,
21085	 => std_logic_vector(to_unsigned(4,8) ,
21086	 => std_logic_vector(to_unsigned(3,8) ,
21087	 => std_logic_vector(to_unsigned(2,8) ,
21088	 => std_logic_vector(to_unsigned(22,8) ,
21089	 => std_logic_vector(to_unsigned(101,8) ,
21090	 => std_logic_vector(to_unsigned(100,8) ,
21091	 => std_logic_vector(to_unsigned(93,8) ,
21092	 => std_logic_vector(to_unsigned(91,8) ,
21093	 => std_logic_vector(to_unsigned(91,8) ,
21094	 => std_logic_vector(to_unsigned(95,8) ,
21095	 => std_logic_vector(to_unsigned(92,8) ,
21096	 => std_logic_vector(to_unsigned(91,8) ,
21097	 => std_logic_vector(to_unsigned(88,8) ,
21098	 => std_logic_vector(to_unsigned(90,8) ,
21099	 => std_logic_vector(to_unsigned(93,8) ,
21100	 => std_logic_vector(to_unsigned(85,8) ,
21101	 => std_logic_vector(to_unsigned(133,8) ,
21102	 => std_logic_vector(to_unsigned(170,8) ,
21103	 => std_logic_vector(to_unsigned(163,8) ,
21104	 => std_logic_vector(to_unsigned(152,8) ,
21105	 => std_logic_vector(to_unsigned(149,8) ,
21106	 => std_logic_vector(to_unsigned(146,8) ,
21107	 => std_logic_vector(to_unsigned(142,8) ,
21108	 => std_logic_vector(to_unsigned(134,8) ,
21109	 => std_logic_vector(to_unsigned(122,8) ,
21110	 => std_logic_vector(to_unsigned(105,8) ,
21111	 => std_logic_vector(to_unsigned(105,8) ,
21112	 => std_logic_vector(to_unsigned(105,8) ,
21113	 => std_logic_vector(to_unsigned(101,8) ,
21114	 => std_logic_vector(to_unsigned(86,8) ,
21115	 => std_logic_vector(to_unsigned(87,8) ,
21116	 => std_logic_vector(to_unsigned(115,8) ,
21117	 => std_logic_vector(to_unsigned(147,8) ,
21118	 => std_logic_vector(to_unsigned(134,8) ,
21119	 => std_logic_vector(to_unsigned(78,8) ,
21120	 => std_logic_vector(to_unsigned(69,8) ,
21121	 => std_logic_vector(to_unsigned(149,8) ,
21122	 => std_logic_vector(to_unsigned(141,8) ,
21123	 => std_logic_vector(to_unsigned(141,8) ,
21124	 => std_logic_vector(to_unsigned(149,8) ,
21125	 => std_logic_vector(to_unsigned(157,8) ,
21126	 => std_logic_vector(to_unsigned(161,8) ,
21127	 => std_logic_vector(to_unsigned(161,8) ,
21128	 => std_logic_vector(to_unsigned(166,8) ,
21129	 => std_logic_vector(to_unsigned(168,8) ,
21130	 => std_logic_vector(to_unsigned(163,8) ,
21131	 => std_logic_vector(to_unsigned(138,8) ,
21132	 => std_logic_vector(to_unsigned(105,8) ,
21133	 => std_logic_vector(to_unsigned(30,8) ,
21134	 => std_logic_vector(to_unsigned(2,8) ,
21135	 => std_logic_vector(to_unsigned(1,8) ,
21136	 => std_logic_vector(to_unsigned(3,8) ,
21137	 => std_logic_vector(to_unsigned(10,8) ,
21138	 => std_logic_vector(to_unsigned(18,8) ,
21139	 => std_logic_vector(to_unsigned(28,8) ,
21140	 => std_logic_vector(to_unsigned(27,8) ,
21141	 => std_logic_vector(to_unsigned(25,8) ,
21142	 => std_logic_vector(to_unsigned(10,8) ,
21143	 => std_logic_vector(to_unsigned(13,8) ,
21144	 => std_logic_vector(to_unsigned(13,8) ,
21145	 => std_logic_vector(to_unsigned(23,8) ,
21146	 => std_logic_vector(to_unsigned(38,8) ,
21147	 => std_logic_vector(to_unsigned(16,8) ,
21148	 => std_logic_vector(to_unsigned(4,8) ,
21149	 => std_logic_vector(to_unsigned(7,8) ,
21150	 => std_logic_vector(to_unsigned(34,8) ,
21151	 => std_logic_vector(to_unsigned(26,8) ,
21152	 => std_logic_vector(to_unsigned(17,8) ,
21153	 => std_logic_vector(to_unsigned(16,8) ,
21154	 => std_logic_vector(to_unsigned(16,8) ,
21155	 => std_logic_vector(to_unsigned(8,8) ,
21156	 => std_logic_vector(to_unsigned(15,8) ,
21157	 => std_logic_vector(to_unsigned(40,8) ,
21158	 => std_logic_vector(to_unsigned(41,8) ,
21159	 => std_logic_vector(to_unsigned(44,8) ,
21160	 => std_logic_vector(to_unsigned(37,8) ,
21161	 => std_logic_vector(to_unsigned(6,8) ,
21162	 => std_logic_vector(to_unsigned(2,8) ,
21163	 => std_logic_vector(to_unsigned(19,8) ,
21164	 => std_logic_vector(to_unsigned(97,8) ,
21165	 => std_logic_vector(to_unsigned(114,8) ,
21166	 => std_logic_vector(to_unsigned(130,8) ,
21167	 => std_logic_vector(to_unsigned(154,8) ,
21168	 => std_logic_vector(to_unsigned(168,8) ,
21169	 => std_logic_vector(to_unsigned(168,8) ,
21170	 => std_logic_vector(to_unsigned(161,8) ,
21171	 => std_logic_vector(to_unsigned(166,8) ,
21172	 => std_logic_vector(to_unsigned(164,8) ,
21173	 => std_logic_vector(to_unsigned(166,8) ,
21174	 => std_logic_vector(to_unsigned(161,8) ,
21175	 => std_logic_vector(to_unsigned(161,8) ,
21176	 => std_logic_vector(to_unsigned(177,8) ,
21177	 => std_logic_vector(to_unsigned(136,8) ,
21178	 => std_logic_vector(to_unsigned(8,8) ,
21179	 => std_logic_vector(to_unsigned(3,8) ,
21180	 => std_logic_vector(to_unsigned(6,8) ,
21181	 => std_logic_vector(to_unsigned(8,8) ,
21182	 => std_logic_vector(to_unsigned(10,8) ,
21183	 => std_logic_vector(to_unsigned(8,8) ,
21184	 => std_logic_vector(to_unsigned(9,8) ,
21185	 => std_logic_vector(to_unsigned(10,8) ,
21186	 => std_logic_vector(to_unsigned(12,8) ,
21187	 => std_logic_vector(to_unsigned(35,8) ,
21188	 => std_logic_vector(to_unsigned(127,8) ,
21189	 => std_logic_vector(to_unsigned(88,8) ,
21190	 => std_logic_vector(to_unsigned(28,8) ,
21191	 => std_logic_vector(to_unsigned(114,8) ,
21192	 => std_logic_vector(to_unsigned(166,8) ,
21193	 => std_logic_vector(to_unsigned(159,8) ,
21194	 => std_logic_vector(to_unsigned(161,8) ,
21195	 => std_logic_vector(to_unsigned(161,8) ,
21196	 => std_logic_vector(to_unsigned(168,8) ,
21197	 => std_logic_vector(to_unsigned(152,8) ,
21198	 => std_logic_vector(to_unsigned(166,8) ,
21199	 => std_logic_vector(to_unsigned(171,8) ,
21200	 => std_logic_vector(to_unsigned(164,8) ,
21201	 => std_logic_vector(to_unsigned(164,8) ,
21202	 => std_logic_vector(to_unsigned(166,8) ,
21203	 => std_logic_vector(to_unsigned(163,8) ,
21204	 => std_logic_vector(to_unsigned(164,8) ,
21205	 => std_logic_vector(to_unsigned(164,8) ,
21206	 => std_logic_vector(to_unsigned(164,8) ,
21207	 => std_logic_vector(to_unsigned(166,8) ,
21208	 => std_logic_vector(to_unsigned(163,8) ,
21209	 => std_logic_vector(to_unsigned(156,8) ,
21210	 => std_logic_vector(to_unsigned(161,8) ,
21211	 => std_logic_vector(to_unsigned(161,8) ,
21212	 => std_logic_vector(to_unsigned(32,8) ,
21213	 => std_logic_vector(to_unsigned(2,8) ,
21214	 => std_logic_vector(to_unsigned(2,8) ,
21215	 => std_logic_vector(to_unsigned(2,8) ,
21216	 => std_logic_vector(to_unsigned(2,8) ,
21217	 => std_logic_vector(to_unsigned(4,8) ,
21218	 => std_logic_vector(to_unsigned(10,8) ,
21219	 => std_logic_vector(to_unsigned(17,8) ,
21220	 => std_logic_vector(to_unsigned(29,8) ,
21221	 => std_logic_vector(to_unsigned(115,8) ,
21222	 => std_logic_vector(to_unsigned(177,8) ,
21223	 => std_logic_vector(to_unsigned(170,8) ,
21224	 => std_logic_vector(to_unsigned(166,8) ,
21225	 => std_logic_vector(to_unsigned(168,8) ,
21226	 => std_logic_vector(to_unsigned(163,8) ,
21227	 => std_logic_vector(to_unsigned(171,8) ,
21228	 => std_logic_vector(to_unsigned(170,8) ,
21229	 => std_logic_vector(to_unsigned(168,8) ,
21230	 => std_logic_vector(to_unsigned(166,8) ,
21231	 => std_logic_vector(to_unsigned(166,8) ,
21232	 => std_logic_vector(to_unsigned(166,8) ,
21233	 => std_logic_vector(to_unsigned(164,8) ,
21234	 => std_logic_vector(to_unsigned(168,8) ,
21235	 => std_logic_vector(to_unsigned(166,8) ,
21236	 => std_logic_vector(to_unsigned(163,8) ,
21237	 => std_logic_vector(to_unsigned(159,8) ,
21238	 => std_logic_vector(to_unsigned(149,8) ,
21239	 => std_logic_vector(to_unsigned(161,8) ,
21240	 => std_logic_vector(to_unsigned(125,8) ,
21241	 => std_logic_vector(to_unsigned(96,8) ,
21242	 => std_logic_vector(to_unsigned(45,8) ,
21243	 => std_logic_vector(to_unsigned(23,8) ,
21244	 => std_logic_vector(to_unsigned(63,8) ,
21245	 => std_logic_vector(to_unsigned(101,8) ,
21246	 => std_logic_vector(to_unsigned(65,8) ,
21247	 => std_logic_vector(to_unsigned(32,8) ,
21248	 => std_logic_vector(to_unsigned(90,8) ,
21249	 => std_logic_vector(to_unsigned(170,8) ,
21250	 => std_logic_vector(to_unsigned(133,8) ,
21251	 => std_logic_vector(to_unsigned(124,8) ,
21252	 => std_logic_vector(to_unsigned(138,8) ,
21253	 => std_logic_vector(to_unsigned(146,8) ,
21254	 => std_logic_vector(to_unsigned(147,8) ,
21255	 => std_logic_vector(to_unsigned(146,8) ,
21256	 => std_logic_vector(to_unsigned(139,8) ,
21257	 => std_logic_vector(to_unsigned(139,8) ,
21258	 => std_logic_vector(to_unsigned(139,8) ,
21259	 => std_logic_vector(to_unsigned(125,8) ,
21260	 => std_logic_vector(to_unsigned(121,8) ,
21261	 => std_logic_vector(to_unsigned(131,8) ,
21262	 => std_logic_vector(to_unsigned(134,8) ,
21263	 => std_logic_vector(to_unsigned(107,8) ,
21264	 => std_logic_vector(to_unsigned(47,8) ,
21265	 => std_logic_vector(to_unsigned(54,8) ,
21266	 => std_logic_vector(to_unsigned(95,8) ,
21267	 => std_logic_vector(to_unsigned(114,8) ,
21268	 => std_logic_vector(to_unsigned(118,8) ,
21269	 => std_logic_vector(to_unsigned(79,8) ,
21270	 => std_logic_vector(to_unsigned(60,8) ,
21271	 => std_logic_vector(to_unsigned(92,8) ,
21272	 => std_logic_vector(to_unsigned(59,8) ,
21273	 => std_logic_vector(to_unsigned(34,8) ,
21274	 => std_logic_vector(to_unsigned(124,8) ,
21275	 => std_logic_vector(to_unsigned(173,8) ,
21276	 => std_logic_vector(to_unsigned(152,8) ,
21277	 => std_logic_vector(to_unsigned(157,8) ,
21278	 => std_logic_vector(to_unsigned(154,8) ,
21279	 => std_logic_vector(to_unsigned(138,8) ,
21280	 => std_logic_vector(to_unsigned(133,8) ,
21281	 => std_logic_vector(to_unsigned(124,8) ,
21282	 => std_logic_vector(to_unsigned(104,8) ,
21283	 => std_logic_vector(to_unsigned(104,8) ,
21284	 => std_logic_vector(to_unsigned(88,8) ,
21285	 => std_logic_vector(to_unsigned(17,8) ,
21286	 => std_logic_vector(to_unsigned(1,8) ,
21287	 => std_logic_vector(to_unsigned(0,8) ,
21288	 => std_logic_vector(to_unsigned(2,8) ,
21289	 => std_logic_vector(to_unsigned(12,8) ,
21290	 => std_logic_vector(to_unsigned(26,8) ,
21291	 => std_logic_vector(to_unsigned(12,8) ,
21292	 => std_logic_vector(to_unsigned(7,8) ,
21293	 => std_logic_vector(to_unsigned(8,8) ,
21294	 => std_logic_vector(to_unsigned(4,8) ,
21295	 => std_logic_vector(to_unsigned(13,8) ,
21296	 => std_logic_vector(to_unsigned(130,8) ,
21297	 => std_logic_vector(to_unsigned(168,8) ,
21298	 => std_logic_vector(to_unsigned(146,8) ,
21299	 => std_logic_vector(to_unsigned(154,8) ,
21300	 => std_logic_vector(to_unsigned(151,8) ,
21301	 => std_logic_vector(to_unsigned(141,8) ,
21302	 => std_logic_vector(to_unsigned(118,8) ,
21303	 => std_logic_vector(to_unsigned(114,8) ,
21304	 => std_logic_vector(to_unsigned(114,8) ,
21305	 => std_logic_vector(to_unsigned(91,8) ,
21306	 => std_logic_vector(to_unsigned(90,8) ,
21307	 => std_logic_vector(to_unsigned(95,8) ,
21308	 => std_logic_vector(to_unsigned(86,8) ,
21309	 => std_logic_vector(to_unsigned(85,8) ,
21310	 => std_logic_vector(to_unsigned(91,8) ,
21311	 => std_logic_vector(to_unsigned(99,8) ,
21312	 => std_logic_vector(to_unsigned(90,8) ,
21313	 => std_logic_vector(to_unsigned(73,8) ,
21314	 => std_logic_vector(to_unsigned(11,8) ,
21315	 => std_logic_vector(to_unsigned(0,8) ,
21316	 => std_logic_vector(to_unsigned(1,8) ,
21317	 => std_logic_vector(to_unsigned(1,8) ,
21318	 => std_logic_vector(to_unsigned(1,8) ,
21319	 => std_logic_vector(to_unsigned(1,8) ,
21320	 => std_logic_vector(to_unsigned(2,8) ,
21321	 => std_logic_vector(to_unsigned(2,8) ,
21322	 => std_logic_vector(to_unsigned(1,8) ,
21323	 => std_logic_vector(to_unsigned(3,8) ,
21324	 => std_logic_vector(to_unsigned(45,8) ,
21325	 => std_logic_vector(to_unsigned(111,8) ,
21326	 => std_logic_vector(to_unsigned(118,8) ,
21327	 => std_logic_vector(to_unsigned(114,8) ,
21328	 => std_logic_vector(to_unsigned(103,8) ,
21329	 => std_logic_vector(to_unsigned(91,8) ,
21330	 => std_logic_vector(to_unsigned(92,8) ,
21331	 => std_logic_vector(to_unsigned(88,8) ,
21332	 => std_logic_vector(to_unsigned(93,8) ,
21333	 => std_logic_vector(to_unsigned(96,8) ,
21334	 => std_logic_vector(to_unsigned(103,8) ,
21335	 => std_logic_vector(to_unsigned(105,8) ,
21336	 => std_logic_vector(to_unsigned(96,8) ,
21337	 => std_logic_vector(to_unsigned(99,8) ,
21338	 => std_logic_vector(to_unsigned(97,8) ,
21339	 => std_logic_vector(to_unsigned(99,8) ,
21340	 => std_logic_vector(to_unsigned(128,8) ,
21341	 => std_logic_vector(to_unsigned(58,8) ,
21342	 => std_logic_vector(to_unsigned(1,8) ,
21343	 => std_logic_vector(to_unsigned(1,8) ,
21344	 => std_logic_vector(to_unsigned(13,8) ,
21345	 => std_logic_vector(to_unsigned(13,8) ,
21346	 => std_logic_vector(to_unsigned(3,8) ,
21347	 => std_logic_vector(to_unsigned(4,8) ,
21348	 => std_logic_vector(to_unsigned(9,8) ,
21349	 => std_logic_vector(to_unsigned(10,8) ,
21350	 => std_logic_vector(to_unsigned(10,8) ,
21351	 => std_logic_vector(to_unsigned(15,8) ,
21352	 => std_logic_vector(to_unsigned(38,8) ,
21353	 => std_logic_vector(to_unsigned(46,8) ,
21354	 => std_logic_vector(to_unsigned(50,8) ,
21355	 => std_logic_vector(to_unsigned(69,8) ,
21356	 => std_logic_vector(to_unsigned(76,8) ,
21357	 => std_logic_vector(to_unsigned(108,8) ,
21358	 => std_logic_vector(to_unsigned(122,8) ,
21359	 => std_logic_vector(to_unsigned(124,8) ,
21360	 => std_logic_vector(to_unsigned(121,8) ,
21361	 => std_logic_vector(to_unsigned(112,8) ,
21362	 => std_logic_vector(to_unsigned(115,8) ,
21363	 => std_logic_vector(to_unsigned(114,8) ,
21364	 => std_logic_vector(to_unsigned(112,8) ,
21365	 => std_logic_vector(to_unsigned(107,8) ,
21366	 => std_logic_vector(to_unsigned(92,8) ,
21367	 => std_logic_vector(to_unsigned(101,8) ,
21368	 => std_logic_vector(to_unsigned(109,8) ,
21369	 => std_logic_vector(to_unsigned(124,8) ,
21370	 => std_logic_vector(to_unsigned(144,8) ,
21371	 => std_logic_vector(to_unsigned(156,8) ,
21372	 => std_logic_vector(to_unsigned(33,8) ,
21373	 => std_logic_vector(to_unsigned(1,8) ,
21374	 => std_logic_vector(to_unsigned(1,8) ,
21375	 => std_logic_vector(to_unsigned(52,8) ,
21376	 => std_logic_vector(to_unsigned(173,8) ,
21377	 => std_logic_vector(to_unsigned(130,8) ,
21378	 => std_logic_vector(to_unsigned(112,8) ,
21379	 => std_logic_vector(to_unsigned(119,8) ,
21380	 => std_logic_vector(to_unsigned(130,8) ,
21381	 => std_logic_vector(to_unsigned(128,8) ,
21382	 => std_logic_vector(to_unsigned(125,8) ,
21383	 => std_logic_vector(to_unsigned(125,8) ,
21384	 => std_logic_vector(to_unsigned(134,8) ,
21385	 => std_logic_vector(to_unsigned(133,8) ,
21386	 => std_logic_vector(to_unsigned(124,8) ,
21387	 => std_logic_vector(to_unsigned(124,8) ,
21388	 => std_logic_vector(to_unsigned(122,8) ,
21389	 => std_logic_vector(to_unsigned(99,8) ,
21390	 => std_logic_vector(to_unsigned(59,8) ,
21391	 => std_logic_vector(to_unsigned(81,8) ,
21392	 => std_logic_vector(to_unsigned(41,8) ,
21393	 => std_logic_vector(to_unsigned(1,8) ,
21394	 => std_logic_vector(to_unsigned(1,8) ,
21395	 => std_logic_vector(to_unsigned(1,8) ,
21396	 => std_logic_vector(to_unsigned(1,8) ,
21397	 => std_logic_vector(to_unsigned(3,8) ,
21398	 => std_logic_vector(to_unsigned(8,8) ,
21399	 => std_logic_vector(to_unsigned(8,8) ,
21400	 => std_logic_vector(to_unsigned(11,8) ,
21401	 => std_logic_vector(to_unsigned(16,8) ,
21402	 => std_logic_vector(to_unsigned(12,8) ,
21403	 => std_logic_vector(to_unsigned(12,8) ,
21404	 => std_logic_vector(to_unsigned(7,8) ,
21405	 => std_logic_vector(to_unsigned(2,8) ,
21406	 => std_logic_vector(to_unsigned(3,8) ,
21407	 => std_logic_vector(to_unsigned(14,8) ,
21408	 => std_logic_vector(to_unsigned(91,8) ,
21409	 => std_logic_vector(to_unsigned(105,8) ,
21410	 => std_logic_vector(to_unsigned(97,8) ,
21411	 => std_logic_vector(to_unsigned(90,8) ,
21412	 => std_logic_vector(to_unsigned(86,8) ,
21413	 => std_logic_vector(to_unsigned(85,8) ,
21414	 => std_logic_vector(to_unsigned(88,8) ,
21415	 => std_logic_vector(to_unsigned(87,8) ,
21416	 => std_logic_vector(to_unsigned(95,8) ,
21417	 => std_logic_vector(to_unsigned(99,8) ,
21418	 => std_logic_vector(to_unsigned(91,8) ,
21419	 => std_logic_vector(to_unsigned(91,8) ,
21420	 => std_logic_vector(to_unsigned(97,8) ,
21421	 => std_logic_vector(to_unsigned(136,8) ,
21422	 => std_logic_vector(to_unsigned(147,8) ,
21423	 => std_logic_vector(to_unsigned(125,8) ,
21424	 => std_logic_vector(to_unsigned(104,8) ,
21425	 => std_logic_vector(to_unsigned(127,8) ,
21426	 => std_logic_vector(to_unsigned(154,8) ,
21427	 => std_logic_vector(to_unsigned(152,8) ,
21428	 => std_logic_vector(to_unsigned(146,8) ,
21429	 => std_logic_vector(to_unsigned(121,8) ,
21430	 => std_logic_vector(to_unsigned(114,8) ,
21431	 => std_logic_vector(to_unsigned(134,8) ,
21432	 => std_logic_vector(to_unsigned(108,8) ,
21433	 => std_logic_vector(to_unsigned(95,8) ,
21434	 => std_logic_vector(to_unsigned(91,8) ,
21435	 => std_logic_vector(to_unsigned(85,8) ,
21436	 => std_logic_vector(to_unsigned(97,8) ,
21437	 => std_logic_vector(to_unsigned(118,8) ,
21438	 => std_logic_vector(to_unsigned(92,8) ,
21439	 => std_logic_vector(to_unsigned(69,8) ,
21440	 => std_logic_vector(to_unsigned(76,8) ,
21441	 => std_logic_vector(to_unsigned(154,8) ,
21442	 => std_logic_vector(to_unsigned(147,8) ,
21443	 => std_logic_vector(to_unsigned(146,8) ,
21444	 => std_logic_vector(to_unsigned(151,8) ,
21445	 => std_logic_vector(to_unsigned(157,8) ,
21446	 => std_logic_vector(to_unsigned(166,8) ,
21447	 => std_logic_vector(to_unsigned(163,8) ,
21448	 => std_logic_vector(to_unsigned(168,8) ,
21449	 => std_logic_vector(to_unsigned(152,8) ,
21450	 => std_logic_vector(to_unsigned(121,8) ,
21451	 => std_logic_vector(to_unsigned(105,8) ,
21452	 => std_logic_vector(to_unsigned(88,8) ,
21453	 => std_logic_vector(to_unsigned(60,8) ,
21454	 => std_logic_vector(to_unsigned(13,8) ,
21455	 => std_logic_vector(to_unsigned(4,8) ,
21456	 => std_logic_vector(to_unsigned(8,8) ,
21457	 => std_logic_vector(to_unsigned(14,8) ,
21458	 => std_logic_vector(to_unsigned(25,8) ,
21459	 => std_logic_vector(to_unsigned(33,8) ,
21460	 => std_logic_vector(to_unsigned(24,8) ,
21461	 => std_logic_vector(to_unsigned(22,8) ,
21462	 => std_logic_vector(to_unsigned(6,8) ,
21463	 => std_logic_vector(to_unsigned(6,8) ,
21464	 => std_logic_vector(to_unsigned(15,8) ,
21465	 => std_logic_vector(to_unsigned(6,8) ,
21466	 => std_logic_vector(to_unsigned(6,8) ,
21467	 => std_logic_vector(to_unsigned(13,8) ,
21468	 => std_logic_vector(to_unsigned(39,8) ,
21469	 => std_logic_vector(to_unsigned(32,8) ,
21470	 => std_logic_vector(to_unsigned(8,8) ,
21471	 => std_logic_vector(to_unsigned(14,8) ,
21472	 => std_logic_vector(to_unsigned(34,8) ,
21473	 => std_logic_vector(to_unsigned(21,8) ,
21474	 => std_logic_vector(to_unsigned(14,8) ,
21475	 => std_logic_vector(to_unsigned(10,8) ,
21476	 => std_logic_vector(to_unsigned(14,8) ,
21477	 => std_logic_vector(to_unsigned(24,8) ,
21478	 => std_logic_vector(to_unsigned(24,8) ,
21479	 => std_logic_vector(to_unsigned(45,8) ,
21480	 => std_logic_vector(to_unsigned(32,8) ,
21481	 => std_logic_vector(to_unsigned(5,8) ,
21482	 => std_logic_vector(to_unsigned(12,8) ,
21483	 => std_logic_vector(to_unsigned(58,8) ,
21484	 => std_logic_vector(to_unsigned(74,8) ,
21485	 => std_logic_vector(to_unsigned(63,8) ,
21486	 => std_logic_vector(to_unsigned(93,8) ,
21487	 => std_logic_vector(to_unsigned(93,8) ,
21488	 => std_logic_vector(to_unsigned(122,8) ,
21489	 => std_logic_vector(to_unsigned(175,8) ,
21490	 => std_logic_vector(to_unsigned(163,8) ,
21491	 => std_logic_vector(to_unsigned(163,8) ,
21492	 => std_logic_vector(to_unsigned(163,8) ,
21493	 => std_logic_vector(to_unsigned(163,8) ,
21494	 => std_logic_vector(to_unsigned(171,8) ,
21495	 => std_logic_vector(to_unsigned(159,8) ,
21496	 => std_logic_vector(to_unsigned(170,8) ,
21497	 => std_logic_vector(to_unsigned(170,8) ,
21498	 => std_logic_vector(to_unsigned(21,8) ,
21499	 => std_logic_vector(to_unsigned(0,8) ,
21500	 => std_logic_vector(to_unsigned(4,8) ,
21501	 => std_logic_vector(to_unsigned(5,8) ,
21502	 => std_logic_vector(to_unsigned(6,8) ,
21503	 => std_logic_vector(to_unsigned(8,8) ,
21504	 => std_logic_vector(to_unsigned(15,8) ,
21505	 => std_logic_vector(to_unsigned(13,8) ,
21506	 => std_logic_vector(to_unsigned(22,8) ,
21507	 => std_logic_vector(to_unsigned(46,8) ,
21508	 => std_logic_vector(to_unsigned(27,8) ,
21509	 => std_logic_vector(to_unsigned(35,8) ,
21510	 => std_logic_vector(to_unsigned(70,8) ,
21511	 => std_logic_vector(to_unsigned(104,8) ,
21512	 => std_logic_vector(to_unsigned(151,8) ,
21513	 => std_logic_vector(to_unsigned(159,8) ,
21514	 => std_logic_vector(to_unsigned(161,8) ,
21515	 => std_logic_vector(to_unsigned(156,8) ,
21516	 => std_logic_vector(to_unsigned(154,8) ,
21517	 => std_logic_vector(to_unsigned(127,8) ,
21518	 => std_logic_vector(to_unsigned(154,8) ,
21519	 => std_logic_vector(to_unsigned(170,8) ,
21520	 => std_logic_vector(to_unsigned(164,8) ,
21521	 => std_logic_vector(to_unsigned(166,8) ,
21522	 => std_logic_vector(to_unsigned(161,8) ,
21523	 => std_logic_vector(to_unsigned(163,8) ,
21524	 => std_logic_vector(to_unsigned(166,8) ,
21525	 => std_logic_vector(to_unsigned(163,8) ,
21526	 => std_logic_vector(to_unsigned(168,8) ,
21527	 => std_logic_vector(to_unsigned(168,8) ,
21528	 => std_logic_vector(to_unsigned(161,8) ,
21529	 => std_logic_vector(to_unsigned(163,8) ,
21530	 => std_logic_vector(to_unsigned(157,8) ,
21531	 => std_logic_vector(to_unsigned(166,8) ,
21532	 => std_logic_vector(to_unsigned(122,8) ,
21533	 => std_logic_vector(to_unsigned(40,8) ,
21534	 => std_logic_vector(to_unsigned(17,8) ,
21535	 => std_logic_vector(to_unsigned(4,8) ,
21536	 => std_logic_vector(to_unsigned(3,8) ,
21537	 => std_logic_vector(to_unsigned(6,8) ,
21538	 => std_logic_vector(to_unsigned(7,8) ,
21539	 => std_logic_vector(to_unsigned(15,8) ,
21540	 => std_logic_vector(to_unsigned(80,8) ,
21541	 => std_logic_vector(to_unsigned(173,8) ,
21542	 => std_logic_vector(to_unsigned(171,8) ,
21543	 => std_logic_vector(to_unsigned(168,8) ,
21544	 => std_logic_vector(to_unsigned(171,8) ,
21545	 => std_logic_vector(to_unsigned(168,8) ,
21546	 => std_logic_vector(to_unsigned(164,8) ,
21547	 => std_logic_vector(to_unsigned(168,8) ,
21548	 => std_logic_vector(to_unsigned(171,8) ,
21549	 => std_logic_vector(to_unsigned(166,8) ,
21550	 => std_logic_vector(to_unsigned(164,8) ,
21551	 => std_logic_vector(to_unsigned(166,8) ,
21552	 => std_logic_vector(to_unsigned(164,8) ,
21553	 => std_logic_vector(to_unsigned(163,8) ,
21554	 => std_logic_vector(to_unsigned(170,8) ,
21555	 => std_logic_vector(to_unsigned(157,8) ,
21556	 => std_logic_vector(to_unsigned(152,8) ,
21557	 => std_logic_vector(to_unsigned(154,8) ,
21558	 => std_logic_vector(to_unsigned(121,8) ,
21559	 => std_logic_vector(to_unsigned(134,8) ,
21560	 => std_logic_vector(to_unsigned(121,8) ,
21561	 => std_logic_vector(to_unsigned(78,8) ,
21562	 => std_logic_vector(to_unsigned(38,8) ,
21563	 => std_logic_vector(to_unsigned(40,8) ,
21564	 => std_logic_vector(to_unsigned(62,8) ,
21565	 => std_logic_vector(to_unsigned(50,8) ,
21566	 => std_logic_vector(to_unsigned(19,8) ,
21567	 => std_logic_vector(to_unsigned(19,8) ,
21568	 => std_logic_vector(to_unsigned(124,8) ,
21569	 => std_logic_vector(to_unsigned(164,8) ,
21570	 => std_logic_vector(to_unsigned(138,8) ,
21571	 => std_logic_vector(to_unsigned(122,8) ,
21572	 => std_logic_vector(to_unsigned(133,8) ,
21573	 => std_logic_vector(to_unsigned(149,8) ,
21574	 => std_logic_vector(to_unsigned(147,8) ,
21575	 => std_logic_vector(to_unsigned(149,8) ,
21576	 => std_logic_vector(to_unsigned(142,8) ,
21577	 => std_logic_vector(to_unsigned(136,8) ,
21578	 => std_logic_vector(to_unsigned(144,8) ,
21579	 => std_logic_vector(to_unsigned(103,8) ,
21580	 => std_logic_vector(to_unsigned(72,8) ,
21581	 => std_logic_vector(to_unsigned(131,8) ,
21582	 => std_logic_vector(to_unsigned(136,8) ,
21583	 => std_logic_vector(to_unsigned(59,8) ,
21584	 => std_logic_vector(to_unsigned(13,8) ,
21585	 => std_logic_vector(to_unsigned(23,8) ,
21586	 => std_logic_vector(to_unsigned(67,8) ,
21587	 => std_logic_vector(to_unsigned(99,8) ,
21588	 => std_logic_vector(to_unsigned(101,8) ,
21589	 => std_logic_vector(to_unsigned(76,8) ,
21590	 => std_logic_vector(to_unsigned(19,8) ,
21591	 => std_logic_vector(to_unsigned(24,8) ,
21592	 => std_logic_vector(to_unsigned(43,8) ,
21593	 => std_logic_vector(to_unsigned(26,8) ,
21594	 => std_logic_vector(to_unsigned(118,8) ,
21595	 => std_logic_vector(to_unsigned(173,8) ,
21596	 => std_logic_vector(to_unsigned(159,8) ,
21597	 => std_logic_vector(to_unsigned(151,8) ,
21598	 => std_logic_vector(to_unsigned(138,8) ,
21599	 => std_logic_vector(to_unsigned(142,8) ,
21600	 => std_logic_vector(to_unsigned(130,8) ,
21601	 => std_logic_vector(to_unsigned(105,8) ,
21602	 => std_logic_vector(to_unsigned(97,8) ,
21603	 => std_logic_vector(to_unsigned(90,8) ,
21604	 => std_logic_vector(to_unsigned(91,8) ,
21605	 => std_logic_vector(to_unsigned(59,8) ,
21606	 => std_logic_vector(to_unsigned(15,8) ,
21607	 => std_logic_vector(to_unsigned(4,8) ,
21608	 => std_logic_vector(to_unsigned(8,8) ,
21609	 => std_logic_vector(to_unsigned(19,8) ,
21610	 => std_logic_vector(to_unsigned(14,8) ,
21611	 => std_logic_vector(to_unsigned(6,8) ,
21612	 => std_logic_vector(to_unsigned(3,8) ,
21613	 => std_logic_vector(to_unsigned(9,8) ,
21614	 => std_logic_vector(to_unsigned(8,8) ,
21615	 => std_logic_vector(to_unsigned(16,8) ,
21616	 => std_logic_vector(to_unsigned(122,8) ,
21617	 => std_logic_vector(to_unsigned(152,8) ,
21618	 => std_logic_vector(to_unsigned(147,8) ,
21619	 => std_logic_vector(to_unsigned(139,8) ,
21620	 => std_logic_vector(to_unsigned(142,8) ,
21621	 => std_logic_vector(to_unsigned(136,8) ,
21622	 => std_logic_vector(to_unsigned(127,8) ,
21623	 => std_logic_vector(to_unsigned(128,8) ,
21624	 => std_logic_vector(to_unsigned(114,8) ,
21625	 => std_logic_vector(to_unsigned(93,8) ,
21626	 => std_logic_vector(to_unsigned(88,8) ,
21627	 => std_logic_vector(to_unsigned(95,8) ,
21628	 => std_logic_vector(to_unsigned(88,8) ,
21629	 => std_logic_vector(to_unsigned(87,8) ,
21630	 => std_logic_vector(to_unsigned(92,8) ,
21631	 => std_logic_vector(to_unsigned(95,8) ,
21632	 => std_logic_vector(to_unsigned(99,8) ,
21633	 => std_logic_vector(to_unsigned(22,8) ,
21634	 => std_logic_vector(to_unsigned(0,8) ,
21635	 => std_logic_vector(to_unsigned(1,8) ,
21636	 => std_logic_vector(to_unsigned(1,8) ,
21637	 => std_logic_vector(to_unsigned(0,8) ,
21638	 => std_logic_vector(to_unsigned(0,8) ,
21639	 => std_logic_vector(to_unsigned(0,8) ,
21640	 => std_logic_vector(to_unsigned(1,8) ,
21641	 => std_logic_vector(to_unsigned(3,8) ,
21642	 => std_logic_vector(to_unsigned(4,8) ,
21643	 => std_logic_vector(to_unsigned(1,8) ,
21644	 => std_logic_vector(to_unsigned(14,8) ,
21645	 => std_logic_vector(to_unsigned(118,8) ,
21646	 => std_logic_vector(to_unsigned(130,8) ,
21647	 => std_logic_vector(to_unsigned(118,8) ,
21648	 => std_logic_vector(to_unsigned(115,8) ,
21649	 => std_logic_vector(to_unsigned(114,8) ,
21650	 => std_logic_vector(to_unsigned(109,8) ,
21651	 => std_logic_vector(to_unsigned(112,8) ,
21652	 => std_logic_vector(to_unsigned(112,8) ,
21653	 => std_logic_vector(to_unsigned(112,8) ,
21654	 => std_logic_vector(to_unsigned(122,8) ,
21655	 => std_logic_vector(to_unsigned(122,8) ,
21656	 => std_logic_vector(to_unsigned(116,8) ,
21657	 => std_logic_vector(to_unsigned(121,8) ,
21658	 => std_logic_vector(to_unsigned(118,8) ,
21659	 => std_logic_vector(to_unsigned(119,8) ,
21660	 => std_logic_vector(to_unsigned(133,8) ,
21661	 => std_logic_vector(to_unsigned(108,8) ,
21662	 => std_logic_vector(to_unsigned(63,8) ,
21663	 => std_logic_vector(to_unsigned(29,8) ,
21664	 => std_logic_vector(to_unsigned(14,8) ,
21665	 => std_logic_vector(to_unsigned(41,8) ,
21666	 => std_logic_vector(to_unsigned(23,8) ,
21667	 => std_logic_vector(to_unsigned(4,8) ,
21668	 => std_logic_vector(to_unsigned(2,8) ,
21669	 => std_logic_vector(to_unsigned(4,8) ,
21670	 => std_logic_vector(to_unsigned(8,8) ,
21671	 => std_logic_vector(to_unsigned(15,8) ,
21672	 => std_logic_vector(to_unsigned(35,8) ,
21673	 => std_logic_vector(to_unsigned(55,8) ,
21674	 => std_logic_vector(to_unsigned(58,8) ,
21675	 => std_logic_vector(to_unsigned(60,8) ,
21676	 => std_logic_vector(to_unsigned(62,8) ,
21677	 => std_logic_vector(to_unsigned(87,8) ,
21678	 => std_logic_vector(to_unsigned(125,8) ,
21679	 => std_logic_vector(to_unsigned(131,8) ,
21680	 => std_logic_vector(to_unsigned(121,8) ,
21681	 => std_logic_vector(to_unsigned(109,8) ,
21682	 => std_logic_vector(to_unsigned(114,8) ,
21683	 => std_logic_vector(to_unsigned(118,8) ,
21684	 => std_logic_vector(to_unsigned(115,8) ,
21685	 => std_logic_vector(to_unsigned(112,8) ,
21686	 => std_logic_vector(to_unsigned(104,8) ,
21687	 => std_logic_vector(to_unsigned(111,8) ,
21688	 => std_logic_vector(to_unsigned(125,8) ,
21689	 => std_logic_vector(to_unsigned(147,8) ,
21690	 => std_logic_vector(to_unsigned(147,8) ,
21691	 => std_logic_vector(to_unsigned(173,8) ,
21692	 => std_logic_vector(to_unsigned(79,8) ,
21693	 => std_logic_vector(to_unsigned(2,8) ,
21694	 => std_logic_vector(to_unsigned(1,8) ,
21695	 => std_logic_vector(to_unsigned(29,8) ,
21696	 => std_logic_vector(to_unsigned(175,8) ,
21697	 => std_logic_vector(to_unsigned(159,8) ,
21698	 => std_logic_vector(to_unsigned(141,8) ,
21699	 => std_logic_vector(to_unsigned(138,8) ,
21700	 => std_logic_vector(to_unsigned(136,8) ,
21701	 => std_logic_vector(to_unsigned(136,8) ,
21702	 => std_logic_vector(to_unsigned(138,8) ,
21703	 => std_logic_vector(to_unsigned(136,8) ,
21704	 => std_logic_vector(to_unsigned(134,8) ,
21705	 => std_logic_vector(to_unsigned(131,8) ,
21706	 => std_logic_vector(to_unsigned(134,8) ,
21707	 => std_logic_vector(to_unsigned(133,8) ,
21708	 => std_logic_vector(to_unsigned(130,8) ,
21709	 => std_logic_vector(to_unsigned(87,8) ,
21710	 => std_logic_vector(to_unsigned(48,8) ,
21711	 => std_logic_vector(to_unsigned(92,8) ,
21712	 => std_logic_vector(to_unsigned(48,8) ,
21713	 => std_logic_vector(to_unsigned(1,8) ,
21714	 => std_logic_vector(to_unsigned(0,8) ,
21715	 => std_logic_vector(to_unsigned(0,8) ,
21716	 => std_logic_vector(to_unsigned(2,8) ,
21717	 => std_logic_vector(to_unsigned(6,8) ,
21718	 => std_logic_vector(to_unsigned(17,8) ,
21719	 => std_logic_vector(to_unsigned(15,8) ,
21720	 => std_logic_vector(to_unsigned(17,8) ,
21721	 => std_logic_vector(to_unsigned(30,8) ,
21722	 => std_logic_vector(to_unsigned(32,8) ,
21723	 => std_logic_vector(to_unsigned(27,8) ,
21724	 => std_logic_vector(to_unsigned(20,8) ,
21725	 => std_logic_vector(to_unsigned(7,8) ,
21726	 => std_logic_vector(to_unsigned(5,8) ,
21727	 => std_logic_vector(to_unsigned(12,8) ,
21728	 => std_logic_vector(to_unsigned(61,8) ,
21729	 => std_logic_vector(to_unsigned(121,8) ,
21730	 => std_logic_vector(to_unsigned(114,8) ,
21731	 => std_logic_vector(to_unsigned(105,8) ,
21732	 => std_logic_vector(to_unsigned(88,8) ,
21733	 => std_logic_vector(to_unsigned(78,8) ,
21734	 => std_logic_vector(to_unsigned(86,8) ,
21735	 => std_logic_vector(to_unsigned(92,8) ,
21736	 => std_logic_vector(to_unsigned(97,8) ,
21737	 => std_logic_vector(to_unsigned(101,8) ,
21738	 => std_logic_vector(to_unsigned(93,8) ,
21739	 => std_logic_vector(to_unsigned(92,8) ,
21740	 => std_logic_vector(to_unsigned(95,8) ,
21741	 => std_logic_vector(to_unsigned(115,8) ,
21742	 => std_logic_vector(to_unsigned(128,8) ,
21743	 => std_logic_vector(to_unsigned(100,8) ,
21744	 => std_logic_vector(to_unsigned(90,8) ,
21745	 => std_logic_vector(to_unsigned(101,8) ,
21746	 => std_logic_vector(to_unsigned(119,8) ,
21747	 => std_logic_vector(to_unsigned(116,8) ,
21748	 => std_logic_vector(to_unsigned(105,8) ,
21749	 => std_logic_vector(to_unsigned(99,8) ,
21750	 => std_logic_vector(to_unsigned(96,8) ,
21751	 => std_logic_vector(to_unsigned(125,8) ,
21752	 => std_logic_vector(to_unsigned(131,8) ,
21753	 => std_logic_vector(to_unsigned(92,8) ,
21754	 => std_logic_vector(to_unsigned(82,8) ,
21755	 => std_logic_vector(to_unsigned(90,8) ,
21756	 => std_logic_vector(to_unsigned(104,8) ,
21757	 => std_logic_vector(to_unsigned(103,8) ,
21758	 => std_logic_vector(to_unsigned(100,8) ,
21759	 => std_logic_vector(to_unsigned(115,8) ,
21760	 => std_logic_vector(to_unsigned(118,8) ,
21761	 => std_logic_vector(to_unsigned(154,8) ,
21762	 => std_logic_vector(to_unsigned(151,8) ,
21763	 => std_logic_vector(to_unsigned(152,8) ,
21764	 => std_logic_vector(to_unsigned(156,8) ,
21765	 => std_logic_vector(to_unsigned(161,8) ,
21766	 => std_logic_vector(to_unsigned(163,8) ,
21767	 => std_logic_vector(to_unsigned(164,8) ,
21768	 => std_logic_vector(to_unsigned(159,8) ,
21769	 => std_logic_vector(to_unsigned(125,8) ,
21770	 => std_logic_vector(to_unsigned(95,8) ,
21771	 => std_logic_vector(to_unsigned(77,8) ,
21772	 => std_logic_vector(to_unsigned(49,8) ,
21773	 => std_logic_vector(to_unsigned(38,8) ,
21774	 => std_logic_vector(to_unsigned(28,8) ,
21775	 => std_logic_vector(to_unsigned(18,8) ,
21776	 => std_logic_vector(to_unsigned(11,8) ,
21777	 => std_logic_vector(to_unsigned(8,8) ,
21778	 => std_logic_vector(to_unsigned(4,8) ,
21779	 => std_logic_vector(to_unsigned(3,8) ,
21780	 => std_logic_vector(to_unsigned(5,8) ,
21781	 => std_logic_vector(to_unsigned(1,8) ,
21782	 => std_logic_vector(to_unsigned(2,8) ,
21783	 => std_logic_vector(to_unsigned(6,8) ,
21784	 => std_logic_vector(to_unsigned(6,8) ,
21785	 => std_logic_vector(to_unsigned(4,8) ,
21786	 => std_logic_vector(to_unsigned(3,8) ,
21787	 => std_logic_vector(to_unsigned(6,8) ,
21788	 => std_logic_vector(to_unsigned(19,8) ,
21789	 => std_logic_vector(to_unsigned(13,8) ,
21790	 => std_logic_vector(to_unsigned(7,8) ,
21791	 => std_logic_vector(to_unsigned(16,8) ,
21792	 => std_logic_vector(to_unsigned(16,8) ,
21793	 => std_logic_vector(to_unsigned(11,8) ,
21794	 => std_logic_vector(to_unsigned(10,8) ,
21795	 => std_logic_vector(to_unsigned(11,8) ,
21796	 => std_logic_vector(to_unsigned(16,8) ,
21797	 => std_logic_vector(to_unsigned(25,8) ,
21798	 => std_logic_vector(to_unsigned(23,8) ,
21799	 => std_logic_vector(to_unsigned(35,8) ,
21800	 => std_logic_vector(to_unsigned(33,8) ,
21801	 => std_logic_vector(to_unsigned(6,8) ,
21802	 => std_logic_vector(to_unsigned(32,8) ,
21803	 => std_logic_vector(to_unsigned(93,8) ,
21804	 => std_logic_vector(to_unsigned(51,8) ,
21805	 => std_logic_vector(to_unsigned(51,8) ,
21806	 => std_logic_vector(to_unsigned(80,8) ,
21807	 => std_logic_vector(to_unsigned(67,8) ,
21808	 => std_logic_vector(to_unsigned(43,8) ,
21809	 => std_logic_vector(to_unsigned(100,8) ,
21810	 => std_logic_vector(to_unsigned(175,8) ,
21811	 => std_logic_vector(to_unsigned(166,8) ,
21812	 => std_logic_vector(to_unsigned(163,8) ,
21813	 => std_logic_vector(to_unsigned(170,8) ,
21814	 => std_logic_vector(to_unsigned(141,8) ,
21815	 => std_logic_vector(to_unsigned(38,8) ,
21816	 => std_logic_vector(to_unsigned(85,8) ,
21817	 => std_logic_vector(to_unsigned(200,8) ,
21818	 => std_logic_vector(to_unsigned(80,8) ,
21819	 => std_logic_vector(to_unsigned(2,8) ,
21820	 => std_logic_vector(to_unsigned(2,8) ,
21821	 => std_logic_vector(to_unsigned(3,8) ,
21822	 => std_logic_vector(to_unsigned(3,8) ,
21823	 => std_logic_vector(to_unsigned(3,8) ,
21824	 => std_logic_vector(to_unsigned(7,8) ,
21825	 => std_logic_vector(to_unsigned(4,8) ,
21826	 => std_logic_vector(to_unsigned(16,8) ,
21827	 => std_logic_vector(to_unsigned(157,8) ,
21828	 => std_logic_vector(to_unsigned(72,8) ,
21829	 => std_logic_vector(to_unsigned(29,8) ,
21830	 => std_logic_vector(to_unsigned(119,8) ,
21831	 => std_logic_vector(to_unsigned(139,8) ,
21832	 => std_logic_vector(to_unsigned(146,8) ,
21833	 => std_logic_vector(to_unsigned(142,8) ,
21834	 => std_logic_vector(to_unsigned(156,8) ,
21835	 => std_logic_vector(to_unsigned(151,8) ,
21836	 => std_logic_vector(to_unsigned(147,8) ,
21837	 => std_logic_vector(to_unsigned(161,8) ,
21838	 => std_logic_vector(to_unsigned(151,8) ,
21839	 => std_logic_vector(to_unsigned(159,8) ,
21840	 => std_logic_vector(to_unsigned(164,8) ,
21841	 => std_logic_vector(to_unsigned(170,8) ,
21842	 => std_logic_vector(to_unsigned(168,8) ,
21843	 => std_logic_vector(to_unsigned(166,8) ,
21844	 => std_logic_vector(to_unsigned(164,8) ,
21845	 => std_logic_vector(to_unsigned(168,8) ,
21846	 => std_logic_vector(to_unsigned(170,8) ,
21847	 => std_logic_vector(to_unsigned(164,8) ,
21848	 => std_logic_vector(to_unsigned(161,8) ,
21849	 => std_logic_vector(to_unsigned(161,8) ,
21850	 => std_logic_vector(to_unsigned(161,8) ,
21851	 => std_logic_vector(to_unsigned(154,8) ,
21852	 => std_logic_vector(to_unsigned(103,8) ,
21853	 => std_logic_vector(to_unsigned(46,8) ,
21854	 => std_logic_vector(to_unsigned(55,8) ,
21855	 => std_logic_vector(to_unsigned(22,8) ,
21856	 => std_logic_vector(to_unsigned(8,8) ,
21857	 => std_logic_vector(to_unsigned(9,8) ,
21858	 => std_logic_vector(to_unsigned(10,8) ,
21859	 => std_logic_vector(to_unsigned(46,8) ,
21860	 => std_logic_vector(to_unsigned(151,8) ,
21861	 => std_logic_vector(to_unsigned(171,8) ,
21862	 => std_logic_vector(to_unsigned(164,8) ,
21863	 => std_logic_vector(to_unsigned(171,8) ,
21864	 => std_logic_vector(to_unsigned(163,8) ,
21865	 => std_logic_vector(to_unsigned(159,8) ,
21866	 => std_logic_vector(to_unsigned(170,8) ,
21867	 => std_logic_vector(to_unsigned(171,8) ,
21868	 => std_logic_vector(to_unsigned(171,8) ,
21869	 => std_logic_vector(to_unsigned(168,8) ,
21870	 => std_logic_vector(to_unsigned(164,8) ,
21871	 => std_logic_vector(to_unsigned(166,8) ,
21872	 => std_logic_vector(to_unsigned(163,8) ,
21873	 => std_logic_vector(to_unsigned(163,8) ,
21874	 => std_logic_vector(to_unsigned(170,8) ,
21875	 => std_logic_vector(to_unsigned(144,8) ,
21876	 => std_logic_vector(to_unsigned(96,8) ,
21877	 => std_logic_vector(to_unsigned(51,8) ,
21878	 => std_logic_vector(to_unsigned(57,8) ,
21879	 => std_logic_vector(to_unsigned(108,8) ,
21880	 => std_logic_vector(to_unsigned(105,8) ,
21881	 => std_logic_vector(to_unsigned(81,8) ,
21882	 => std_logic_vector(to_unsigned(67,8) ,
21883	 => std_logic_vector(to_unsigned(69,8) ,
21884	 => std_logic_vector(to_unsigned(92,8) ,
21885	 => std_logic_vector(to_unsigned(38,8) ,
21886	 => std_logic_vector(to_unsigned(10,8) ,
21887	 => std_logic_vector(to_unsigned(52,8) ,
21888	 => std_logic_vector(to_unsigned(181,8) ,
21889	 => std_logic_vector(to_unsigned(157,8) ,
21890	 => std_logic_vector(to_unsigned(141,8) ,
21891	 => std_logic_vector(to_unsigned(125,8) ,
21892	 => std_logic_vector(to_unsigned(131,8) ,
21893	 => std_logic_vector(to_unsigned(147,8) ,
21894	 => std_logic_vector(to_unsigned(151,8) ,
21895	 => std_logic_vector(to_unsigned(149,8) ,
21896	 => std_logic_vector(to_unsigned(144,8) ,
21897	 => std_logic_vector(to_unsigned(141,8) ,
21898	 => std_logic_vector(to_unsigned(149,8) ,
21899	 => std_logic_vector(to_unsigned(116,8) ,
21900	 => std_logic_vector(to_unsigned(28,8) ,
21901	 => std_logic_vector(to_unsigned(45,8) ,
21902	 => std_logic_vector(to_unsigned(38,8) ,
21903	 => std_logic_vector(to_unsigned(8,8) ,
21904	 => std_logic_vector(to_unsigned(6,8) ,
21905	 => std_logic_vector(to_unsigned(10,8) ,
21906	 => std_logic_vector(to_unsigned(21,8) ,
21907	 => std_logic_vector(to_unsigned(40,8) ,
21908	 => std_logic_vector(to_unsigned(43,8) ,
21909	 => std_logic_vector(to_unsigned(35,8) ,
21910	 => std_logic_vector(to_unsigned(26,8) ,
21911	 => std_logic_vector(to_unsigned(8,8) ,
21912	 => std_logic_vector(to_unsigned(0,8) ,
21913	 => std_logic_vector(to_unsigned(14,8) ,
21914	 => std_logic_vector(to_unsigned(139,8) ,
21915	 => std_logic_vector(to_unsigned(152,8) ,
21916	 => std_logic_vector(to_unsigned(156,8) ,
21917	 => std_logic_vector(to_unsigned(149,8) ,
21918	 => std_logic_vector(to_unsigned(139,8) ,
21919	 => std_logic_vector(to_unsigned(152,8) ,
21920	 => std_logic_vector(to_unsigned(138,8) ,
21921	 => std_logic_vector(to_unsigned(99,8) ,
21922	 => std_logic_vector(to_unsigned(93,8) ,
21923	 => std_logic_vector(to_unsigned(91,8) ,
21924	 => std_logic_vector(to_unsigned(87,8) ,
21925	 => std_logic_vector(to_unsigned(39,8) ,
21926	 => std_logic_vector(to_unsigned(15,8) ,
21927	 => std_logic_vector(to_unsigned(9,8) ,
21928	 => std_logic_vector(to_unsigned(7,8) ,
21929	 => std_logic_vector(to_unsigned(8,8) ,
21930	 => std_logic_vector(to_unsigned(5,8) ,
21931	 => std_logic_vector(to_unsigned(7,8) ,
21932	 => std_logic_vector(to_unsigned(9,8) ,
21933	 => std_logic_vector(to_unsigned(5,8) ,
21934	 => std_logic_vector(to_unsigned(3,8) ,
21935	 => std_logic_vector(to_unsigned(12,8) ,
21936	 => std_logic_vector(to_unsigned(64,8) ,
21937	 => std_logic_vector(to_unsigned(121,8) ,
21938	 => std_logic_vector(to_unsigned(152,8) ,
21939	 => std_logic_vector(to_unsigned(142,8) ,
21940	 => std_logic_vector(to_unsigned(146,8) ,
21941	 => std_logic_vector(to_unsigned(118,8) ,
21942	 => std_logic_vector(to_unsigned(105,8) ,
21943	 => std_logic_vector(to_unsigned(125,8) ,
21944	 => std_logic_vector(to_unsigned(112,8) ,
21945	 => std_logic_vector(to_unsigned(101,8) ,
21946	 => std_logic_vector(to_unsigned(91,8) ,
21947	 => std_logic_vector(to_unsigned(92,8) ,
21948	 => std_logic_vector(to_unsigned(95,8) ,
21949	 => std_logic_vector(to_unsigned(91,8) ,
21950	 => std_logic_vector(to_unsigned(91,8) ,
21951	 => std_logic_vector(to_unsigned(104,8) ,
21952	 => std_logic_vector(to_unsigned(93,8) ,
21953	 => std_logic_vector(to_unsigned(6,8) ,
21954	 => std_logic_vector(to_unsigned(0,8) ,
21955	 => std_logic_vector(to_unsigned(1,8) ,
21956	 => std_logic_vector(to_unsigned(0,8) ,
21957	 => std_logic_vector(to_unsigned(0,8) ,
21958	 => std_logic_vector(to_unsigned(1,8) ,
21959	 => std_logic_vector(to_unsigned(1,8) ,
21960	 => std_logic_vector(to_unsigned(2,8) ,
21961	 => std_logic_vector(to_unsigned(4,8) ,
21962	 => std_logic_vector(to_unsigned(5,8) ,
21963	 => std_logic_vector(to_unsigned(3,8) ,
21964	 => std_logic_vector(to_unsigned(13,8) ,
21965	 => std_logic_vector(to_unsigned(78,8) ,
21966	 => std_logic_vector(to_unsigned(114,8) ,
21967	 => std_logic_vector(to_unsigned(119,8) ,
21968	 => std_logic_vector(to_unsigned(122,8) ,
21969	 => std_logic_vector(to_unsigned(116,8) ,
21970	 => std_logic_vector(to_unsigned(114,8) ,
21971	 => std_logic_vector(to_unsigned(118,8) ,
21972	 => std_logic_vector(to_unsigned(115,8) ,
21973	 => std_logic_vector(to_unsigned(119,8) ,
21974	 => std_logic_vector(to_unsigned(119,8) ,
21975	 => std_logic_vector(to_unsigned(124,8) ,
21976	 => std_logic_vector(to_unsigned(128,8) ,
21977	 => std_logic_vector(to_unsigned(128,8) ,
21978	 => std_logic_vector(to_unsigned(127,8) ,
21979	 => std_logic_vector(to_unsigned(127,8) ,
21980	 => std_logic_vector(to_unsigned(127,8) ,
21981	 => std_logic_vector(to_unsigned(127,8) ,
21982	 => std_logic_vector(to_unsigned(168,8) ,
21983	 => std_logic_vector(to_unsigned(80,8) ,
21984	 => std_logic_vector(to_unsigned(3,8) ,
21985	 => std_logic_vector(to_unsigned(10,8) ,
21986	 => std_logic_vector(to_unsigned(24,8) ,
21987	 => std_logic_vector(to_unsigned(28,8) ,
21988	 => std_logic_vector(to_unsigned(14,8) ,
21989	 => std_logic_vector(to_unsigned(3,8) ,
21990	 => std_logic_vector(to_unsigned(2,8) ,
21991	 => std_logic_vector(to_unsigned(7,8) ,
21992	 => std_logic_vector(to_unsigned(16,8) ,
21993	 => std_logic_vector(to_unsigned(36,8) ,
21994	 => std_logic_vector(to_unsigned(44,8) ,
21995	 => std_logic_vector(to_unsigned(40,8) ,
21996	 => std_logic_vector(to_unsigned(58,8) ,
21997	 => std_logic_vector(to_unsigned(69,8) ,
21998	 => std_logic_vector(to_unsigned(112,8) ,
21999	 => std_logic_vector(to_unsigned(130,8) ,
22000	 => std_logic_vector(to_unsigned(118,8) ,
22001	 => std_logic_vector(to_unsigned(115,8) ,
22002	 => std_logic_vector(to_unsigned(121,8) ,
22003	 => std_logic_vector(to_unsigned(116,8) ,
22004	 => std_logic_vector(to_unsigned(114,8) ,
22005	 => std_logic_vector(to_unsigned(116,8) ,
22006	 => std_logic_vector(to_unsigned(134,8) ,
22007	 => std_logic_vector(to_unsigned(142,8) ,
22008	 => std_logic_vector(to_unsigned(154,8) ,
22009	 => std_logic_vector(to_unsigned(149,8) ,
22010	 => std_logic_vector(to_unsigned(128,8) ,
22011	 => std_logic_vector(to_unsigned(157,8) ,
22012	 => std_logic_vector(to_unsigned(122,8) ,
22013	 => std_logic_vector(to_unsigned(6,8) ,
22014	 => std_logic_vector(to_unsigned(1,8) ,
22015	 => std_logic_vector(to_unsigned(13,8) ,
22016	 => std_logic_vector(to_unsigned(138,8) ,
22017	 => std_logic_vector(to_unsigned(173,8) ,
22018	 => std_logic_vector(to_unsigned(159,8) ,
22019	 => std_logic_vector(to_unsigned(151,8) ,
22020	 => std_logic_vector(to_unsigned(146,8) ,
22021	 => std_logic_vector(to_unsigned(149,8) ,
22022	 => std_logic_vector(to_unsigned(149,8) ,
22023	 => std_logic_vector(to_unsigned(149,8) ,
22024	 => std_logic_vector(to_unsigned(146,8) ,
22025	 => std_logic_vector(to_unsigned(144,8) ,
22026	 => std_logic_vector(to_unsigned(147,8) ,
22027	 => std_logic_vector(to_unsigned(146,8) ,
22028	 => std_logic_vector(to_unsigned(141,8) ,
22029	 => std_logic_vector(to_unsigned(124,8) ,
22030	 => std_logic_vector(to_unsigned(119,8) ,
22031	 => std_logic_vector(to_unsigned(111,8) ,
22032	 => std_logic_vector(to_unsigned(108,8) ,
22033	 => std_logic_vector(to_unsigned(66,8) ,
22034	 => std_logic_vector(to_unsigned(24,8) ,
22035	 => std_logic_vector(to_unsigned(5,8) ,
22036	 => std_logic_vector(to_unsigned(5,8) ,
22037	 => std_logic_vector(to_unsigned(7,8) ,
22038	 => std_logic_vector(to_unsigned(10,8) ,
22039	 => std_logic_vector(to_unsigned(13,8) ,
22040	 => std_logic_vector(to_unsigned(8,8) ,
22041	 => std_logic_vector(to_unsigned(8,8) ,
22042	 => std_logic_vector(to_unsigned(13,8) ,
22043	 => std_logic_vector(to_unsigned(18,8) ,
22044	 => std_logic_vector(to_unsigned(38,8) ,
22045	 => std_logic_vector(to_unsigned(33,8) ,
22046	 => std_logic_vector(to_unsigned(9,8) ,
22047	 => std_logic_vector(to_unsigned(6,8) ,
22048	 => std_logic_vector(to_unsigned(51,8) ,
22049	 => std_logic_vector(to_unsigned(124,8) ,
22050	 => std_logic_vector(to_unsigned(118,8) ,
22051	 => std_logic_vector(to_unsigned(114,8) ,
22052	 => std_logic_vector(to_unsigned(101,8) ,
22053	 => std_logic_vector(to_unsigned(77,8) ,
22054	 => std_logic_vector(to_unsigned(80,8) ,
22055	 => std_logic_vector(to_unsigned(97,8) ,
22056	 => std_logic_vector(to_unsigned(105,8) ,
22057	 => std_logic_vector(to_unsigned(107,8) ,
22058	 => std_logic_vector(to_unsigned(95,8) ,
22059	 => std_logic_vector(to_unsigned(95,8) ,
22060	 => std_logic_vector(to_unsigned(97,8) ,
22061	 => std_logic_vector(to_unsigned(97,8) ,
22062	 => std_logic_vector(to_unsigned(130,8) ,
22063	 => std_logic_vector(to_unsigned(131,8) ,
22064	 => std_logic_vector(to_unsigned(108,8) ,
22065	 => std_logic_vector(to_unsigned(90,8) ,
22066	 => std_logic_vector(to_unsigned(103,8) ,
22067	 => std_logic_vector(to_unsigned(122,8) ,
22068	 => std_logic_vector(to_unsigned(114,8) ,
22069	 => std_logic_vector(to_unsigned(122,8) ,
22070	 => std_logic_vector(to_unsigned(115,8) ,
22071	 => std_logic_vector(to_unsigned(108,8) ,
22072	 => std_logic_vector(to_unsigned(124,8) ,
22073	 => std_logic_vector(to_unsigned(115,8) ,
22074	 => std_logic_vector(to_unsigned(99,8) ,
22075	 => std_logic_vector(to_unsigned(91,8) ,
22076	 => std_logic_vector(to_unsigned(109,8) ,
22077	 => std_logic_vector(to_unsigned(115,8) ,
22078	 => std_logic_vector(to_unsigned(109,8) ,
22079	 => std_logic_vector(to_unsigned(141,8) ,
22080	 => std_logic_vector(to_unsigned(163,8) ,
22081	 => std_logic_vector(to_unsigned(156,8) ,
22082	 => std_logic_vector(to_unsigned(154,8) ,
22083	 => std_logic_vector(to_unsigned(154,8) ,
22084	 => std_logic_vector(to_unsigned(157,8) ,
22085	 => std_logic_vector(to_unsigned(159,8) ,
22086	 => std_logic_vector(to_unsigned(159,8) ,
22087	 => std_logic_vector(to_unsigned(170,8) ,
22088	 => std_logic_vector(to_unsigned(136,8) ,
22089	 => std_logic_vector(to_unsigned(85,8) ,
22090	 => std_logic_vector(to_unsigned(65,8) ,
22091	 => std_logic_vector(to_unsigned(52,8) ,
22092	 => std_logic_vector(to_unsigned(45,8) ,
22093	 => std_logic_vector(to_unsigned(31,8) ,
22094	 => std_logic_vector(to_unsigned(12,8) ,
22095	 => std_logic_vector(to_unsigned(16,8) ,
22096	 => std_logic_vector(to_unsigned(13,8) ,
22097	 => std_logic_vector(to_unsigned(12,8) ,
22098	 => std_logic_vector(to_unsigned(6,8) ,
22099	 => std_logic_vector(to_unsigned(6,8) ,
22100	 => std_logic_vector(to_unsigned(28,8) ,
22101	 => std_logic_vector(to_unsigned(14,8) ,
22102	 => std_logic_vector(to_unsigned(4,8) ,
22103	 => std_logic_vector(to_unsigned(3,8) ,
22104	 => std_logic_vector(to_unsigned(4,8) ,
22105	 => std_logic_vector(to_unsigned(7,8) ,
22106	 => std_logic_vector(to_unsigned(3,8) ,
22107	 => std_logic_vector(to_unsigned(2,8) ,
22108	 => std_logic_vector(to_unsigned(2,8) ,
22109	 => std_logic_vector(to_unsigned(5,8) ,
22110	 => std_logic_vector(to_unsigned(7,8) ,
22111	 => std_logic_vector(to_unsigned(4,8) ,
22112	 => std_logic_vector(to_unsigned(7,8) ,
22113	 => std_logic_vector(to_unsigned(10,8) ,
22114	 => std_logic_vector(to_unsigned(8,8) ,
22115	 => std_logic_vector(to_unsigned(8,8) ,
22116	 => std_logic_vector(to_unsigned(14,8) ,
22117	 => std_logic_vector(to_unsigned(32,8) ,
22118	 => std_logic_vector(to_unsigned(41,8) ,
22119	 => std_logic_vector(to_unsigned(45,8) ,
22120	 => std_logic_vector(to_unsigned(32,8) ,
22121	 => std_logic_vector(to_unsigned(8,8) ,
22122	 => std_logic_vector(to_unsigned(19,8) ,
22123	 => std_logic_vector(to_unsigned(25,8) ,
22124	 => std_logic_vector(to_unsigned(32,8) ,
22125	 => std_logic_vector(to_unsigned(56,8) ,
22126	 => std_logic_vector(to_unsigned(46,8) ,
22127	 => std_logic_vector(to_unsigned(51,8) ,
22128	 => std_logic_vector(to_unsigned(37,8) ,
22129	 => std_logic_vector(to_unsigned(30,8) ,
22130	 => std_logic_vector(to_unsigned(131,8) ,
22131	 => std_logic_vector(to_unsigned(177,8) ,
22132	 => std_logic_vector(to_unsigned(171,8) ,
22133	 => std_logic_vector(to_unsigned(152,8) ,
22134	 => std_logic_vector(to_unsigned(40,8) ,
22135	 => std_logic_vector(to_unsigned(2,8) ,
22136	 => std_logic_vector(to_unsigned(20,8) ,
22137	 => std_logic_vector(to_unsigned(166,8) ,
22138	 => std_logic_vector(to_unsigned(175,8) ,
22139	 => std_logic_vector(to_unsigned(50,8) ,
22140	 => std_logic_vector(to_unsigned(5,8) ,
22141	 => std_logic_vector(to_unsigned(4,8) ,
22142	 => std_logic_vector(to_unsigned(2,8) ,
22143	 => std_logic_vector(to_unsigned(2,8) ,
22144	 => std_logic_vector(to_unsigned(2,8) ,
22145	 => std_logic_vector(to_unsigned(6,8) ,
22146	 => std_logic_vector(to_unsigned(41,8) ,
22147	 => std_logic_vector(to_unsigned(64,8) ,
22148	 => std_logic_vector(to_unsigned(15,8) ,
22149	 => std_logic_vector(to_unsigned(12,8) ,
22150	 => std_logic_vector(to_unsigned(62,8) ,
22151	 => std_logic_vector(to_unsigned(141,8) ,
22152	 => std_logic_vector(to_unsigned(138,8) ,
22153	 => std_logic_vector(to_unsigned(127,8) ,
22154	 => std_logic_vector(to_unsigned(122,8) ,
22155	 => std_logic_vector(to_unsigned(115,8) ,
22156	 => std_logic_vector(to_unsigned(121,8) ,
22157	 => std_logic_vector(to_unsigned(149,8) ,
22158	 => std_logic_vector(to_unsigned(144,8) ,
22159	 => std_logic_vector(to_unsigned(152,8) ,
22160	 => std_logic_vector(to_unsigned(154,8) ,
22161	 => std_logic_vector(to_unsigned(159,8) ,
22162	 => std_logic_vector(to_unsigned(170,8) ,
22163	 => std_logic_vector(to_unsigned(163,8) ,
22164	 => std_logic_vector(to_unsigned(170,8) ,
22165	 => std_logic_vector(to_unsigned(166,8) ,
22166	 => std_logic_vector(to_unsigned(168,8) ,
22167	 => std_logic_vector(to_unsigned(164,8) ,
22168	 => std_logic_vector(to_unsigned(159,8) ,
22169	 => std_logic_vector(to_unsigned(161,8) ,
22170	 => std_logic_vector(to_unsigned(156,8) ,
22171	 => std_logic_vector(to_unsigned(141,8) ,
22172	 => std_logic_vector(to_unsigned(119,8) ,
22173	 => std_logic_vector(to_unsigned(90,8) ,
22174	 => std_logic_vector(to_unsigned(101,8) ,
22175	 => std_logic_vector(to_unsigned(53,8) ,
22176	 => std_logic_vector(to_unsigned(13,8) ,
22177	 => std_logic_vector(to_unsigned(28,8) ,
22178	 => std_logic_vector(to_unsigned(71,8) ,
22179	 => std_logic_vector(to_unsigned(168,8) ,
22180	 => std_logic_vector(to_unsigned(179,8) ,
22181	 => std_logic_vector(to_unsigned(159,8) ,
22182	 => std_logic_vector(to_unsigned(170,8) ,
22183	 => std_logic_vector(to_unsigned(173,8) ,
22184	 => std_logic_vector(to_unsigned(149,8) ,
22185	 => std_logic_vector(to_unsigned(139,8) ,
22186	 => std_logic_vector(to_unsigned(166,8) ,
22187	 => std_logic_vector(to_unsigned(170,8) ,
22188	 => std_logic_vector(to_unsigned(171,8) ,
22189	 => std_logic_vector(to_unsigned(171,8) ,
22190	 => std_logic_vector(to_unsigned(166,8) ,
22191	 => std_logic_vector(to_unsigned(164,8) ,
22192	 => std_logic_vector(to_unsigned(159,8) ,
22193	 => std_logic_vector(to_unsigned(164,8) ,
22194	 => std_logic_vector(to_unsigned(159,8) ,
22195	 => std_logic_vector(to_unsigned(95,8) ,
22196	 => std_logic_vector(to_unsigned(45,8) ,
22197	 => std_logic_vector(to_unsigned(30,8) ,
22198	 => std_logic_vector(to_unsigned(56,8) ,
22199	 => std_logic_vector(to_unsigned(68,8) ,
22200	 => std_logic_vector(to_unsigned(66,8) ,
22201	 => std_logic_vector(to_unsigned(55,8) ,
22202	 => std_logic_vector(to_unsigned(57,8) ,
22203	 => std_logic_vector(to_unsigned(60,8) ,
22204	 => std_logic_vector(to_unsigned(29,8) ,
22205	 => std_logic_vector(to_unsigned(16,8) ,
22206	 => std_logic_vector(to_unsigned(37,8) ,
22207	 => std_logic_vector(to_unsigned(85,8) ,
22208	 => std_logic_vector(to_unsigned(163,8) ,
22209	 => std_logic_vector(to_unsigned(156,8) ,
22210	 => std_logic_vector(to_unsigned(142,8) ,
22211	 => std_logic_vector(to_unsigned(133,8) ,
22212	 => std_logic_vector(to_unsigned(138,8) ,
22213	 => std_logic_vector(to_unsigned(146,8) ,
22214	 => std_logic_vector(to_unsigned(147,8) ,
22215	 => std_logic_vector(to_unsigned(149,8) ,
22216	 => std_logic_vector(to_unsigned(147,8) ,
22217	 => std_logic_vector(to_unsigned(147,8) ,
22218	 => std_logic_vector(to_unsigned(146,8) ,
22219	 => std_logic_vector(to_unsigned(144,8) ,
22220	 => std_logic_vector(to_unsigned(60,8) ,
22221	 => std_logic_vector(to_unsigned(9,8) ,
22222	 => std_logic_vector(to_unsigned(2,8) ,
22223	 => std_logic_vector(to_unsigned(4,8) ,
22224	 => std_logic_vector(to_unsigned(19,8) ,
22225	 => std_logic_vector(to_unsigned(31,8) ,
22226	 => std_logic_vector(to_unsigned(35,8) ,
22227	 => std_logic_vector(to_unsigned(43,8) ,
22228	 => std_logic_vector(to_unsigned(62,8) ,
22229	 => std_logic_vector(to_unsigned(64,8) ,
22230	 => std_logic_vector(to_unsigned(55,8) ,
22231	 => std_logic_vector(to_unsigned(16,8) ,
22232	 => std_logic_vector(to_unsigned(3,8) ,
22233	 => std_logic_vector(to_unsigned(39,8) ,
22234	 => std_logic_vector(to_unsigned(152,8) ,
22235	 => std_logic_vector(to_unsigned(142,8) ,
22236	 => std_logic_vector(to_unsigned(157,8) ,
22237	 => std_logic_vector(to_unsigned(159,8) ,
22238	 => std_logic_vector(to_unsigned(157,8) ,
22239	 => std_logic_vector(to_unsigned(161,8) ,
22240	 => std_logic_vector(to_unsigned(134,8) ,
22241	 => std_logic_vector(to_unsigned(95,8) ,
22242	 => std_logic_vector(to_unsigned(91,8) ,
22243	 => std_logic_vector(to_unsigned(93,8) ,
22244	 => std_logic_vector(to_unsigned(107,8) ,
22245	 => std_logic_vector(to_unsigned(38,8) ,
22246	 => std_logic_vector(to_unsigned(3,8) ,
22247	 => std_logic_vector(to_unsigned(3,8) ,
22248	 => std_logic_vector(to_unsigned(3,8) ,
22249	 => std_logic_vector(to_unsigned(4,8) ,
22250	 => std_logic_vector(to_unsigned(5,8) ,
22251	 => std_logic_vector(to_unsigned(6,8) ,
22252	 => std_logic_vector(to_unsigned(10,8) ,
22253	 => std_logic_vector(to_unsigned(6,8) ,
22254	 => std_logic_vector(to_unsigned(3,8) ,
22255	 => std_logic_vector(to_unsigned(11,8) ,
22256	 => std_logic_vector(to_unsigned(29,8) ,
22257	 => std_logic_vector(to_unsigned(36,8) ,
22258	 => std_logic_vector(to_unsigned(46,8) ,
22259	 => std_logic_vector(to_unsigned(60,8) ,
22260	 => std_logic_vector(to_unsigned(91,8) ,
22261	 => std_logic_vector(to_unsigned(115,8) ,
22262	 => std_logic_vector(to_unsigned(124,8) ,
22263	 => std_logic_vector(to_unsigned(138,8) ,
22264	 => std_logic_vector(to_unsigned(125,8) ,
22265	 => std_logic_vector(to_unsigned(111,8) ,
22266	 => std_logic_vector(to_unsigned(93,8) ,
22267	 => std_logic_vector(to_unsigned(96,8) ,
22268	 => std_logic_vector(to_unsigned(107,8) ,
22269	 => std_logic_vector(to_unsigned(114,8) ,
22270	 => std_logic_vector(to_unsigned(114,8) ,
22271	 => std_logic_vector(to_unsigned(127,8) ,
22272	 => std_logic_vector(to_unsigned(70,8) ,
22273	 => std_logic_vector(to_unsigned(2,8) ,
22274	 => std_logic_vector(to_unsigned(0,8) ,
22275	 => std_logic_vector(to_unsigned(1,8) ,
22276	 => std_logic_vector(to_unsigned(1,8) ,
22277	 => std_logic_vector(to_unsigned(1,8) ,
22278	 => std_logic_vector(to_unsigned(1,8) ,
22279	 => std_logic_vector(to_unsigned(3,8) ,
22280	 => std_logic_vector(to_unsigned(3,8) ,
22281	 => std_logic_vector(to_unsigned(1,8) ,
22282	 => std_logic_vector(to_unsigned(2,8) ,
22283	 => std_logic_vector(to_unsigned(3,8) ,
22284	 => std_logic_vector(to_unsigned(2,8) ,
22285	 => std_logic_vector(to_unsigned(7,8) ,
22286	 => std_logic_vector(to_unsigned(46,8) ,
22287	 => std_logic_vector(to_unsigned(141,8) ,
22288	 => std_logic_vector(to_unsigned(124,8) ,
22289	 => std_logic_vector(to_unsigned(124,8) ,
22290	 => std_logic_vector(to_unsigned(121,8) ,
22291	 => std_logic_vector(to_unsigned(116,8) ,
22292	 => std_logic_vector(to_unsigned(119,8) ,
22293	 => std_logic_vector(to_unsigned(124,8) ,
22294	 => std_logic_vector(to_unsigned(118,8) ,
22295	 => std_logic_vector(to_unsigned(118,8) ,
22296	 => std_logic_vector(to_unsigned(124,8) ,
22297	 => std_logic_vector(to_unsigned(125,8) ,
22298	 => std_logic_vector(to_unsigned(122,8) ,
22299	 => std_logic_vector(to_unsigned(125,8) ,
22300	 => std_logic_vector(to_unsigned(130,8) ,
22301	 => std_logic_vector(to_unsigned(127,8) ,
22302	 => std_logic_vector(to_unsigned(134,8) ,
22303	 => std_logic_vector(to_unsigned(33,8) ,
22304	 => std_logic_vector(to_unsigned(3,8) ,
22305	 => std_logic_vector(to_unsigned(3,8) ,
22306	 => std_logic_vector(to_unsigned(3,8) ,
22307	 => std_logic_vector(to_unsigned(8,8) ,
22308	 => std_logic_vector(to_unsigned(19,8) ,
22309	 => std_logic_vector(to_unsigned(14,8) ,
22310	 => std_logic_vector(to_unsigned(7,8) ,
22311	 => std_logic_vector(to_unsigned(3,8) ,
22312	 => std_logic_vector(to_unsigned(2,8) ,
22313	 => std_logic_vector(to_unsigned(6,8) ,
22314	 => std_logic_vector(to_unsigned(13,8) ,
22315	 => std_logic_vector(to_unsigned(14,8) ,
22316	 => std_logic_vector(to_unsigned(44,8) ,
22317	 => std_logic_vector(to_unsigned(58,8) ,
22318	 => std_logic_vector(to_unsigned(78,8) ,
22319	 => std_logic_vector(to_unsigned(136,8) ,
22320	 => std_logic_vector(to_unsigned(136,8) ,
22321	 => std_logic_vector(to_unsigned(133,8) ,
22322	 => std_logic_vector(to_unsigned(138,8) ,
22323	 => std_logic_vector(to_unsigned(138,8) ,
22324	 => std_logic_vector(to_unsigned(127,8) ,
22325	 => std_logic_vector(to_unsigned(133,8) ,
22326	 => std_logic_vector(to_unsigned(144,8) ,
22327	 => std_logic_vector(to_unsigned(142,8) ,
22328	 => std_logic_vector(to_unsigned(152,8) ,
22329	 => std_logic_vector(to_unsigned(157,8) ,
22330	 => std_logic_vector(to_unsigned(147,8) ,
22331	 => std_logic_vector(to_unsigned(146,8) ,
22332	 => std_logic_vector(to_unsigned(157,8) ,
22333	 => std_logic_vector(to_unsigned(25,8) ,
22334	 => std_logic_vector(to_unsigned(1,8) ,
22335	 => std_logic_vector(to_unsigned(3,8) ,
22336	 => std_logic_vector(to_unsigned(84,8) ,
22337	 => std_logic_vector(to_unsigned(179,8) ,
22338	 => std_logic_vector(to_unsigned(144,8) ,
22339	 => std_logic_vector(to_unsigned(157,8) ,
22340	 => std_logic_vector(to_unsigned(159,8) ,
22341	 => std_logic_vector(to_unsigned(161,8) ,
22342	 => std_logic_vector(to_unsigned(151,8) ,
22343	 => std_logic_vector(to_unsigned(154,8) ,
22344	 => std_logic_vector(to_unsigned(152,8) ,
22345	 => std_logic_vector(to_unsigned(152,8) ,
22346	 => std_logic_vector(to_unsigned(156,8) ,
22347	 => std_logic_vector(to_unsigned(163,8) ,
22348	 => std_logic_vector(to_unsigned(159,8) ,
22349	 => std_logic_vector(to_unsigned(142,8) ,
22350	 => std_logic_vector(to_unsigned(125,8) ,
22351	 => std_logic_vector(to_unsigned(116,8) ,
22352	 => std_logic_vector(to_unsigned(122,8) ,
22353	 => std_logic_vector(to_unsigned(147,8) ,
22354	 => std_logic_vector(to_unsigned(141,8) ,
22355	 => std_logic_vector(to_unsigned(45,8) ,
22356	 => std_logic_vector(to_unsigned(4,8) ,
22357	 => std_logic_vector(to_unsigned(3,8) ,
22358	 => std_logic_vector(to_unsigned(1,8) ,
22359	 => std_logic_vector(to_unsigned(3,8) ,
22360	 => std_logic_vector(to_unsigned(6,8) ,
22361	 => std_logic_vector(to_unsigned(1,8) ,
22362	 => std_logic_vector(to_unsigned(1,8) ,
22363	 => std_logic_vector(to_unsigned(6,8) ,
22364	 => std_logic_vector(to_unsigned(33,8) ,
22365	 => std_logic_vector(to_unsigned(31,8) ,
22366	 => std_logic_vector(to_unsigned(14,8) ,
22367	 => std_logic_vector(to_unsigned(8,8) ,
22368	 => std_logic_vector(to_unsigned(55,8) ,
22369	 => std_logic_vector(to_unsigned(111,8) ,
22370	 => std_logic_vector(to_unsigned(109,8) ,
22371	 => std_logic_vector(to_unsigned(119,8) ,
22372	 => std_logic_vector(to_unsigned(107,8) ,
22373	 => std_logic_vector(to_unsigned(86,8) ,
22374	 => std_logic_vector(to_unsigned(85,8) ,
22375	 => std_logic_vector(to_unsigned(104,8) ,
22376	 => std_logic_vector(to_unsigned(138,8) ,
22377	 => std_logic_vector(to_unsigned(109,8) ,
22378	 => std_logic_vector(to_unsigned(92,8) ,
22379	 => std_logic_vector(to_unsigned(90,8) ,
22380	 => std_logic_vector(to_unsigned(105,8) ,
22381	 => std_logic_vector(to_unsigned(107,8) ,
22382	 => std_logic_vector(to_unsigned(131,8) ,
22383	 => std_logic_vector(to_unsigned(156,8) ,
22384	 => std_logic_vector(to_unsigned(124,8) ,
22385	 => std_logic_vector(to_unsigned(104,8) ,
22386	 => std_logic_vector(to_unsigned(115,8) ,
22387	 => std_logic_vector(to_unsigned(157,8) ,
22388	 => std_logic_vector(to_unsigned(154,8) ,
22389	 => std_logic_vector(to_unsigned(157,8) ,
22390	 => std_logic_vector(to_unsigned(159,8) ,
22391	 => std_logic_vector(to_unsigned(118,8) ,
22392	 => std_logic_vector(to_unsigned(119,8) ,
22393	 => std_logic_vector(to_unsigned(139,8) ,
22394	 => std_logic_vector(to_unsigned(119,8) ,
22395	 => std_logic_vector(to_unsigned(100,8) ,
22396	 => std_logic_vector(to_unsigned(100,8) ,
22397	 => std_logic_vector(to_unsigned(111,8) ,
22398	 => std_logic_vector(to_unsigned(103,8) ,
22399	 => std_logic_vector(to_unsigned(119,8) ,
22400	 => std_logic_vector(to_unsigned(147,8) ,
22401	 => std_logic_vector(to_unsigned(154,8) ,
22402	 => std_logic_vector(to_unsigned(154,8) ,
22403	 => std_logic_vector(to_unsigned(156,8) ,
22404	 => std_logic_vector(to_unsigned(159,8) ,
22405	 => std_logic_vector(to_unsigned(157,8) ,
22406	 => std_logic_vector(to_unsigned(157,8) ,
22407	 => std_logic_vector(to_unsigned(163,8) ,
22408	 => std_logic_vector(to_unsigned(111,8) ,
22409	 => std_logic_vector(to_unsigned(52,8) ,
22410	 => std_logic_vector(to_unsigned(41,8) ,
22411	 => std_logic_vector(to_unsigned(42,8) ,
22412	 => std_logic_vector(to_unsigned(38,8) ,
22413	 => std_logic_vector(to_unsigned(20,8) ,
22414	 => std_logic_vector(to_unsigned(14,8) ,
22415	 => std_logic_vector(to_unsigned(37,8) ,
22416	 => std_logic_vector(to_unsigned(17,8) ,
22417	 => std_logic_vector(to_unsigned(4,8) ,
22418	 => std_logic_vector(to_unsigned(8,8) ,
22419	 => std_logic_vector(to_unsigned(12,8) ,
22420	 => std_logic_vector(to_unsigned(41,8) ,
22421	 => std_logic_vector(to_unsigned(30,8) ,
22422	 => std_logic_vector(to_unsigned(5,8) ,
22423	 => std_logic_vector(to_unsigned(2,8) ,
22424	 => std_logic_vector(to_unsigned(3,8) ,
22425	 => std_logic_vector(to_unsigned(8,8) ,
22426	 => std_logic_vector(to_unsigned(4,8) ,
22427	 => std_logic_vector(to_unsigned(2,8) ,
22428	 => std_logic_vector(to_unsigned(2,8) ,
22429	 => std_logic_vector(to_unsigned(6,8) ,
22430	 => std_logic_vector(to_unsigned(7,8) ,
22431	 => std_logic_vector(to_unsigned(9,8) ,
22432	 => std_logic_vector(to_unsigned(7,8) ,
22433	 => std_logic_vector(to_unsigned(3,8) ,
22434	 => std_logic_vector(to_unsigned(2,8) ,
22435	 => std_logic_vector(to_unsigned(3,8) ,
22436	 => std_logic_vector(to_unsigned(7,8) ,
22437	 => std_logic_vector(to_unsigned(15,8) ,
22438	 => std_logic_vector(to_unsigned(43,8) ,
22439	 => std_logic_vector(to_unsigned(59,8) ,
22440	 => std_logic_vector(to_unsigned(16,8) ,
22441	 => std_logic_vector(to_unsigned(5,8) ,
22442	 => std_logic_vector(to_unsigned(14,8) ,
22443	 => std_logic_vector(to_unsigned(15,8) ,
22444	 => std_logic_vector(to_unsigned(37,8) ,
22445	 => std_logic_vector(to_unsigned(46,8) ,
22446	 => std_logic_vector(to_unsigned(37,8) ,
22447	 => std_logic_vector(to_unsigned(36,8) ,
22448	 => std_logic_vector(to_unsigned(39,8) ,
22449	 => std_logic_vector(to_unsigned(24,8) ,
22450	 => std_logic_vector(to_unsigned(58,8) ,
22451	 => std_logic_vector(to_unsigned(161,8) ,
22452	 => std_logic_vector(to_unsigned(173,8) ,
22453	 => std_logic_vector(to_unsigned(163,8) ,
22454	 => std_logic_vector(to_unsigned(45,8) ,
22455	 => std_logic_vector(to_unsigned(5,8) ,
22456	 => std_logic_vector(to_unsigned(36,8) ,
22457	 => std_logic_vector(to_unsigned(177,8) ,
22458	 => std_logic_vector(to_unsigned(156,8) ,
22459	 => std_logic_vector(to_unsigned(43,8) ,
22460	 => std_logic_vector(to_unsigned(20,8) ,
22461	 => std_logic_vector(to_unsigned(24,8) ,
22462	 => std_logic_vector(to_unsigned(10,8) ,
22463	 => std_logic_vector(to_unsigned(12,8) ,
22464	 => std_logic_vector(to_unsigned(11,8) ,
22465	 => std_logic_vector(to_unsigned(29,8) ,
22466	 => std_logic_vector(to_unsigned(28,8) ,
22467	 => std_logic_vector(to_unsigned(2,8) ,
22468	 => std_logic_vector(to_unsigned(2,8) ,
22469	 => std_logic_vector(to_unsigned(3,8) ,
22470	 => std_logic_vector(to_unsigned(6,8) ,
22471	 => std_logic_vector(to_unsigned(69,8) ,
22472	 => std_logic_vector(to_unsigned(154,8) ,
22473	 => std_logic_vector(to_unsigned(152,8) ,
22474	 => std_logic_vector(to_unsigned(105,8) ,
22475	 => std_logic_vector(to_unsigned(80,8) ,
22476	 => std_logic_vector(to_unsigned(112,8) ,
22477	 => std_logic_vector(to_unsigned(119,8) ,
22478	 => std_logic_vector(to_unsigned(138,8) ,
22479	 => std_logic_vector(to_unsigned(146,8) ,
22480	 => std_logic_vector(to_unsigned(156,8) ,
22481	 => std_logic_vector(to_unsigned(152,8) ,
22482	 => std_logic_vector(to_unsigned(68,8) ,
22483	 => std_logic_vector(to_unsigned(97,8) ,
22484	 => std_logic_vector(to_unsigned(175,8) ,
22485	 => std_logic_vector(to_unsigned(166,8) ,
22486	 => std_logic_vector(to_unsigned(159,8) ,
22487	 => std_logic_vector(to_unsigned(164,8) ,
22488	 => std_logic_vector(to_unsigned(154,8) ,
22489	 => std_logic_vector(to_unsigned(164,8) ,
22490	 => std_logic_vector(to_unsigned(156,8) ,
22491	 => std_logic_vector(to_unsigned(134,8) ,
22492	 => std_logic_vector(to_unsigned(154,8) ,
22493	 => std_logic_vector(to_unsigned(173,8) ,
22494	 => std_logic_vector(to_unsigned(177,8) ,
22495	 => std_logic_vector(to_unsigned(105,8) ,
22496	 => std_logic_vector(to_unsigned(26,8) ,
22497	 => std_logic_vector(to_unsigned(108,8) ,
22498	 => std_logic_vector(to_unsigned(73,8) ,
22499	 => std_logic_vector(to_unsigned(73,8) ,
22500	 => std_logic_vector(to_unsigned(146,8) ,
22501	 => std_logic_vector(to_unsigned(163,8) ,
22502	 => std_logic_vector(to_unsigned(166,8) ,
22503	 => std_logic_vector(to_unsigned(166,8) ,
22504	 => std_logic_vector(to_unsigned(159,8) ,
22505	 => std_logic_vector(to_unsigned(157,8) ,
22506	 => std_logic_vector(to_unsigned(166,8) ,
22507	 => std_logic_vector(to_unsigned(168,8) ,
22508	 => std_logic_vector(to_unsigned(170,8) ,
22509	 => std_logic_vector(to_unsigned(171,8) ,
22510	 => std_logic_vector(to_unsigned(164,8) ,
22511	 => std_logic_vector(to_unsigned(152,8) ,
22512	 => std_logic_vector(to_unsigned(149,8) ,
22513	 => std_logic_vector(to_unsigned(170,8) ,
22514	 => std_logic_vector(to_unsigned(134,8) ,
22515	 => std_logic_vector(to_unsigned(29,8) ,
22516	 => std_logic_vector(to_unsigned(24,8) ,
22517	 => std_logic_vector(to_unsigned(43,8) ,
22518	 => std_logic_vector(to_unsigned(33,8) ,
22519	 => std_logic_vector(to_unsigned(29,8) ,
22520	 => std_logic_vector(to_unsigned(51,8) ,
22521	 => std_logic_vector(to_unsigned(34,8) ,
22522	 => std_logic_vector(to_unsigned(18,8) ,
22523	 => std_logic_vector(to_unsigned(18,8) ,
22524	 => std_logic_vector(to_unsigned(18,8) ,
22525	 => std_logic_vector(to_unsigned(27,8) ,
22526	 => std_logic_vector(to_unsigned(37,8) ,
22527	 => std_logic_vector(to_unsigned(95,8) ,
22528	 => std_logic_vector(to_unsigned(166,8) ,
22529	 => std_logic_vector(to_unsigned(161,8) ,
22530	 => std_logic_vector(to_unsigned(147,8) ,
22531	 => std_logic_vector(to_unsigned(128,8) ,
22532	 => std_logic_vector(to_unsigned(139,8) ,
22533	 => std_logic_vector(to_unsigned(151,8) ,
22534	 => std_logic_vector(to_unsigned(147,8) ,
22535	 => std_logic_vector(to_unsigned(149,8) ,
22536	 => std_logic_vector(to_unsigned(149,8) ,
22537	 => std_logic_vector(to_unsigned(152,8) ,
22538	 => std_logic_vector(to_unsigned(142,8) ,
22539	 => std_logic_vector(to_unsigned(133,8) ,
22540	 => std_logic_vector(to_unsigned(146,8) ,
22541	 => std_logic_vector(to_unsigned(107,8) ,
22542	 => std_logic_vector(to_unsigned(70,8) ,
22543	 => std_logic_vector(to_unsigned(22,8) ,
22544	 => std_logic_vector(to_unsigned(2,8) ,
22545	 => std_logic_vector(to_unsigned(3,8) ,
22546	 => std_logic_vector(to_unsigned(4,8) ,
22547	 => std_logic_vector(to_unsigned(3,8) ,
22548	 => std_logic_vector(to_unsigned(4,8) ,
22549	 => std_logic_vector(to_unsigned(3,8) ,
22550	 => std_logic_vector(to_unsigned(8,8) ,
22551	 => std_logic_vector(to_unsigned(12,8) ,
22552	 => std_logic_vector(to_unsigned(19,8) ,
22553	 => std_logic_vector(to_unsigned(119,8) ,
22554	 => std_logic_vector(to_unsigned(171,8) ,
22555	 => std_logic_vector(to_unsigned(157,8) ,
22556	 => std_logic_vector(to_unsigned(159,8) ,
22557	 => std_logic_vector(to_unsigned(157,8) ,
22558	 => std_logic_vector(to_unsigned(157,8) ,
22559	 => std_logic_vector(to_unsigned(163,8) ,
22560	 => std_logic_vector(to_unsigned(134,8) ,
22561	 => std_logic_vector(to_unsigned(105,8) ,
22562	 => std_logic_vector(to_unsigned(112,8) ,
22563	 => std_logic_vector(to_unsigned(105,8) ,
22564	 => std_logic_vector(to_unsigned(118,8) ,
22565	 => std_logic_vector(to_unsigned(109,8) ,
22566	 => std_logic_vector(to_unsigned(10,8) ,
22567	 => std_logic_vector(to_unsigned(1,8) ,
22568	 => std_logic_vector(to_unsigned(3,8) ,
22569	 => std_logic_vector(to_unsigned(7,8) ,
22570	 => std_logic_vector(to_unsigned(5,8) ,
22571	 => std_logic_vector(to_unsigned(4,8) ,
22572	 => std_logic_vector(to_unsigned(5,8) ,
22573	 => std_logic_vector(to_unsigned(3,8) ,
22574	 => std_logic_vector(to_unsigned(5,8) ,
22575	 => std_logic_vector(to_unsigned(11,8) ,
22576	 => std_logic_vector(to_unsigned(19,8) ,
22577	 => std_logic_vector(to_unsigned(16,8) ,
22578	 => std_logic_vector(to_unsigned(11,8) ,
22579	 => std_logic_vector(to_unsigned(16,8) ,
22580	 => std_logic_vector(to_unsigned(32,8) ,
22581	 => std_logic_vector(to_unsigned(59,8) ,
22582	 => std_logic_vector(to_unsigned(109,8) ,
22583	 => std_logic_vector(to_unsigned(141,8) ,
22584	 => std_logic_vector(to_unsigned(125,8) ,
22585	 => std_logic_vector(to_unsigned(114,8) ,
22586	 => std_logic_vector(to_unsigned(95,8) ,
22587	 => std_logic_vector(to_unsigned(103,8) ,
22588	 => std_logic_vector(to_unsigned(127,8) ,
22589	 => std_logic_vector(to_unsigned(130,8) ,
22590	 => std_logic_vector(to_unsigned(121,8) ,
22591	 => std_logic_vector(to_unsigned(127,8) ,
22592	 => std_logic_vector(to_unsigned(58,8) ,
22593	 => std_logic_vector(to_unsigned(1,8) ,
22594	 => std_logic_vector(to_unsigned(0,8) ,
22595	 => std_logic_vector(to_unsigned(0,8) ,
22596	 => std_logic_vector(to_unsigned(1,8) ,
22597	 => std_logic_vector(to_unsigned(1,8) ,
22598	 => std_logic_vector(to_unsigned(1,8) ,
22599	 => std_logic_vector(to_unsigned(2,8) ,
22600	 => std_logic_vector(to_unsigned(1,8) ,
22601	 => std_logic_vector(to_unsigned(1,8) ,
22602	 => std_logic_vector(to_unsigned(3,8) ,
22603	 => std_logic_vector(to_unsigned(3,8) ,
22604	 => std_logic_vector(to_unsigned(3,8) ,
22605	 => std_logic_vector(to_unsigned(2,8) ,
22606	 => std_logic_vector(to_unsigned(48,8) ,
22607	 => std_logic_vector(to_unsigned(152,8) ,
22608	 => std_logic_vector(to_unsigned(133,8) ,
22609	 => std_logic_vector(to_unsigned(128,8) ,
22610	 => std_logic_vector(to_unsigned(130,8) ,
22611	 => std_logic_vector(to_unsigned(134,8) ,
22612	 => std_logic_vector(to_unsigned(134,8) ,
22613	 => std_logic_vector(to_unsigned(133,8) ,
22614	 => std_logic_vector(to_unsigned(133,8) ,
22615	 => std_logic_vector(to_unsigned(130,8) ,
22616	 => std_logic_vector(to_unsigned(128,8) ,
22617	 => std_logic_vector(to_unsigned(131,8) ,
22618	 => std_logic_vector(to_unsigned(131,8) ,
22619	 => std_logic_vector(to_unsigned(130,8) ,
22620	 => std_logic_vector(to_unsigned(124,8) ,
22621	 => std_logic_vector(to_unsigned(130,8) ,
22622	 => std_logic_vector(to_unsigned(134,8) ,
22623	 => std_logic_vector(to_unsigned(26,8) ,
22624	 => std_logic_vector(to_unsigned(3,8) ,
22625	 => std_logic_vector(to_unsigned(6,8) ,
22626	 => std_logic_vector(to_unsigned(3,8) ,
22627	 => std_logic_vector(to_unsigned(2,8) ,
22628	 => std_logic_vector(to_unsigned(2,8) ,
22629	 => std_logic_vector(to_unsigned(7,8) ,
22630	 => std_logic_vector(to_unsigned(7,8) ,
22631	 => std_logic_vector(to_unsigned(2,8) ,
22632	 => std_logic_vector(to_unsigned(2,8) ,
22633	 => std_logic_vector(to_unsigned(2,8) ,
22634	 => std_logic_vector(to_unsigned(3,8) ,
22635	 => std_logic_vector(to_unsigned(4,8) ,
22636	 => std_logic_vector(to_unsigned(9,8) ,
22637	 => std_logic_vector(to_unsigned(10,8) ,
22638	 => std_logic_vector(to_unsigned(57,8) ,
22639	 => std_logic_vector(to_unsigned(147,8) ,
22640	 => std_logic_vector(to_unsigned(134,8) ,
22641	 => std_logic_vector(to_unsigned(144,8) ,
22642	 => std_logic_vector(to_unsigned(146,8) ,
22643	 => std_logic_vector(to_unsigned(142,8) ,
22644	 => std_logic_vector(to_unsigned(142,8) ,
22645	 => std_logic_vector(to_unsigned(144,8) ,
22646	 => std_logic_vector(to_unsigned(141,8) ,
22647	 => std_logic_vector(to_unsigned(144,8) ,
22648	 => std_logic_vector(to_unsigned(151,8) ,
22649	 => std_logic_vector(to_unsigned(159,8) ,
22650	 => std_logic_vector(to_unsigned(157,8) ,
22651	 => std_logic_vector(to_unsigned(147,8) ,
22652	 => std_logic_vector(to_unsigned(163,8) ,
22653	 => std_logic_vector(to_unsigned(46,8) ,
22654	 => std_logic_vector(to_unsigned(1,8) ,
22655	 => std_logic_vector(to_unsigned(2,8) ,
22656	 => std_logic_vector(to_unsigned(36,8) ,
22657	 => std_logic_vector(to_unsigned(104,8) ,
22658	 => std_logic_vector(to_unsigned(96,8) ,
22659	 => std_logic_vector(to_unsigned(157,8) ,
22660	 => std_logic_vector(to_unsigned(157,8) ,
22661	 => std_logic_vector(to_unsigned(161,8) ,
22662	 => std_logic_vector(to_unsigned(156,8) ,
22663	 => std_logic_vector(to_unsigned(154,8) ,
22664	 => std_logic_vector(to_unsigned(151,8) ,
22665	 => std_logic_vector(to_unsigned(147,8) ,
22666	 => std_logic_vector(to_unsigned(152,8) ,
22667	 => std_logic_vector(to_unsigned(161,8) ,
22668	 => std_logic_vector(to_unsigned(157,8) ,
22669	 => std_logic_vector(to_unsigned(141,8) ,
22670	 => std_logic_vector(to_unsigned(136,8) ,
22671	 => std_logic_vector(to_unsigned(138,8) ,
22672	 => std_logic_vector(to_unsigned(133,8) ,
22673	 => std_logic_vector(to_unsigned(125,8) ,
22674	 => std_logic_vector(to_unsigned(130,8) ,
22675	 => std_logic_vector(to_unsigned(100,8) ,
22676	 => std_logic_vector(to_unsigned(9,8) ,
22677	 => std_logic_vector(to_unsigned(2,8) ,
22678	 => std_logic_vector(to_unsigned(2,8) ,
22679	 => std_logic_vector(to_unsigned(6,8) ,
22680	 => std_logic_vector(to_unsigned(27,8) ,
22681	 => std_logic_vector(to_unsigned(18,8) ,
22682	 => std_logic_vector(to_unsigned(27,8) ,
22683	 => std_logic_vector(to_unsigned(31,8) ,
22684	 => std_logic_vector(to_unsigned(30,8) ,
22685	 => std_logic_vector(to_unsigned(12,8) ,
22686	 => std_logic_vector(to_unsigned(10,8) ,
22687	 => std_logic_vector(to_unsigned(24,8) ,
22688	 => std_logic_vector(to_unsigned(78,8) ,
22689	 => std_logic_vector(to_unsigned(99,8) ,
22690	 => std_logic_vector(to_unsigned(101,8) ,
22691	 => std_logic_vector(to_unsigned(104,8) ,
22692	 => std_logic_vector(to_unsigned(99,8) ,
22693	 => std_logic_vector(to_unsigned(91,8) ,
22694	 => std_logic_vector(to_unsigned(88,8) ,
22695	 => std_logic_vector(to_unsigned(109,8) ,
22696	 => std_logic_vector(to_unsigned(134,8) ,
22697	 => std_logic_vector(to_unsigned(109,8) ,
22698	 => std_logic_vector(to_unsigned(103,8) ,
22699	 => std_logic_vector(to_unsigned(87,8) ,
22700	 => std_logic_vector(to_unsigned(108,8) ,
22701	 => std_logic_vector(to_unsigned(136,8) ,
22702	 => std_logic_vector(to_unsigned(118,8) ,
22703	 => std_logic_vector(to_unsigned(121,8) ,
22704	 => std_logic_vector(to_unsigned(134,8) ,
22705	 => std_logic_vector(to_unsigned(136,8) ,
22706	 => std_logic_vector(to_unsigned(116,8) ,
22707	 => std_logic_vector(to_unsigned(125,8) ,
22708	 => std_logic_vector(to_unsigned(159,8) ,
22709	 => std_logic_vector(to_unsigned(159,8) ,
22710	 => std_logic_vector(to_unsigned(161,8) ,
22711	 => std_logic_vector(to_unsigned(154,8) ,
22712	 => std_logic_vector(to_unsigned(133,8) ,
22713	 => std_logic_vector(to_unsigned(121,8) ,
22714	 => std_logic_vector(to_unsigned(122,8) ,
22715	 => std_logic_vector(to_unsigned(124,8) ,
22716	 => std_logic_vector(to_unsigned(125,8) ,
22717	 => std_logic_vector(to_unsigned(111,8) ,
22718	 => std_logic_vector(to_unsigned(109,8) ,
22719	 => std_logic_vector(to_unsigned(131,8) ,
22720	 => std_logic_vector(to_unsigned(146,8) ,
22721	 => std_logic_vector(to_unsigned(154,8) ,
22722	 => std_logic_vector(to_unsigned(156,8) ,
22723	 => std_logic_vector(to_unsigned(157,8) ,
22724	 => std_logic_vector(to_unsigned(159,8) ,
22725	 => std_logic_vector(to_unsigned(156,8) ,
22726	 => std_logic_vector(to_unsigned(156,8) ,
22727	 => std_logic_vector(to_unsigned(156,8) ,
22728	 => std_logic_vector(to_unsigned(84,8) ,
22729	 => std_logic_vector(to_unsigned(37,8) ,
22730	 => std_logic_vector(to_unsigned(30,8) ,
22731	 => std_logic_vector(to_unsigned(30,8) ,
22732	 => std_logic_vector(to_unsigned(24,8) ,
22733	 => std_logic_vector(to_unsigned(23,8) ,
22734	 => std_logic_vector(to_unsigned(37,8) ,
22735	 => std_logic_vector(to_unsigned(43,8) ,
22736	 => std_logic_vector(to_unsigned(4,8) ,
22737	 => std_logic_vector(to_unsigned(1,8) ,
22738	 => std_logic_vector(to_unsigned(3,8) ,
22739	 => std_logic_vector(to_unsigned(5,8) ,
22740	 => std_logic_vector(to_unsigned(20,8) ,
22741	 => std_logic_vector(to_unsigned(17,8) ,
22742	 => std_logic_vector(to_unsigned(4,8) ,
22743	 => std_logic_vector(to_unsigned(3,8) ,
22744	 => std_logic_vector(to_unsigned(1,8) ,
22745	 => std_logic_vector(to_unsigned(10,8) ,
22746	 => std_logic_vector(to_unsigned(11,8) ,
22747	 => std_logic_vector(to_unsigned(3,8) ,
22748	 => std_logic_vector(to_unsigned(3,8) ,
22749	 => std_logic_vector(to_unsigned(3,8) ,
22750	 => std_logic_vector(to_unsigned(5,8) ,
22751	 => std_logic_vector(to_unsigned(7,8) ,
22752	 => std_logic_vector(to_unsigned(3,8) ,
22753	 => std_logic_vector(to_unsigned(1,8) ,
22754	 => std_logic_vector(to_unsigned(1,8) ,
22755	 => std_logic_vector(to_unsigned(1,8) ,
22756	 => std_logic_vector(to_unsigned(8,8) ,
22757	 => std_logic_vector(to_unsigned(7,8) ,
22758	 => std_logic_vector(to_unsigned(6,8) ,
22759	 => std_logic_vector(to_unsigned(25,8) ,
22760	 => std_logic_vector(to_unsigned(7,8) ,
22761	 => std_logic_vector(to_unsigned(6,8) ,
22762	 => std_logic_vector(to_unsigned(10,8) ,
22763	 => std_logic_vector(to_unsigned(26,8) ,
22764	 => std_logic_vector(to_unsigned(46,8) ,
22765	 => std_logic_vector(to_unsigned(31,8) ,
22766	 => std_logic_vector(to_unsigned(41,8) ,
22767	 => std_logic_vector(to_unsigned(43,8) ,
22768	 => std_logic_vector(to_unsigned(43,8) ,
22769	 => std_logic_vector(to_unsigned(27,8) ,
22770	 => std_logic_vector(to_unsigned(16,8) ,
22771	 => std_logic_vector(to_unsigned(92,8) ,
22772	 => std_logic_vector(to_unsigned(171,8) ,
22773	 => std_logic_vector(to_unsigned(179,8) ,
22774	 => std_logic_vector(to_unsigned(136,8) ,
22775	 => std_logic_vector(to_unsigned(86,8) ,
22776	 => std_logic_vector(to_unsigned(147,8) ,
22777	 => std_logic_vector(to_unsigned(151,8) ,
22778	 => std_logic_vector(to_unsigned(90,8) ,
22779	 => std_logic_vector(to_unsigned(88,8) ,
22780	 => std_logic_vector(to_unsigned(92,8) ,
22781	 => std_logic_vector(to_unsigned(91,8) ,
22782	 => std_logic_vector(to_unsigned(50,8) ,
22783	 => std_logic_vector(to_unsigned(15,8) ,
22784	 => std_logic_vector(to_unsigned(7,8) ,
22785	 => std_logic_vector(to_unsigned(4,8) ,
22786	 => std_logic_vector(to_unsigned(1,8) ,
22787	 => std_logic_vector(to_unsigned(2,8) ,
22788	 => std_logic_vector(to_unsigned(5,8) ,
22789	 => std_logic_vector(to_unsigned(4,8) ,
22790	 => std_logic_vector(to_unsigned(3,8) ,
22791	 => std_logic_vector(to_unsigned(13,8) ,
22792	 => std_logic_vector(to_unsigned(107,8) ,
22793	 => std_logic_vector(to_unsigned(164,8) ,
22794	 => std_logic_vector(to_unsigned(103,8) ,
22795	 => std_logic_vector(to_unsigned(35,8) ,
22796	 => std_logic_vector(to_unsigned(96,8) ,
22797	 => std_logic_vector(to_unsigned(133,8) ,
22798	 => std_logic_vector(to_unsigned(138,8) ,
22799	 => std_logic_vector(to_unsigned(125,8) ,
22800	 => std_logic_vector(to_unsigned(179,8) ,
22801	 => std_logic_vector(to_unsigned(100,8) ,
22802	 => std_logic_vector(to_unsigned(12,8) ,
22803	 => std_logic_vector(to_unsigned(29,8) ,
22804	 => std_logic_vector(to_unsigned(91,8) ,
22805	 => std_logic_vector(to_unsigned(170,8) ,
22806	 => std_logic_vector(to_unsigned(171,8) ,
22807	 => std_logic_vector(to_unsigned(161,8) ,
22808	 => std_logic_vector(to_unsigned(157,8) ,
22809	 => std_logic_vector(to_unsigned(166,8) ,
22810	 => std_logic_vector(to_unsigned(159,8) ,
22811	 => std_logic_vector(to_unsigned(142,8) ,
22812	 => std_logic_vector(to_unsigned(154,8) ,
22813	 => std_logic_vector(to_unsigned(164,8) ,
22814	 => std_logic_vector(to_unsigned(171,8) ,
22815	 => std_logic_vector(to_unsigned(156,8) ,
22816	 => std_logic_vector(to_unsigned(90,8) ,
22817	 => std_logic_vector(to_unsigned(154,8) ,
22818	 => std_logic_vector(to_unsigned(87,8) ,
22819	 => std_logic_vector(to_unsigned(81,8) ,
22820	 => std_logic_vector(to_unsigned(144,8) ,
22821	 => std_logic_vector(to_unsigned(170,8) ,
22822	 => std_logic_vector(to_unsigned(168,8) ,
22823	 => std_logic_vector(to_unsigned(161,8) ,
22824	 => std_logic_vector(to_unsigned(164,8) ,
22825	 => std_logic_vector(to_unsigned(164,8) ,
22826	 => std_logic_vector(to_unsigned(152,8) ,
22827	 => std_logic_vector(to_unsigned(170,8) ,
22828	 => std_logic_vector(to_unsigned(171,8) ,
22829	 => std_logic_vector(to_unsigned(161,8) ,
22830	 => std_logic_vector(to_unsigned(163,8) ,
22831	 => std_logic_vector(to_unsigned(154,8) ,
22832	 => std_logic_vector(to_unsigned(149,8) ,
22833	 => std_logic_vector(to_unsigned(157,8) ,
22834	 => std_logic_vector(to_unsigned(147,8) ,
22835	 => std_logic_vector(to_unsigned(40,8) ,
22836	 => std_logic_vector(to_unsigned(8,8) ,
22837	 => std_logic_vector(to_unsigned(3,8) ,
22838	 => std_logic_vector(to_unsigned(6,8) ,
22839	 => std_logic_vector(to_unsigned(15,8) ,
22840	 => std_logic_vector(to_unsigned(9,8) ,
22841	 => std_logic_vector(to_unsigned(8,8) ,
22842	 => std_logic_vector(to_unsigned(25,8) ,
22843	 => std_logic_vector(to_unsigned(64,8) ,
22844	 => std_logic_vector(to_unsigned(57,8) ,
22845	 => std_logic_vector(to_unsigned(28,8) ,
22846	 => std_logic_vector(to_unsigned(10,8) ,
22847	 => std_logic_vector(to_unsigned(71,8) ,
22848	 => std_logic_vector(to_unsigned(171,8) ,
22849	 => std_logic_vector(to_unsigned(157,8) ,
22850	 => std_logic_vector(to_unsigned(139,8) ,
22851	 => std_logic_vector(to_unsigned(134,8) ,
22852	 => std_logic_vector(to_unsigned(144,8) ,
22853	 => std_logic_vector(to_unsigned(151,8) ,
22854	 => std_logic_vector(to_unsigned(152,8) ,
22855	 => std_logic_vector(to_unsigned(154,8) ,
22856	 => std_logic_vector(to_unsigned(154,8) ,
22857	 => std_logic_vector(to_unsigned(152,8) ,
22858	 => std_logic_vector(to_unsigned(144,8) ,
22859	 => std_logic_vector(to_unsigned(138,8) ,
22860	 => std_logic_vector(to_unsigned(134,8) ,
22861	 => std_logic_vector(to_unsigned(154,8) ,
22862	 => std_logic_vector(to_unsigned(192,8) ,
22863	 => std_logic_vector(to_unsigned(70,8) ,
22864	 => std_logic_vector(to_unsigned(1,8) ,
22865	 => std_logic_vector(to_unsigned(1,8) ,
22866	 => std_logic_vector(to_unsigned(3,8) ,
22867	 => std_logic_vector(to_unsigned(3,8) ,
22868	 => std_logic_vector(to_unsigned(1,8) ,
22869	 => std_logic_vector(to_unsigned(2,8) ,
22870	 => std_logic_vector(to_unsigned(15,8) ,
22871	 => std_logic_vector(to_unsigned(19,8) ,
22872	 => std_logic_vector(to_unsigned(49,8) ,
22873	 => std_logic_vector(to_unsigned(168,8) ,
22874	 => std_logic_vector(to_unsigned(161,8) ,
22875	 => std_logic_vector(to_unsigned(157,8) ,
22876	 => std_logic_vector(to_unsigned(157,8) ,
22877	 => std_logic_vector(to_unsigned(156,8) ,
22878	 => std_logic_vector(to_unsigned(152,8) ,
22879	 => std_logic_vector(to_unsigned(156,8) ,
22880	 => std_logic_vector(to_unsigned(136,8) ,
22881	 => std_logic_vector(to_unsigned(114,8) ,
22882	 => std_logic_vector(to_unsigned(121,8) ,
22883	 => std_logic_vector(to_unsigned(109,8) ,
22884	 => std_logic_vector(to_unsigned(99,8) ,
22885	 => std_logic_vector(to_unsigned(116,8) ,
22886	 => std_logic_vector(to_unsigned(51,8) ,
22887	 => std_logic_vector(to_unsigned(4,8) ,
22888	 => std_logic_vector(to_unsigned(3,8) ,
22889	 => std_logic_vector(to_unsigned(5,8) ,
22890	 => std_logic_vector(to_unsigned(4,8) ,
22891	 => std_logic_vector(to_unsigned(2,8) ,
22892	 => std_logic_vector(to_unsigned(2,8) ,
22893	 => std_logic_vector(to_unsigned(3,8) ,
22894	 => std_logic_vector(to_unsigned(5,8) ,
22895	 => std_logic_vector(to_unsigned(10,8) ,
22896	 => std_logic_vector(to_unsigned(18,8) ,
22897	 => std_logic_vector(to_unsigned(30,8) ,
22898	 => std_logic_vector(to_unsigned(32,8) ,
22899	 => std_logic_vector(to_unsigned(31,8) ,
22900	 => std_logic_vector(to_unsigned(22,8) ,
22901	 => std_logic_vector(to_unsigned(16,8) ,
22902	 => std_logic_vector(to_unsigned(26,8) ,
22903	 => std_logic_vector(to_unsigned(64,8) ,
22904	 => std_logic_vector(to_unsigned(103,8) ,
22905	 => std_logic_vector(to_unsigned(115,8) ,
22906	 => std_logic_vector(to_unsigned(128,8) ,
22907	 => std_logic_vector(to_unsigned(130,8) ,
22908	 => std_logic_vector(to_unsigned(131,8) ,
22909	 => std_logic_vector(to_unsigned(121,8) ,
22910	 => std_logic_vector(to_unsigned(115,8) ,
22911	 => std_logic_vector(to_unsigned(115,8) ,
22912	 => std_logic_vector(to_unsigned(86,8) ,
22913	 => std_logic_vector(to_unsigned(6,8) ,
22914	 => std_logic_vector(to_unsigned(0,8) ,
22915	 => std_logic_vector(to_unsigned(1,8) ,
22916	 => std_logic_vector(to_unsigned(1,8) ,
22917	 => std_logic_vector(to_unsigned(1,8) ,
22918	 => std_logic_vector(to_unsigned(1,8) ,
22919	 => std_logic_vector(to_unsigned(3,8) ,
22920	 => std_logic_vector(to_unsigned(2,8) ,
22921	 => std_logic_vector(to_unsigned(2,8) ,
22922	 => std_logic_vector(to_unsigned(8,8) ,
22923	 => std_logic_vector(to_unsigned(52,8) ,
22924	 => std_logic_vector(to_unsigned(60,8) ,
22925	 => std_logic_vector(to_unsigned(17,8) ,
22926	 => std_logic_vector(to_unsigned(76,8) ,
22927	 => std_logic_vector(to_unsigned(151,8) ,
22928	 => std_logic_vector(to_unsigned(128,8) ,
22929	 => std_logic_vector(to_unsigned(136,8) ,
22930	 => std_logic_vector(to_unsigned(136,8) ,
22931	 => std_logic_vector(to_unsigned(134,8) ,
22932	 => std_logic_vector(to_unsigned(138,8) ,
22933	 => std_logic_vector(to_unsigned(134,8) ,
22934	 => std_logic_vector(to_unsigned(136,8) ,
22935	 => std_logic_vector(to_unsigned(136,8) ,
22936	 => std_logic_vector(to_unsigned(136,8) ,
22937	 => std_logic_vector(to_unsigned(139,8) ,
22938	 => std_logic_vector(to_unsigned(134,8) ,
22939	 => std_logic_vector(to_unsigned(133,8) ,
22940	 => std_logic_vector(to_unsigned(125,8) ,
22941	 => std_logic_vector(to_unsigned(134,8) ,
22942	 => std_logic_vector(to_unsigned(125,8) ,
22943	 => std_logic_vector(to_unsigned(18,8) ,
22944	 => std_logic_vector(to_unsigned(4,8) ,
22945	 => std_logic_vector(to_unsigned(8,8) ,
22946	 => std_logic_vector(to_unsigned(7,8) ,
22947	 => std_logic_vector(to_unsigned(9,8) ,
22948	 => std_logic_vector(to_unsigned(8,8) ,
22949	 => std_logic_vector(to_unsigned(4,8) ,
22950	 => std_logic_vector(to_unsigned(2,8) ,
22951	 => std_logic_vector(to_unsigned(1,8) ,
22952	 => std_logic_vector(to_unsigned(1,8) ,
22953	 => std_logic_vector(to_unsigned(2,8) ,
22954	 => std_logic_vector(to_unsigned(1,8) ,
22955	 => std_logic_vector(to_unsigned(5,8) ,
22956	 => std_logic_vector(to_unsigned(18,8) ,
22957	 => std_logic_vector(to_unsigned(33,8) ,
22958	 => std_logic_vector(to_unsigned(109,8) ,
22959	 => std_logic_vector(to_unsigned(144,8) ,
22960	 => std_logic_vector(to_unsigned(138,8) ,
22961	 => std_logic_vector(to_unsigned(134,8) ,
22962	 => std_logic_vector(to_unsigned(130,8) ,
22963	 => std_logic_vector(to_unsigned(128,8) ,
22964	 => std_logic_vector(to_unsigned(133,8) ,
22965	 => std_logic_vector(to_unsigned(147,8) ,
22966	 => std_logic_vector(to_unsigned(144,8) ,
22967	 => std_logic_vector(to_unsigned(152,8) ,
22968	 => std_logic_vector(to_unsigned(152,8) ,
22969	 => std_logic_vector(to_unsigned(152,8) ,
22970	 => std_logic_vector(to_unsigned(152,8) ,
22971	 => std_logic_vector(to_unsigned(147,8) ,
22972	 => std_logic_vector(to_unsigned(164,8) ,
22973	 => std_logic_vector(to_unsigned(78,8) ,
22974	 => std_logic_vector(to_unsigned(3,8) ,
22975	 => std_logic_vector(to_unsigned(2,8) ,
22976	 => std_logic_vector(to_unsigned(15,8) ,
22977	 => std_logic_vector(to_unsigned(71,8) ,
22978	 => std_logic_vector(to_unsigned(109,8) ,
22979	 => std_logic_vector(to_unsigned(163,8) ,
22980	 => std_logic_vector(to_unsigned(156,8) ,
22981	 => std_logic_vector(to_unsigned(152,8) ,
22982	 => std_logic_vector(to_unsigned(157,8) ,
22983	 => std_logic_vector(to_unsigned(157,8) ,
22984	 => std_logic_vector(to_unsigned(152,8) ,
22985	 => std_logic_vector(to_unsigned(151,8) ,
22986	 => std_logic_vector(to_unsigned(152,8) ,
22987	 => std_logic_vector(to_unsigned(156,8) ,
22988	 => std_logic_vector(to_unsigned(154,8) ,
22989	 => std_logic_vector(to_unsigned(146,8) ,
22990	 => std_logic_vector(to_unsigned(142,8) ,
22991	 => std_logic_vector(to_unsigned(142,8) ,
22992	 => std_logic_vector(to_unsigned(141,8) ,
22993	 => std_logic_vector(to_unsigned(136,8) ,
22994	 => std_logic_vector(to_unsigned(127,8) ,
22995	 => std_logic_vector(to_unsigned(122,8) ,
22996	 => std_logic_vector(to_unsigned(27,8) ,
22997	 => std_logic_vector(to_unsigned(5,8) ,
22998	 => std_logic_vector(to_unsigned(3,8) ,
22999	 => std_logic_vector(to_unsigned(15,8) ,
23000	 => std_logic_vector(to_unsigned(59,8) ,
23001	 => std_logic_vector(to_unsigned(22,8) ,
23002	 => std_logic_vector(to_unsigned(21,8) ,
23003	 => std_logic_vector(to_unsigned(34,8) ,
23004	 => std_logic_vector(to_unsigned(17,8) ,
23005	 => std_logic_vector(to_unsigned(9,8) ,
23006	 => std_logic_vector(to_unsigned(10,8) ,
23007	 => std_logic_vector(to_unsigned(45,8) ,
23008	 => std_logic_vector(to_unsigned(97,8) ,
23009	 => std_logic_vector(to_unsigned(99,8) ,
23010	 => std_logic_vector(to_unsigned(97,8) ,
23011	 => std_logic_vector(to_unsigned(91,8) ,
23012	 => std_logic_vector(to_unsigned(93,8) ,
23013	 => std_logic_vector(to_unsigned(97,8) ,
23014	 => std_logic_vector(to_unsigned(100,8) ,
23015	 => std_logic_vector(to_unsigned(104,8) ,
23016	 => std_logic_vector(to_unsigned(97,8) ,
23017	 => std_logic_vector(to_unsigned(101,8) ,
23018	 => std_logic_vector(to_unsigned(95,8) ,
23019	 => std_logic_vector(to_unsigned(81,8) ,
23020	 => std_logic_vector(to_unsigned(91,8) ,
23021	 => std_logic_vector(to_unsigned(139,8) ,
23022	 => std_logic_vector(to_unsigned(119,8) ,
23023	 => std_logic_vector(to_unsigned(97,8) ,
23024	 => std_logic_vector(to_unsigned(141,8) ,
23025	 => std_logic_vector(to_unsigned(164,8) ,
23026	 => std_logic_vector(to_unsigned(127,8) ,
23027	 => std_logic_vector(to_unsigned(96,8) ,
23028	 => std_logic_vector(to_unsigned(138,8) ,
23029	 => std_logic_vector(to_unsigned(164,8) ,
23030	 => std_logic_vector(to_unsigned(154,8) ,
23031	 => std_logic_vector(to_unsigned(161,8) ,
23032	 => std_logic_vector(to_unsigned(152,8) ,
23033	 => std_logic_vector(to_unsigned(115,8) ,
23034	 => std_logic_vector(to_unsigned(125,8) ,
23035	 => std_logic_vector(to_unsigned(146,8) ,
23036	 => std_logic_vector(to_unsigned(151,8) ,
23037	 => std_logic_vector(to_unsigned(109,8) ,
23038	 => std_logic_vector(to_unsigned(109,8) ,
23039	 => std_logic_vector(to_unsigned(139,8) ,
23040	 => std_logic_vector(to_unsigned(136,8) ,
23041	 => std_logic_vector(to_unsigned(157,8) ,
23042	 => std_logic_vector(to_unsigned(157,8) ,
23043	 => std_logic_vector(to_unsigned(157,8) ,
23044	 => std_logic_vector(to_unsigned(157,8) ,
23045	 => std_logic_vector(to_unsigned(157,8) ,
23046	 => std_logic_vector(to_unsigned(161,8) ,
23047	 => std_logic_vector(to_unsigned(141,8) ,
23048	 => std_logic_vector(to_unsigned(49,8) ,
23049	 => std_logic_vector(to_unsigned(45,8) ,
23050	 => std_logic_vector(to_unsigned(23,8) ,
23051	 => std_logic_vector(to_unsigned(23,8) ,
23052	 => std_logic_vector(to_unsigned(26,8) ,
23053	 => std_logic_vector(to_unsigned(18,8) ,
23054	 => std_logic_vector(to_unsigned(6,8) ,
23055	 => std_logic_vector(to_unsigned(4,8) ,
23056	 => std_logic_vector(to_unsigned(2,8) ,
23057	 => std_logic_vector(to_unsigned(1,8) ,
23058	 => std_logic_vector(to_unsigned(11,8) ,
23059	 => std_logic_vector(to_unsigned(38,8) ,
23060	 => std_logic_vector(to_unsigned(19,8) ,
23061	 => std_logic_vector(to_unsigned(11,8) ,
23062	 => std_logic_vector(to_unsigned(2,8) ,
23063	 => std_logic_vector(to_unsigned(1,8) ,
23064	 => std_logic_vector(to_unsigned(0,8) ,
23065	 => std_logic_vector(to_unsigned(3,8) ,
23066	 => std_logic_vector(to_unsigned(10,8) ,
23067	 => std_logic_vector(to_unsigned(5,8) ,
23068	 => std_logic_vector(to_unsigned(2,8) ,
23069	 => std_logic_vector(to_unsigned(3,8) ,
23070	 => std_logic_vector(to_unsigned(3,8) ,
23071	 => std_logic_vector(to_unsigned(3,8) ,
23072	 => std_logic_vector(to_unsigned(1,8) ,
23073	 => std_logic_vector(to_unsigned(4,8) ,
23074	 => std_logic_vector(to_unsigned(6,8) ,
23075	 => std_logic_vector(to_unsigned(8,8) ,
23076	 => std_logic_vector(to_unsigned(30,8) ,
23077	 => std_logic_vector(to_unsigned(19,8) ,
23078	 => std_logic_vector(to_unsigned(1,8) ,
23079	 => std_logic_vector(to_unsigned(1,8) ,
23080	 => std_logic_vector(to_unsigned(4,8) ,
23081	 => std_logic_vector(to_unsigned(12,8) ,
23082	 => std_logic_vector(to_unsigned(12,8) ,
23083	 => std_logic_vector(to_unsigned(29,8) ,
23084	 => std_logic_vector(to_unsigned(35,8) ,
23085	 => std_logic_vector(to_unsigned(26,8) ,
23086	 => std_logic_vector(to_unsigned(30,8) ,
23087	 => std_logic_vector(to_unsigned(32,8) ,
23088	 => std_logic_vector(to_unsigned(43,8) ,
23089	 => std_logic_vector(to_unsigned(31,8) ,
23090	 => std_logic_vector(to_unsigned(5,8) ,
23091	 => std_logic_vector(to_unsigned(38,8) ,
23092	 => std_logic_vector(to_unsigned(181,8) ,
23093	 => std_logic_vector(to_unsigned(164,8) ,
23094	 => std_logic_vector(to_unsigned(171,8) ,
23095	 => std_logic_vector(to_unsigned(173,8) ,
23096	 => std_logic_vector(to_unsigned(112,8) ,
23097	 => std_logic_vector(to_unsigned(22,8) ,
23098	 => std_logic_vector(to_unsigned(12,8) ,
23099	 => std_logic_vector(to_unsigned(39,8) ,
23100	 => std_logic_vector(to_unsigned(24,8) ,
23101	 => std_logic_vector(to_unsigned(11,8) ,
23102	 => std_logic_vector(to_unsigned(7,8) ,
23103	 => std_logic_vector(to_unsigned(2,8) ,
23104	 => std_logic_vector(to_unsigned(3,8) ,
23105	 => std_logic_vector(to_unsigned(4,8) ,
23106	 => std_logic_vector(to_unsigned(4,8) ,
23107	 => std_logic_vector(to_unsigned(5,8) ,
23108	 => std_logic_vector(to_unsigned(5,8) ,
23109	 => std_logic_vector(to_unsigned(4,8) ,
23110	 => std_logic_vector(to_unsigned(8,8) ,
23111	 => std_logic_vector(to_unsigned(4,8) ,
23112	 => std_logic_vector(to_unsigned(38,8) ,
23113	 => std_logic_vector(to_unsigned(146,8) ,
23114	 => std_logic_vector(to_unsigned(86,8) ,
23115	 => std_logic_vector(to_unsigned(14,8) ,
23116	 => std_logic_vector(to_unsigned(54,8) ,
23117	 => std_logic_vector(to_unsigned(115,8) ,
23118	 => std_logic_vector(to_unsigned(138,8) ,
23119	 => std_logic_vector(to_unsigned(118,8) ,
23120	 => std_logic_vector(to_unsigned(122,8) ,
23121	 => std_logic_vector(to_unsigned(30,8) ,
23122	 => std_logic_vector(to_unsigned(10,8) ,
23123	 => std_logic_vector(to_unsigned(14,8) ,
23124	 => std_logic_vector(to_unsigned(25,8) ,
23125	 => std_logic_vector(to_unsigned(86,8) ,
23126	 => std_logic_vector(to_unsigned(151,8) ,
23127	 => std_logic_vector(to_unsigned(166,8) ,
23128	 => std_logic_vector(to_unsigned(163,8) ,
23129	 => std_logic_vector(to_unsigned(147,8) ,
23130	 => std_logic_vector(to_unsigned(141,8) ,
23131	 => std_logic_vector(to_unsigned(156,8) ,
23132	 => std_logic_vector(to_unsigned(161,8) ,
23133	 => std_logic_vector(to_unsigned(168,8) ,
23134	 => std_logic_vector(to_unsigned(170,8) ,
23135	 => std_logic_vector(to_unsigned(128,8) ,
23136	 => std_logic_vector(to_unsigned(99,8) ,
23137	 => std_logic_vector(to_unsigned(156,8) ,
23138	 => std_logic_vector(to_unsigned(168,8) ,
23139	 => std_logic_vector(to_unsigned(179,8) ,
23140	 => std_logic_vector(to_unsigned(170,8) ,
23141	 => std_logic_vector(to_unsigned(168,8) ,
23142	 => std_logic_vector(to_unsigned(170,8) ,
23143	 => std_logic_vector(to_unsigned(156,8) ,
23144	 => std_logic_vector(to_unsigned(144,8) ,
23145	 => std_logic_vector(to_unsigned(144,8) ,
23146	 => std_logic_vector(to_unsigned(136,8) ,
23147	 => std_logic_vector(to_unsigned(124,8) ,
23148	 => std_logic_vector(to_unsigned(157,8) ,
23149	 => std_logic_vector(to_unsigned(163,8) ,
23150	 => std_logic_vector(to_unsigned(163,8) ,
23151	 => std_logic_vector(to_unsigned(164,8) ,
23152	 => std_logic_vector(to_unsigned(157,8) ,
23153	 => std_logic_vector(to_unsigned(154,8) ,
23154	 => std_logic_vector(to_unsigned(163,8) ,
23155	 => std_logic_vector(to_unsigned(127,8) ,
23156	 => std_logic_vector(to_unsigned(25,8) ,
23157	 => std_logic_vector(to_unsigned(2,8) ,
23158	 => std_logic_vector(to_unsigned(0,8) ,
23159	 => std_logic_vector(to_unsigned(1,8) ,
23160	 => std_logic_vector(to_unsigned(4,8) ,
23161	 => std_logic_vector(to_unsigned(6,8) ,
23162	 => std_logic_vector(to_unsigned(9,8) ,
23163	 => std_logic_vector(to_unsigned(22,8) ,
23164	 => std_logic_vector(to_unsigned(21,8) ,
23165	 => std_logic_vector(to_unsigned(16,8) ,
23166	 => std_logic_vector(to_unsigned(11,8) ,
23167	 => std_logic_vector(to_unsigned(51,8) ,
23168	 => std_logic_vector(to_unsigned(166,8) ,
23169	 => std_logic_vector(to_unsigned(161,8) ,
23170	 => std_logic_vector(to_unsigned(138,8) ,
23171	 => std_logic_vector(to_unsigned(130,8) ,
23172	 => std_logic_vector(to_unsigned(144,8) ,
23173	 => std_logic_vector(to_unsigned(149,8) ,
23174	 => std_logic_vector(to_unsigned(152,8) ,
23175	 => std_logic_vector(to_unsigned(156,8) ,
23176	 => std_logic_vector(to_unsigned(156,8) ,
23177	 => std_logic_vector(to_unsigned(154,8) ,
23178	 => std_logic_vector(to_unsigned(147,8) ,
23179	 => std_logic_vector(to_unsigned(142,8) ,
23180	 => std_logic_vector(to_unsigned(139,8) ,
23181	 => std_logic_vector(to_unsigned(139,8) ,
23182	 => std_logic_vector(to_unsigned(168,8) ,
23183	 => std_logic_vector(to_unsigned(88,8) ,
23184	 => std_logic_vector(to_unsigned(6,8) ,
23185	 => std_logic_vector(to_unsigned(5,8) ,
23186	 => std_logic_vector(to_unsigned(9,8) ,
23187	 => std_logic_vector(to_unsigned(13,8) ,
23188	 => std_logic_vector(to_unsigned(18,8) ,
23189	 => std_logic_vector(to_unsigned(21,8) ,
23190	 => std_logic_vector(to_unsigned(19,8) ,
23191	 => std_logic_vector(to_unsigned(17,8) ,
23192	 => std_logic_vector(to_unsigned(45,8) ,
23193	 => std_logic_vector(to_unsigned(141,8) ,
23194	 => std_logic_vector(to_unsigned(164,8) ,
23195	 => std_logic_vector(to_unsigned(156,8) ,
23196	 => std_logic_vector(to_unsigned(156,8) ,
23197	 => std_logic_vector(to_unsigned(157,8) ,
23198	 => std_logic_vector(to_unsigned(154,8) ,
23199	 => std_logic_vector(to_unsigned(156,8) ,
23200	 => std_logic_vector(to_unsigned(138,8) ,
23201	 => std_logic_vector(to_unsigned(108,8) ,
23202	 => std_logic_vector(to_unsigned(104,8) ,
23203	 => std_logic_vector(to_unsigned(100,8) ,
23204	 => std_logic_vector(to_unsigned(97,8) ,
23205	 => std_logic_vector(to_unsigned(107,8) ,
23206	 => std_logic_vector(to_unsigned(95,8) ,
23207	 => std_logic_vector(to_unsigned(9,8) ,
23208	 => std_logic_vector(to_unsigned(2,8) ,
23209	 => std_logic_vector(to_unsigned(3,8) ,
23210	 => std_logic_vector(to_unsigned(3,8) ,
23211	 => std_logic_vector(to_unsigned(2,8) ,
23212	 => std_logic_vector(to_unsigned(3,8) ,
23213	 => std_logic_vector(to_unsigned(6,8) ,
23214	 => std_logic_vector(to_unsigned(9,8) ,
23215	 => std_logic_vector(to_unsigned(10,8) ,
23216	 => std_logic_vector(to_unsigned(17,8) ,
23217	 => std_logic_vector(to_unsigned(37,8) ,
23218	 => std_logic_vector(to_unsigned(44,8) ,
23219	 => std_logic_vector(to_unsigned(36,8) ,
23220	 => std_logic_vector(to_unsigned(24,8) ,
23221	 => std_logic_vector(to_unsigned(16,8) ,
23222	 => std_logic_vector(to_unsigned(22,8) ,
23223	 => std_logic_vector(to_unsigned(40,8) ,
23224	 => std_logic_vector(to_unsigned(63,8) ,
23225	 => std_logic_vector(to_unsigned(87,8) ,
23226	 => std_logic_vector(to_unsigned(130,8) ,
23227	 => std_logic_vector(to_unsigned(147,8) ,
23228	 => std_logic_vector(to_unsigned(125,8) ,
23229	 => std_logic_vector(to_unsigned(116,8) ,
23230	 => std_logic_vector(to_unsigned(111,8) ,
23231	 => std_logic_vector(to_unsigned(121,8) ,
23232	 => std_logic_vector(to_unsigned(116,8) ,
23233	 => std_logic_vector(to_unsigned(11,8) ,
23234	 => std_logic_vector(to_unsigned(0,8) ,
23235	 => std_logic_vector(to_unsigned(1,8) ,
23236	 => std_logic_vector(to_unsigned(1,8) ,
23237	 => std_logic_vector(to_unsigned(3,8) ,
23238	 => std_logic_vector(to_unsigned(3,8) ,
23239	 => std_logic_vector(to_unsigned(3,8) ,
23240	 => std_logic_vector(to_unsigned(2,8) ,
23241	 => std_logic_vector(to_unsigned(4,8) ,
23242	 => std_logic_vector(to_unsigned(36,8) ,
23243	 => std_logic_vector(to_unsigned(90,8) ,
23244	 => std_logic_vector(to_unsigned(71,8) ,
23245	 => std_logic_vector(to_unsigned(49,8) ,
23246	 => std_logic_vector(to_unsigned(104,8) ,
23247	 => std_logic_vector(to_unsigned(139,8) ,
23248	 => std_logic_vector(to_unsigned(131,8) ,
23249	 => std_logic_vector(to_unsigned(142,8) ,
23250	 => std_logic_vector(to_unsigned(138,8) ,
23251	 => std_logic_vector(to_unsigned(133,8) ,
23252	 => std_logic_vector(to_unsigned(133,8) ,
23253	 => std_logic_vector(to_unsigned(133,8) ,
23254	 => std_logic_vector(to_unsigned(134,8) ,
23255	 => std_logic_vector(to_unsigned(136,8) ,
23256	 => std_logic_vector(to_unsigned(138,8) ,
23257	 => std_logic_vector(to_unsigned(139,8) ,
23258	 => std_logic_vector(to_unsigned(138,8) ,
23259	 => std_logic_vector(to_unsigned(139,8) ,
23260	 => std_logic_vector(to_unsigned(138,8) ,
23261	 => std_logic_vector(to_unsigned(136,8) ,
23262	 => std_logic_vector(to_unsigned(136,8) ,
23263	 => std_logic_vector(to_unsigned(32,8) ,
23264	 => std_logic_vector(to_unsigned(4,8) ,
23265	 => std_logic_vector(to_unsigned(9,8) ,
23266	 => std_logic_vector(to_unsigned(11,8) ,
23267	 => std_logic_vector(to_unsigned(22,8) ,
23268	 => std_logic_vector(to_unsigned(22,8) ,
23269	 => std_logic_vector(to_unsigned(12,8) ,
23270	 => std_logic_vector(to_unsigned(13,8) ,
23271	 => std_logic_vector(to_unsigned(3,8) ,
23272	 => std_logic_vector(to_unsigned(1,8) ,
23273	 => std_logic_vector(to_unsigned(3,8) ,
23274	 => std_logic_vector(to_unsigned(4,8) ,
23275	 => std_logic_vector(to_unsigned(54,8) ,
23276	 => std_logic_vector(to_unsigned(151,8) ,
23277	 => std_logic_vector(to_unsigned(144,8) ,
23278	 => std_logic_vector(to_unsigned(144,8) ,
23279	 => std_logic_vector(to_unsigned(136,8) ,
23280	 => std_logic_vector(to_unsigned(147,8) ,
23281	 => std_logic_vector(to_unsigned(133,8) ,
23282	 => std_logic_vector(to_unsigned(122,8) ,
23283	 => std_logic_vector(to_unsigned(136,8) ,
23284	 => std_logic_vector(to_unsigned(142,8) ,
23285	 => std_logic_vector(to_unsigned(146,8) ,
23286	 => std_logic_vector(to_unsigned(139,8) ,
23287	 => std_logic_vector(to_unsigned(139,8) ,
23288	 => std_logic_vector(to_unsigned(151,8) ,
23289	 => std_logic_vector(to_unsigned(151,8) ,
23290	 => std_logic_vector(to_unsigned(157,8) ,
23291	 => std_logic_vector(to_unsigned(139,8) ,
23292	 => std_logic_vector(to_unsigned(118,8) ,
23293	 => std_logic_vector(to_unsigned(81,8) ,
23294	 => std_logic_vector(to_unsigned(7,8) ,
23295	 => std_logic_vector(to_unsigned(1,8) ,
23296	 => std_logic_vector(to_unsigned(7,8) ,
23297	 => std_logic_vector(to_unsigned(86,8) ,
23298	 => std_logic_vector(to_unsigned(166,8) ,
23299	 => std_logic_vector(to_unsigned(154,8) ,
23300	 => std_logic_vector(to_unsigned(159,8) ,
23301	 => std_logic_vector(to_unsigned(163,8) ,
23302	 => std_logic_vector(to_unsigned(159,8) ,
23303	 => std_logic_vector(to_unsigned(159,8) ,
23304	 => std_logic_vector(to_unsigned(159,8) ,
23305	 => std_logic_vector(to_unsigned(161,8) ,
23306	 => std_logic_vector(to_unsigned(161,8) ,
23307	 => std_logic_vector(to_unsigned(159,8) ,
23308	 => std_logic_vector(to_unsigned(159,8) ,
23309	 => std_logic_vector(to_unsigned(161,8) ,
23310	 => std_logic_vector(to_unsigned(154,8) ,
23311	 => std_logic_vector(to_unsigned(157,8) ,
23312	 => std_logic_vector(to_unsigned(147,8) ,
23313	 => std_logic_vector(to_unsigned(149,8) ,
23314	 => std_logic_vector(to_unsigned(141,8) ,
23315	 => std_logic_vector(to_unsigned(138,8) ,
23316	 => std_logic_vector(to_unsigned(64,8) ,
23317	 => std_logic_vector(to_unsigned(5,8) ,
23318	 => std_logic_vector(to_unsigned(3,8) ,
23319	 => std_logic_vector(to_unsigned(15,8) ,
23320	 => std_logic_vector(to_unsigned(25,8) ,
23321	 => std_logic_vector(to_unsigned(8,8) ,
23322	 => std_logic_vector(to_unsigned(7,8) ,
23323	 => std_logic_vector(to_unsigned(13,8) ,
23324	 => std_logic_vector(to_unsigned(13,8) ,
23325	 => std_logic_vector(to_unsigned(9,8) ,
23326	 => std_logic_vector(to_unsigned(36,8) ,
23327	 => std_logic_vector(to_unsigned(108,8) ,
23328	 => std_logic_vector(to_unsigned(97,8) ,
23329	 => std_logic_vector(to_unsigned(103,8) ,
23330	 => std_logic_vector(to_unsigned(105,8) ,
23331	 => std_logic_vector(to_unsigned(97,8) ,
23332	 => std_logic_vector(to_unsigned(109,8) ,
23333	 => std_logic_vector(to_unsigned(116,8) ,
23334	 => std_logic_vector(to_unsigned(119,8) ,
23335	 => std_logic_vector(to_unsigned(101,8) ,
23336	 => std_logic_vector(to_unsigned(87,8) ,
23337	 => std_logic_vector(to_unsigned(92,8) ,
23338	 => std_logic_vector(to_unsigned(86,8) ,
23339	 => std_logic_vector(to_unsigned(85,8) ,
23340	 => std_logic_vector(to_unsigned(80,8) ,
23341	 => std_logic_vector(to_unsigned(119,8) ,
23342	 => std_logic_vector(to_unsigned(144,8) ,
23343	 => std_logic_vector(to_unsigned(96,8) ,
23344	 => std_logic_vector(to_unsigned(93,8) ,
23345	 => std_logic_vector(to_unsigned(111,8) ,
23346	 => std_logic_vector(to_unsigned(114,8) ,
23347	 => std_logic_vector(to_unsigned(103,8) ,
23348	 => std_logic_vector(to_unsigned(104,8) ,
23349	 => std_logic_vector(to_unsigned(136,8) ,
23350	 => std_logic_vector(to_unsigned(163,8) ,
23351	 => std_logic_vector(to_unsigned(157,8) ,
23352	 => std_logic_vector(to_unsigned(163,8) ,
23353	 => std_logic_vector(to_unsigned(133,8) ,
23354	 => std_logic_vector(to_unsigned(121,8) ,
23355	 => std_logic_vector(to_unsigned(127,8) ,
23356	 => std_logic_vector(to_unsigned(134,8) ,
23357	 => std_logic_vector(to_unsigned(131,8) ,
23358	 => std_logic_vector(to_unsigned(116,8) ,
23359	 => std_logic_vector(to_unsigned(108,8) ,
23360	 => std_logic_vector(to_unsigned(104,8) ,
23361	 => std_logic_vector(to_unsigned(159,8) ,
23362	 => std_logic_vector(to_unsigned(161,8) ,
23363	 => std_logic_vector(to_unsigned(157,8) ,
23364	 => std_logic_vector(to_unsigned(156,8) ,
23365	 => std_logic_vector(to_unsigned(159,8) ,
23366	 => std_logic_vector(to_unsigned(168,8) ,
23367	 => std_logic_vector(to_unsigned(130,8) ,
23368	 => std_logic_vector(to_unsigned(44,8) ,
23369	 => std_logic_vector(to_unsigned(53,8) ,
23370	 => std_logic_vector(to_unsigned(51,8) ,
23371	 => std_logic_vector(to_unsigned(15,8) ,
23372	 => std_logic_vector(to_unsigned(17,8) ,
23373	 => std_logic_vector(to_unsigned(20,8) ,
23374	 => std_logic_vector(to_unsigned(7,8) ,
23375	 => std_logic_vector(to_unsigned(6,8) ,
23376	 => std_logic_vector(to_unsigned(10,8) ,
23377	 => std_logic_vector(to_unsigned(8,8) ,
23378	 => std_logic_vector(to_unsigned(62,8) ,
23379	 => std_logic_vector(to_unsigned(76,8) ,
23380	 => std_logic_vector(to_unsigned(14,8) ,
23381	 => std_logic_vector(to_unsigned(32,8) ,
23382	 => std_logic_vector(to_unsigned(4,8) ,
23383	 => std_logic_vector(to_unsigned(0,8) ,
23384	 => std_logic_vector(to_unsigned(3,8) ,
23385	 => std_logic_vector(to_unsigned(2,8) ,
23386	 => std_logic_vector(to_unsigned(2,8) ,
23387	 => std_logic_vector(to_unsigned(4,8) ,
23388	 => std_logic_vector(to_unsigned(4,8) ,
23389	 => std_logic_vector(to_unsigned(2,8) ,
23390	 => std_logic_vector(to_unsigned(3,8) ,
23391	 => std_logic_vector(to_unsigned(7,8) ,
23392	 => std_logic_vector(to_unsigned(2,8) ,
23393	 => std_logic_vector(to_unsigned(2,8) ,
23394	 => std_logic_vector(to_unsigned(10,8) ,
23395	 => std_logic_vector(to_unsigned(9,8) ,
23396	 => std_logic_vector(to_unsigned(49,8) ,
23397	 => std_logic_vector(to_unsigned(27,8) ,
23398	 => std_logic_vector(to_unsigned(2,8) ,
23399	 => std_logic_vector(to_unsigned(2,8) ,
23400	 => std_logic_vector(to_unsigned(7,8) ,
23401	 => std_logic_vector(to_unsigned(18,8) ,
23402	 => std_logic_vector(to_unsigned(14,8) ,
23403	 => std_logic_vector(to_unsigned(17,8) ,
23404	 => std_logic_vector(to_unsigned(20,8) ,
23405	 => std_logic_vector(to_unsigned(24,8) ,
23406	 => std_logic_vector(to_unsigned(36,8) ,
23407	 => std_logic_vector(to_unsigned(37,8) ,
23408	 => std_logic_vector(to_unsigned(37,8) ,
23409	 => std_logic_vector(to_unsigned(29,8) ,
23410	 => std_logic_vector(to_unsigned(10,8) ,
23411	 => std_logic_vector(to_unsigned(68,8) ,
23412	 => std_logic_vector(to_unsigned(190,8) ,
23413	 => std_logic_vector(to_unsigned(161,8) ,
23414	 => std_logic_vector(to_unsigned(157,8) ,
23415	 => std_logic_vector(to_unsigned(170,8) ,
23416	 => std_logic_vector(to_unsigned(91,8) ,
23417	 => std_logic_vector(to_unsigned(6,8) ,
23418	 => std_logic_vector(to_unsigned(2,8) ,
23419	 => std_logic_vector(to_unsigned(3,8) ,
23420	 => std_logic_vector(to_unsigned(2,8) ,
23421	 => std_logic_vector(to_unsigned(3,8) ,
23422	 => std_logic_vector(to_unsigned(3,8) ,
23423	 => std_logic_vector(to_unsigned(5,8) ,
23424	 => std_logic_vector(to_unsigned(6,8) ,
23425	 => std_logic_vector(to_unsigned(8,8) ,
23426	 => std_logic_vector(to_unsigned(6,8) ,
23427	 => std_logic_vector(to_unsigned(4,8) ,
23428	 => std_logic_vector(to_unsigned(11,8) ,
23429	 => std_logic_vector(to_unsigned(6,8) ,
23430	 => std_logic_vector(to_unsigned(6,8) ,
23431	 => std_logic_vector(to_unsigned(4,8) ,
23432	 => std_logic_vector(to_unsigned(8,8) ,
23433	 => std_logic_vector(to_unsigned(85,8) ,
23434	 => std_logic_vector(to_unsigned(74,8) ,
23435	 => std_logic_vector(to_unsigned(5,8) ,
23436	 => std_logic_vector(to_unsigned(15,8) ,
23437	 => std_logic_vector(to_unsigned(104,8) ,
23438	 => std_logic_vector(to_unsigned(152,8) ,
23439	 => std_logic_vector(to_unsigned(130,8) ,
23440	 => std_logic_vector(to_unsigned(36,8) ,
23441	 => std_logic_vector(to_unsigned(8,8) ,
23442	 => std_logic_vector(to_unsigned(17,8) ,
23443	 => std_logic_vector(to_unsigned(22,8) ,
23444	 => std_logic_vector(to_unsigned(27,8) ,
23445	 => std_logic_vector(to_unsigned(45,8) ,
23446	 => std_logic_vector(to_unsigned(87,8) ,
23447	 => std_logic_vector(to_unsigned(163,8) ,
23448	 => std_logic_vector(to_unsigned(170,8) ,
23449	 => std_logic_vector(to_unsigned(139,8) ,
23450	 => std_logic_vector(to_unsigned(115,8) ,
23451	 => std_logic_vector(to_unsigned(141,8) ,
23452	 => std_logic_vector(to_unsigned(166,8) ,
23453	 => std_logic_vector(to_unsigned(161,8) ,
23454	 => std_logic_vector(to_unsigned(175,8) ,
23455	 => std_logic_vector(to_unsigned(124,8) ,
23456	 => std_logic_vector(to_unsigned(115,8) ,
23457	 => std_logic_vector(to_unsigned(164,8) ,
23458	 => std_logic_vector(to_unsigned(166,8) ,
23459	 => std_logic_vector(to_unsigned(168,8) ,
23460	 => std_logic_vector(to_unsigned(166,8) ,
23461	 => std_logic_vector(to_unsigned(163,8) ,
23462	 => std_logic_vector(to_unsigned(163,8) ,
23463	 => std_logic_vector(to_unsigned(128,8) ,
23464	 => std_logic_vector(to_unsigned(111,8) ,
23465	 => std_logic_vector(to_unsigned(127,8) ,
23466	 => std_logic_vector(to_unsigned(136,8) ,
23467	 => std_logic_vector(to_unsigned(115,8) ,
23468	 => std_logic_vector(to_unsigned(151,8) ,
23469	 => std_logic_vector(to_unsigned(157,8) ,
23470	 => std_logic_vector(to_unsigned(161,8) ,
23471	 => std_logic_vector(to_unsigned(163,8) ,
23472	 => std_logic_vector(to_unsigned(159,8) ,
23473	 => std_logic_vector(to_unsigned(156,8) ,
23474	 => std_logic_vector(to_unsigned(152,8) ,
23475	 => std_logic_vector(to_unsigned(198,8) ,
23476	 => std_logic_vector(to_unsigned(78,8) ,
23477	 => std_logic_vector(to_unsigned(2,8) ,
23478	 => std_logic_vector(to_unsigned(0,8) ,
23479	 => std_logic_vector(to_unsigned(1,8) ,
23480	 => std_logic_vector(to_unsigned(4,8) ,
23481	 => std_logic_vector(to_unsigned(5,8) ,
23482	 => std_logic_vector(to_unsigned(5,8) ,
23483	 => std_logic_vector(to_unsigned(8,8) ,
23484	 => std_logic_vector(to_unsigned(11,8) ,
23485	 => std_logic_vector(to_unsigned(9,8) ,
23486	 => std_logic_vector(to_unsigned(5,8) ,
23487	 => std_logic_vector(to_unsigned(39,8) ,
23488	 => std_logic_vector(to_unsigned(109,8) ,
23489	 => std_logic_vector(to_unsigned(134,8) ,
23490	 => std_logic_vector(to_unsigned(161,8) ,
23491	 => std_logic_vector(to_unsigned(144,8) ,
23492	 => std_logic_vector(to_unsigned(144,8) ,
23493	 => std_logic_vector(to_unsigned(152,8) ,
23494	 => std_logic_vector(to_unsigned(152,8) ,
23495	 => std_logic_vector(to_unsigned(156,8) ,
23496	 => std_logic_vector(to_unsigned(154,8) ,
23497	 => std_logic_vector(to_unsigned(152,8) ,
23498	 => std_logic_vector(to_unsigned(154,8) ,
23499	 => std_logic_vector(to_unsigned(156,8) ,
23500	 => std_logic_vector(to_unsigned(151,8) ,
23501	 => std_logic_vector(to_unsigned(146,8) ,
23502	 => std_logic_vector(to_unsigned(157,8) ,
23503	 => std_logic_vector(to_unsigned(141,8) ,
23504	 => std_logic_vector(to_unsigned(14,8) ,
23505	 => std_logic_vector(to_unsigned(2,8) ,
23506	 => std_logic_vector(to_unsigned(20,8) ,
23507	 => std_logic_vector(to_unsigned(29,8) ,
23508	 => std_logic_vector(to_unsigned(15,8) ,
23509	 => std_logic_vector(to_unsigned(12,8) ,
23510	 => std_logic_vector(to_unsigned(14,8) ,
23511	 => std_logic_vector(to_unsigned(15,8) ,
23512	 => std_logic_vector(to_unsigned(30,8) ,
23513	 => std_logic_vector(to_unsigned(86,8) ,
23514	 => std_logic_vector(to_unsigned(133,8) ,
23515	 => std_logic_vector(to_unsigned(151,8) ,
23516	 => std_logic_vector(to_unsigned(161,8) ,
23517	 => std_logic_vector(to_unsigned(159,8) ,
23518	 => std_logic_vector(to_unsigned(156,8) ,
23519	 => std_logic_vector(to_unsigned(161,8) ,
23520	 => std_logic_vector(to_unsigned(144,8) ,
23521	 => std_logic_vector(to_unsigned(107,8) ,
23522	 => std_logic_vector(to_unsigned(99,8) ,
23523	 => std_logic_vector(to_unsigned(99,8) ,
23524	 => std_logic_vector(to_unsigned(109,8) ,
23525	 => std_logic_vector(to_unsigned(84,8) ,
23526	 => std_logic_vector(to_unsigned(29,8) ,
23527	 => std_logic_vector(to_unsigned(3,8) ,
23528	 => std_logic_vector(to_unsigned(2,8) ,
23529	 => std_logic_vector(to_unsigned(3,8) ,
23530	 => std_logic_vector(to_unsigned(2,8) ,
23531	 => std_logic_vector(to_unsigned(4,8) ,
23532	 => std_logic_vector(to_unsigned(7,8) ,
23533	 => std_logic_vector(to_unsigned(10,8) ,
23534	 => std_logic_vector(to_unsigned(11,8) ,
23535	 => std_logic_vector(to_unsigned(8,8) ,
23536	 => std_logic_vector(to_unsigned(15,8) ,
23537	 => std_logic_vector(to_unsigned(37,8) ,
23538	 => std_logic_vector(to_unsigned(43,8) ,
23539	 => std_logic_vector(to_unsigned(46,8) ,
23540	 => std_logic_vector(to_unsigned(43,8) ,
23541	 => std_logic_vector(to_unsigned(22,8) ,
23542	 => std_logic_vector(to_unsigned(28,8) ,
23543	 => std_logic_vector(to_unsigned(52,8) ,
23544	 => std_logic_vector(to_unsigned(61,8) ,
23545	 => std_logic_vector(to_unsigned(61,8) ,
23546	 => std_logic_vector(to_unsigned(78,8) ,
23547	 => std_logic_vector(to_unsigned(139,8) ,
23548	 => std_logic_vector(to_unsigned(136,8) ,
23549	 => std_logic_vector(to_unsigned(114,8) ,
23550	 => std_logic_vector(to_unsigned(111,8) ,
23551	 => std_logic_vector(to_unsigned(133,8) ,
23552	 => std_logic_vector(to_unsigned(127,8) ,
23553	 => std_logic_vector(to_unsigned(17,8) ,
23554	 => std_logic_vector(to_unsigned(0,8) ,
23555	 => std_logic_vector(to_unsigned(0,8) ,
23556	 => std_logic_vector(to_unsigned(0,8) ,
23557	 => std_logic_vector(to_unsigned(2,8) ,
23558	 => std_logic_vector(to_unsigned(1,8) ,
23559	 => std_logic_vector(to_unsigned(1,8) ,
23560	 => std_logic_vector(to_unsigned(3,8) ,
23561	 => std_logic_vector(to_unsigned(27,8) ,
23562	 => std_logic_vector(to_unsigned(59,8) ,
23563	 => std_logic_vector(to_unsigned(41,8) ,
23564	 => std_logic_vector(to_unsigned(44,8) ,
23565	 => std_logic_vector(to_unsigned(72,8) ,
23566	 => std_logic_vector(to_unsigned(131,8) ,
23567	 => std_logic_vector(to_unsigned(136,8) ,
23568	 => std_logic_vector(to_unsigned(136,8) ,
23569	 => std_logic_vector(to_unsigned(141,8) ,
23570	 => std_logic_vector(to_unsigned(133,8) ,
23571	 => std_logic_vector(to_unsigned(139,8) ,
23572	 => std_logic_vector(to_unsigned(139,8) ,
23573	 => std_logic_vector(to_unsigned(133,8) ,
23574	 => std_logic_vector(to_unsigned(133,8) ,
23575	 => std_logic_vector(to_unsigned(139,8) ,
23576	 => std_logic_vector(to_unsigned(139,8) ,
23577	 => std_logic_vector(to_unsigned(138,8) ,
23578	 => std_logic_vector(to_unsigned(136,8) ,
23579	 => std_logic_vector(to_unsigned(134,8) ,
23580	 => std_logic_vector(to_unsigned(139,8) ,
23581	 => std_logic_vector(to_unsigned(131,8) ,
23582	 => std_logic_vector(to_unsigned(146,8) ,
23583	 => std_logic_vector(to_unsigned(101,8) ,
23584	 => std_logic_vector(to_unsigned(7,8) ,
23585	 => std_logic_vector(to_unsigned(1,8) ,
23586	 => std_logic_vector(to_unsigned(2,8) ,
23587	 => std_logic_vector(to_unsigned(7,8) ,
23588	 => std_logic_vector(to_unsigned(18,8) ,
23589	 => std_logic_vector(to_unsigned(29,8) ,
23590	 => std_logic_vector(to_unsigned(23,8) ,
23591	 => std_logic_vector(to_unsigned(8,8) ,
23592	 => std_logic_vector(to_unsigned(5,8) ,
23593	 => std_logic_vector(to_unsigned(2,8) ,
23594	 => std_logic_vector(to_unsigned(5,8) ,
23595	 => std_logic_vector(to_unsigned(122,8) ,
23596	 => std_logic_vector(to_unsigned(161,8) ,
23597	 => std_logic_vector(to_unsigned(131,8) ,
23598	 => std_logic_vector(to_unsigned(142,8) ,
23599	 => std_logic_vector(to_unsigned(142,8) ,
23600	 => std_logic_vector(to_unsigned(141,8) ,
23601	 => std_logic_vector(to_unsigned(131,8) ,
23602	 => std_logic_vector(to_unsigned(119,8) ,
23603	 => std_logic_vector(to_unsigned(131,8) ,
23604	 => std_logic_vector(to_unsigned(149,8) ,
23605	 => std_logic_vector(to_unsigned(163,8) ,
23606	 => std_logic_vector(to_unsigned(157,8) ,
23607	 => std_logic_vector(to_unsigned(144,8) ,
23608	 => std_logic_vector(to_unsigned(147,8) ,
23609	 => std_logic_vector(to_unsigned(130,8) ,
23610	 => std_logic_vector(to_unsigned(111,8) ,
23611	 => std_logic_vector(to_unsigned(78,8) ,
23612	 => std_logic_vector(to_unsigned(50,8) ,
23613	 => std_logic_vector(to_unsigned(26,8) ,
23614	 => std_logic_vector(to_unsigned(9,8) ,
23615	 => std_logic_vector(to_unsigned(4,8) ,
23616	 => std_logic_vector(to_unsigned(4,8) ,
23617	 => std_logic_vector(to_unsigned(26,8) ,
23618	 => std_logic_vector(to_unsigned(62,8) ,
23619	 => std_logic_vector(to_unsigned(131,8) ,
23620	 => std_logic_vector(to_unsigned(171,8) ,
23621	 => std_logic_vector(to_unsigned(163,8) ,
23622	 => std_logic_vector(to_unsigned(166,8) ,
23623	 => std_logic_vector(to_unsigned(159,8) ,
23624	 => std_logic_vector(to_unsigned(161,8) ,
23625	 => std_logic_vector(to_unsigned(163,8) ,
23626	 => std_logic_vector(to_unsigned(163,8) ,
23627	 => std_logic_vector(to_unsigned(164,8) ,
23628	 => std_logic_vector(to_unsigned(159,8) ,
23629	 => std_logic_vector(to_unsigned(161,8) ,
23630	 => std_logic_vector(to_unsigned(159,8) ,
23631	 => std_logic_vector(to_unsigned(159,8) ,
23632	 => std_logic_vector(to_unsigned(159,8) ,
23633	 => std_logic_vector(to_unsigned(156,8) ,
23634	 => std_logic_vector(to_unsigned(151,8) ,
23635	 => std_logic_vector(to_unsigned(139,8) ,
23636	 => std_logic_vector(to_unsigned(118,8) ,
23637	 => std_logic_vector(to_unsigned(13,8) ,
23638	 => std_logic_vector(to_unsigned(1,8) ,
23639	 => std_logic_vector(to_unsigned(4,8) ,
23640	 => std_logic_vector(to_unsigned(1,8) ,
23641	 => std_logic_vector(to_unsigned(8,8) ,
23642	 => std_logic_vector(to_unsigned(18,8) ,
23643	 => std_logic_vector(to_unsigned(10,8) ,
23644	 => std_logic_vector(to_unsigned(14,8) ,
23645	 => std_logic_vector(to_unsigned(14,8) ,
23646	 => std_logic_vector(to_unsigned(29,8) ,
23647	 => std_logic_vector(to_unsigned(100,8) ,
23648	 => std_logic_vector(to_unsigned(115,8) ,
23649	 => std_logic_vector(to_unsigned(104,8) ,
23650	 => std_logic_vector(to_unsigned(114,8) ,
23651	 => std_logic_vector(to_unsigned(115,8) ,
23652	 => std_logic_vector(to_unsigned(104,8) ,
23653	 => std_logic_vector(to_unsigned(104,8) ,
23654	 => std_logic_vector(to_unsigned(97,8) ,
23655	 => std_logic_vector(to_unsigned(88,8) ,
23656	 => std_logic_vector(to_unsigned(91,8) ,
23657	 => std_logic_vector(to_unsigned(95,8) ,
23658	 => std_logic_vector(to_unsigned(93,8) ,
23659	 => std_logic_vector(to_unsigned(92,8) ,
23660	 => std_logic_vector(to_unsigned(87,8) ,
23661	 => std_logic_vector(to_unsigned(97,8) ,
23662	 => std_logic_vector(to_unsigned(119,8) ,
23663	 => std_logic_vector(to_unsigned(101,8) ,
23664	 => std_logic_vector(to_unsigned(84,8) ,
23665	 => std_logic_vector(to_unsigned(95,8) ,
23666	 => std_logic_vector(to_unsigned(105,8) ,
23667	 => std_logic_vector(to_unsigned(109,8) ,
23668	 => std_logic_vector(to_unsigned(95,8) ,
23669	 => std_logic_vector(to_unsigned(111,8) ,
23670	 => std_logic_vector(to_unsigned(159,8) ,
23671	 => std_logic_vector(to_unsigned(164,8) ,
23672	 => std_logic_vector(to_unsigned(159,8) ,
23673	 => std_logic_vector(to_unsigned(142,8) ,
23674	 => std_logic_vector(to_unsigned(130,8) ,
23675	 => std_logic_vector(to_unsigned(125,8) ,
23676	 => std_logic_vector(to_unsigned(121,8) ,
23677	 => std_logic_vector(to_unsigned(130,8) ,
23678	 => std_logic_vector(to_unsigned(122,8) ,
23679	 => std_logic_vector(to_unsigned(103,8) ,
23680	 => std_logic_vector(to_unsigned(99,8) ,
23681	 => std_logic_vector(to_unsigned(163,8) ,
23682	 => std_logic_vector(to_unsigned(164,8) ,
23683	 => std_logic_vector(to_unsigned(163,8) ,
23684	 => std_logic_vector(to_unsigned(159,8) ,
23685	 => std_logic_vector(to_unsigned(159,8) ,
23686	 => std_logic_vector(to_unsigned(168,8) ,
23687	 => std_logic_vector(to_unsigned(138,8) ,
23688	 => std_logic_vector(to_unsigned(49,8) ,
23689	 => std_logic_vector(to_unsigned(25,8) ,
23690	 => std_logic_vector(to_unsigned(53,8) ,
23691	 => std_logic_vector(to_unsigned(35,8) ,
23692	 => std_logic_vector(to_unsigned(4,8) ,
23693	 => std_logic_vector(to_unsigned(9,8) ,
23694	 => std_logic_vector(to_unsigned(11,8) ,
23695	 => std_logic_vector(to_unsigned(8,8) ,
23696	 => std_logic_vector(to_unsigned(11,8) ,
23697	 => std_logic_vector(to_unsigned(43,8) ,
23698	 => std_logic_vector(to_unsigned(79,8) ,
23699	 => std_logic_vector(to_unsigned(103,8) ,
23700	 => std_logic_vector(to_unsigned(21,8) ,
23701	 => std_logic_vector(to_unsigned(20,8) ,
23702	 => std_logic_vector(to_unsigned(11,8) ,
23703	 => std_logic_vector(to_unsigned(0,8) ,
23704	 => std_logic_vector(to_unsigned(1,8) ,
23705	 => std_logic_vector(to_unsigned(2,8) ,
23706	 => std_logic_vector(to_unsigned(5,8) ,
23707	 => std_logic_vector(to_unsigned(4,8) ,
23708	 => std_logic_vector(to_unsigned(4,8) ,
23709	 => std_logic_vector(to_unsigned(1,8) ,
23710	 => std_logic_vector(to_unsigned(3,8) ,
23711	 => std_logic_vector(to_unsigned(10,8) ,
23712	 => std_logic_vector(to_unsigned(4,8) ,
23713	 => std_logic_vector(to_unsigned(2,8) ,
23714	 => std_logic_vector(to_unsigned(8,8) ,
23715	 => std_logic_vector(to_unsigned(10,8) ,
23716	 => std_logic_vector(to_unsigned(27,8) ,
23717	 => std_logic_vector(to_unsigned(27,8) ,
23718	 => std_logic_vector(to_unsigned(3,8) ,
23719	 => std_logic_vector(to_unsigned(2,8) ,
23720	 => std_logic_vector(to_unsigned(7,8) ,
23721	 => std_logic_vector(to_unsigned(12,8) ,
23722	 => std_logic_vector(to_unsigned(9,8) ,
23723	 => std_logic_vector(to_unsigned(9,8) ,
23724	 => std_logic_vector(to_unsigned(16,8) ,
23725	 => std_logic_vector(to_unsigned(34,8) ,
23726	 => std_logic_vector(to_unsigned(41,8) ,
23727	 => std_logic_vector(to_unsigned(43,8) ,
23728	 => std_logic_vector(to_unsigned(42,8) ,
23729	 => std_logic_vector(to_unsigned(30,8) ,
23730	 => std_logic_vector(to_unsigned(43,8) ,
23731	 => std_logic_vector(to_unsigned(154,8) ,
23732	 => std_logic_vector(to_unsigned(177,8) ,
23733	 => std_logic_vector(to_unsigned(161,8) ,
23734	 => std_logic_vector(to_unsigned(156,8) ,
23735	 => std_logic_vector(to_unsigned(181,8) ,
23736	 => std_logic_vector(to_unsigned(104,8) ,
23737	 => std_logic_vector(to_unsigned(6,8) ,
23738	 => std_logic_vector(to_unsigned(4,8) ,
23739	 => std_logic_vector(to_unsigned(6,8) ,
23740	 => std_logic_vector(to_unsigned(7,8) ,
23741	 => std_logic_vector(to_unsigned(6,8) ,
23742	 => std_logic_vector(to_unsigned(3,8) ,
23743	 => std_logic_vector(to_unsigned(4,8) ,
23744	 => std_logic_vector(to_unsigned(5,8) ,
23745	 => std_logic_vector(to_unsigned(6,8) ,
23746	 => std_logic_vector(to_unsigned(3,8) ,
23747	 => std_logic_vector(to_unsigned(2,8) ,
23748	 => std_logic_vector(to_unsigned(6,8) ,
23749	 => std_logic_vector(to_unsigned(6,8) ,
23750	 => std_logic_vector(to_unsigned(6,8) ,
23751	 => std_logic_vector(to_unsigned(8,8) ,
23752	 => std_logic_vector(to_unsigned(3,8) ,
23753	 => std_logic_vector(to_unsigned(17,8) ,
23754	 => std_logic_vector(to_unsigned(90,8) ,
23755	 => std_logic_vector(to_unsigned(41,8) ,
23756	 => std_logic_vector(to_unsigned(1,8) ,
23757	 => std_logic_vector(to_unsigned(58,8) ,
23758	 => std_logic_vector(to_unsigned(130,8) ,
23759	 => std_logic_vector(to_unsigned(32,8) ,
23760	 => std_logic_vector(to_unsigned(4,8) ,
23761	 => std_logic_vector(to_unsigned(11,8) ,
23762	 => std_logic_vector(to_unsigned(15,8) ,
23763	 => std_logic_vector(to_unsigned(27,8) ,
23764	 => std_logic_vector(to_unsigned(35,8) ,
23765	 => std_logic_vector(to_unsigned(38,8) ,
23766	 => std_logic_vector(to_unsigned(48,8) ,
23767	 => std_logic_vector(to_unsigned(119,8) ,
23768	 => std_logic_vector(to_unsigned(166,8) ,
23769	 => std_logic_vector(to_unsigned(146,8) ,
23770	 => std_logic_vector(to_unsigned(116,8) ,
23771	 => std_logic_vector(to_unsigned(128,8) ,
23772	 => std_logic_vector(to_unsigned(166,8) ,
23773	 => std_logic_vector(to_unsigned(164,8) ,
23774	 => std_logic_vector(to_unsigned(166,8) ,
23775	 => std_logic_vector(to_unsigned(163,8) ,
23776	 => std_logic_vector(to_unsigned(161,8) ,
23777	 => std_logic_vector(to_unsigned(161,8) ,
23778	 => std_logic_vector(to_unsigned(166,8) ,
23779	 => std_logic_vector(to_unsigned(166,8) ,
23780	 => std_logic_vector(to_unsigned(161,8) ,
23781	 => std_logic_vector(to_unsigned(164,8) ,
23782	 => std_logic_vector(to_unsigned(159,8) ,
23783	 => std_logic_vector(to_unsigned(128,8) ,
23784	 => std_logic_vector(to_unsigned(125,8) ,
23785	 => std_logic_vector(to_unsigned(138,8) ,
23786	 => std_logic_vector(to_unsigned(127,8) ,
23787	 => std_logic_vector(to_unsigned(139,8) ,
23788	 => std_logic_vector(to_unsigned(157,8) ,
23789	 => std_logic_vector(to_unsigned(149,8) ,
23790	 => std_logic_vector(to_unsigned(159,8) ,
23791	 => std_logic_vector(to_unsigned(161,8) ,
23792	 => std_logic_vector(to_unsigned(156,8) ,
23793	 => std_logic_vector(to_unsigned(161,8) ,
23794	 => std_logic_vector(to_unsigned(166,8) ,
23795	 => std_logic_vector(to_unsigned(76,8) ,
23796	 => std_logic_vector(to_unsigned(12,8) ,
23797	 => std_logic_vector(to_unsigned(5,8) ,
23798	 => std_logic_vector(to_unsigned(4,8) ,
23799	 => std_logic_vector(to_unsigned(3,8) ,
23800	 => std_logic_vector(to_unsigned(4,8) ,
23801	 => std_logic_vector(to_unsigned(5,8) ,
23802	 => std_logic_vector(to_unsigned(7,8) ,
23803	 => std_logic_vector(to_unsigned(4,8) ,
23804	 => std_logic_vector(to_unsigned(4,8) ,
23805	 => std_logic_vector(to_unsigned(4,8) ,
23806	 => std_logic_vector(to_unsigned(6,8) ,
23807	 => std_logic_vector(to_unsigned(30,8) ,
23808	 => std_logic_vector(to_unsigned(37,8) ,
23809	 => std_logic_vector(to_unsigned(40,8) ,
23810	 => std_logic_vector(to_unsigned(84,8) ,
23811	 => std_logic_vector(to_unsigned(144,8) ,
23812	 => std_logic_vector(to_unsigned(159,8) ,
23813	 => std_logic_vector(to_unsigned(156,8) ,
23814	 => std_logic_vector(to_unsigned(156,8) ,
23815	 => std_logic_vector(to_unsigned(159,8) ,
23816	 => std_logic_vector(to_unsigned(159,8) ,
23817	 => std_logic_vector(to_unsigned(159,8) ,
23818	 => std_logic_vector(to_unsigned(156,8) ,
23819	 => std_logic_vector(to_unsigned(152,8) ,
23820	 => std_logic_vector(to_unsigned(152,8) ,
23821	 => std_logic_vector(to_unsigned(144,8) ,
23822	 => std_logic_vector(to_unsigned(166,8) ,
23823	 => std_logic_vector(to_unsigned(147,8) ,
23824	 => std_logic_vector(to_unsigned(15,8) ,
23825	 => std_logic_vector(to_unsigned(1,8) ,
23826	 => std_logic_vector(to_unsigned(14,8) ,
23827	 => std_logic_vector(to_unsigned(20,8) ,
23828	 => std_logic_vector(to_unsigned(10,8) ,
23829	 => std_logic_vector(to_unsigned(6,8) ,
23830	 => std_logic_vector(to_unsigned(8,8) ,
23831	 => std_logic_vector(to_unsigned(9,8) ,
23832	 => std_logic_vector(to_unsigned(22,8) ,
23833	 => std_logic_vector(to_unsigned(39,8) ,
23834	 => std_logic_vector(to_unsigned(55,8) ,
23835	 => std_logic_vector(to_unsigned(93,8) ,
23836	 => std_logic_vector(to_unsigned(136,8) ,
23837	 => std_logic_vector(to_unsigned(154,8) ,
23838	 => std_logic_vector(to_unsigned(151,8) ,
23839	 => std_logic_vector(to_unsigned(157,8) ,
23840	 => std_logic_vector(to_unsigned(144,8) ,
23841	 => std_logic_vector(to_unsigned(119,8) ,
23842	 => std_logic_vector(to_unsigned(109,8) ,
23843	 => std_logic_vector(to_unsigned(108,8) ,
23844	 => std_logic_vector(to_unsigned(86,8) ,
23845	 => std_logic_vector(to_unsigned(21,8) ,
23846	 => std_logic_vector(to_unsigned(5,8) ,
23847	 => std_logic_vector(to_unsigned(8,8) ,
23848	 => std_logic_vector(to_unsigned(7,8) ,
23849	 => std_logic_vector(to_unsigned(5,8) ,
23850	 => std_logic_vector(to_unsigned(3,8) ,
23851	 => std_logic_vector(to_unsigned(2,8) ,
23852	 => std_logic_vector(to_unsigned(6,8) ,
23853	 => std_logic_vector(to_unsigned(11,8) ,
23854	 => std_logic_vector(to_unsigned(11,8) ,
23855	 => std_logic_vector(to_unsigned(11,8) ,
23856	 => std_logic_vector(to_unsigned(16,8) ,
23857	 => std_logic_vector(to_unsigned(30,8) ,
23858	 => std_logic_vector(to_unsigned(32,8) ,
23859	 => std_logic_vector(to_unsigned(39,8) ,
23860	 => std_logic_vector(to_unsigned(37,8) ,
23861	 => std_logic_vector(to_unsigned(17,8) ,
23862	 => std_logic_vector(to_unsigned(23,8) ,
23863	 => std_logic_vector(to_unsigned(41,8) ,
23864	 => std_logic_vector(to_unsigned(63,8) ,
23865	 => std_logic_vector(to_unsigned(48,8) ,
23866	 => std_logic_vector(to_unsigned(41,8) ,
23867	 => std_logic_vector(to_unsigned(99,8) ,
23868	 => std_logic_vector(to_unsigned(122,8) ,
23869	 => std_logic_vector(to_unsigned(114,8) ,
23870	 => std_logic_vector(to_unsigned(112,8) ,
23871	 => std_logic_vector(to_unsigned(111,8) ,
23872	 => std_logic_vector(to_unsigned(121,8) ,
23873	 => std_logic_vector(to_unsigned(67,8) ,
23874	 => std_logic_vector(to_unsigned(4,8) ,
23875	 => std_logic_vector(to_unsigned(1,8) ,
23876	 => std_logic_vector(to_unsigned(1,8) ,
23877	 => std_logic_vector(to_unsigned(2,8) ,
23878	 => std_logic_vector(to_unsigned(2,8) ,
23879	 => std_logic_vector(to_unsigned(3,8) ,
23880	 => std_logic_vector(to_unsigned(19,8) ,
23881	 => std_logic_vector(to_unsigned(51,8) ,
23882	 => std_logic_vector(to_unsigned(46,8) ,
23883	 => std_logic_vector(to_unsigned(41,8) ,
23884	 => std_logic_vector(to_unsigned(34,8) ,
23885	 => std_logic_vector(to_unsigned(57,8) ,
23886	 => std_logic_vector(to_unsigned(133,8) ,
23887	 => std_logic_vector(to_unsigned(141,8) ,
23888	 => std_logic_vector(to_unsigned(130,8) ,
23889	 => std_logic_vector(to_unsigned(133,8) ,
23890	 => std_logic_vector(to_unsigned(131,8) ,
23891	 => std_logic_vector(to_unsigned(133,8) ,
23892	 => std_logic_vector(to_unsigned(138,8) ,
23893	 => std_logic_vector(to_unsigned(134,8) ,
23894	 => std_logic_vector(to_unsigned(131,8) ,
23895	 => std_logic_vector(to_unsigned(134,8) ,
23896	 => std_logic_vector(to_unsigned(136,8) ,
23897	 => std_logic_vector(to_unsigned(134,8) ,
23898	 => std_logic_vector(to_unsigned(138,8) ,
23899	 => std_logic_vector(to_unsigned(136,8) ,
23900	 => std_logic_vector(to_unsigned(139,8) ,
23901	 => std_logic_vector(to_unsigned(134,8) ,
23902	 => std_logic_vector(to_unsigned(138,8) ,
23903	 => std_logic_vector(to_unsigned(116,8) ,
23904	 => std_logic_vector(to_unsigned(20,8) ,
23905	 => std_logic_vector(to_unsigned(8,8) ,
23906	 => std_logic_vector(to_unsigned(4,8) ,
23907	 => std_logic_vector(to_unsigned(3,8) ,
23908	 => std_logic_vector(to_unsigned(10,8) ,
23909	 => std_logic_vector(to_unsigned(17,8) ,
23910	 => std_logic_vector(to_unsigned(12,8) ,
23911	 => std_logic_vector(to_unsigned(5,8) ,
23912	 => std_logic_vector(to_unsigned(9,8) ,
23913	 => std_logic_vector(to_unsigned(13,8) ,
23914	 => std_logic_vector(to_unsigned(48,8) ,
23915	 => std_logic_vector(to_unsigned(159,8) ,
23916	 => std_logic_vector(to_unsigned(146,8) ,
23917	 => std_logic_vector(to_unsigned(141,8) ,
23918	 => std_logic_vector(to_unsigned(141,8) ,
23919	 => std_logic_vector(to_unsigned(141,8) ,
23920	 => std_logic_vector(to_unsigned(141,8) ,
23921	 => std_logic_vector(to_unsigned(128,8) ,
23922	 => std_logic_vector(to_unsigned(86,8) ,
23923	 => std_logic_vector(to_unsigned(100,8) ,
23924	 => std_logic_vector(to_unsigned(108,8) ,
23925	 => std_logic_vector(to_unsigned(96,8) ,
23926	 => std_logic_vector(to_unsigned(80,8) ,
23927	 => std_logic_vector(to_unsigned(51,8) ,
23928	 => std_logic_vector(to_unsigned(34,8) ,
23929	 => std_logic_vector(to_unsigned(27,8) ,
23930	 => std_logic_vector(to_unsigned(27,8) ,
23931	 => std_logic_vector(to_unsigned(13,8) ,
23932	 => std_logic_vector(to_unsigned(4,8) ,
23933	 => std_logic_vector(to_unsigned(3,8) ,
23934	 => std_logic_vector(to_unsigned(3,8) ,
23935	 => std_logic_vector(to_unsigned(7,8) ,
23936	 => std_logic_vector(to_unsigned(8,8) ,
23937	 => std_logic_vector(to_unsigned(4,8) ,
23938	 => std_logic_vector(to_unsigned(23,8) ,
23939	 => std_logic_vector(to_unsigned(152,8) ,
23940	 => std_logic_vector(to_unsigned(170,8) ,
23941	 => std_logic_vector(to_unsigned(157,8) ,
23942	 => std_logic_vector(to_unsigned(163,8) ,
23943	 => std_logic_vector(to_unsigned(163,8) ,
23944	 => std_logic_vector(to_unsigned(164,8) ,
23945	 => std_logic_vector(to_unsigned(164,8) ,
23946	 => std_logic_vector(to_unsigned(166,8) ,
23947	 => std_logic_vector(to_unsigned(159,8) ,
23948	 => std_logic_vector(to_unsigned(161,8) ,
23949	 => std_logic_vector(to_unsigned(163,8) ,
23950	 => std_logic_vector(to_unsigned(163,8) ,
23951	 => std_logic_vector(to_unsigned(161,8) ,
23952	 => std_logic_vector(to_unsigned(164,8) ,
23953	 => std_logic_vector(to_unsigned(154,8) ,
23954	 => std_logic_vector(to_unsigned(146,8) ,
23955	 => std_logic_vector(to_unsigned(133,8) ,
23956	 => std_logic_vector(to_unsigned(161,8) ,
23957	 => std_logic_vector(to_unsigned(62,8) ,
23958	 => std_logic_vector(to_unsigned(3,8) ,
23959	 => std_logic_vector(to_unsigned(4,8) ,
23960	 => std_logic_vector(to_unsigned(5,8) ,
23961	 => std_logic_vector(to_unsigned(11,8) ,
23962	 => std_logic_vector(to_unsigned(14,8) ,
23963	 => std_logic_vector(to_unsigned(11,8) ,
23964	 => std_logic_vector(to_unsigned(14,8) ,
23965	 => std_logic_vector(to_unsigned(19,8) ,
23966	 => std_logic_vector(to_unsigned(5,8) ,
23967	 => std_logic_vector(to_unsigned(45,8) ,
23968	 => std_logic_vector(to_unsigned(159,8) ,
23969	 => std_logic_vector(to_unsigned(130,8) ,
23970	 => std_logic_vector(to_unsigned(124,8) ,
23971	 => std_logic_vector(to_unsigned(119,8) ,
23972	 => std_logic_vector(to_unsigned(101,8) ,
23973	 => std_logic_vector(to_unsigned(104,8) ,
23974	 => std_logic_vector(to_unsigned(101,8) ,
23975	 => std_logic_vector(to_unsigned(90,8) ,
23976	 => std_logic_vector(to_unsigned(93,8) ,
23977	 => std_logic_vector(to_unsigned(101,8) ,
23978	 => std_logic_vector(to_unsigned(96,8) ,
23979	 => std_logic_vector(to_unsigned(92,8) ,
23980	 => std_logic_vector(to_unsigned(92,8) ,
23981	 => std_logic_vector(to_unsigned(96,8) ,
23982	 => std_logic_vector(to_unsigned(105,8) ,
23983	 => std_logic_vector(to_unsigned(107,8) ,
23984	 => std_logic_vector(to_unsigned(97,8) ,
23985	 => std_logic_vector(to_unsigned(97,8) ,
23986	 => std_logic_vector(to_unsigned(103,8) ,
23987	 => std_logic_vector(to_unsigned(105,8) ,
23988	 => std_logic_vector(to_unsigned(103,8) ,
23989	 => std_logic_vector(to_unsigned(104,8) ,
23990	 => std_logic_vector(to_unsigned(127,8) ,
23991	 => std_logic_vector(to_unsigned(161,8) ,
23992	 => std_logic_vector(to_unsigned(163,8) ,
23993	 => std_logic_vector(to_unsigned(138,8) ,
23994	 => std_logic_vector(to_unsigned(127,8) ,
23995	 => std_logic_vector(to_unsigned(121,8) ,
23996	 => std_logic_vector(to_unsigned(111,8) ,
23997	 => std_logic_vector(to_unsigned(116,8) ,
23998	 => std_logic_vector(to_unsigned(115,8) ,
23999	 => std_logic_vector(to_unsigned(111,8) ,
24000	 => std_logic_vector(to_unsigned(105,8) ,
24001	 => std_logic_vector(to_unsigned(166,8) ,
24002	 => std_logic_vector(to_unsigned(168,8) ,
24003	 => std_logic_vector(to_unsigned(168,8) ,
24004	 => std_logic_vector(to_unsigned(163,8) ,
24005	 => std_logic_vector(to_unsigned(161,8) ,
24006	 => std_logic_vector(to_unsigned(166,8) ,
24007	 => std_logic_vector(to_unsigned(119,8) ,
24008	 => std_logic_vector(to_unsigned(49,8) ,
24009	 => std_logic_vector(to_unsigned(23,8) ,
24010	 => std_logic_vector(to_unsigned(20,8) ,
24011	 => std_logic_vector(to_unsigned(49,8) ,
24012	 => std_logic_vector(to_unsigned(13,8) ,
24013	 => std_logic_vector(to_unsigned(2,8) ,
24014	 => std_logic_vector(to_unsigned(3,8) ,
24015	 => std_logic_vector(to_unsigned(7,8) ,
24016	 => std_logic_vector(to_unsigned(5,8) ,
24017	 => std_logic_vector(to_unsigned(52,8) ,
24018	 => std_logic_vector(to_unsigned(37,8) ,
24019	 => std_logic_vector(to_unsigned(33,8) ,
24020	 => std_logic_vector(to_unsigned(34,8) ,
24021	 => std_logic_vector(to_unsigned(40,8) ,
24022	 => std_logic_vector(to_unsigned(96,8) ,
24023	 => std_logic_vector(to_unsigned(67,8) ,
24024	 => std_logic_vector(to_unsigned(25,8) ,
24025	 => std_logic_vector(to_unsigned(4,8) ,
24026	 => std_logic_vector(to_unsigned(2,8) ,
24027	 => std_logic_vector(to_unsigned(4,8) ,
24028	 => std_logic_vector(to_unsigned(3,8) ,
24029	 => std_logic_vector(to_unsigned(1,8) ,
24030	 => std_logic_vector(to_unsigned(2,8) ,
24031	 => std_logic_vector(to_unsigned(8,8) ,
24032	 => std_logic_vector(to_unsigned(8,8) ,
24033	 => std_logic_vector(to_unsigned(4,8) ,
24034	 => std_logic_vector(to_unsigned(2,8) ,
24035	 => std_logic_vector(to_unsigned(19,8) ,
24036	 => std_logic_vector(to_unsigned(57,8) ,
24037	 => std_logic_vector(to_unsigned(42,8) ,
24038	 => std_logic_vector(to_unsigned(3,8) ,
24039	 => std_logic_vector(to_unsigned(1,8) ,
24040	 => std_logic_vector(to_unsigned(3,8) ,
24041	 => std_logic_vector(to_unsigned(7,8) ,
24042	 => std_logic_vector(to_unsigned(7,8) ,
24043	 => std_logic_vector(to_unsigned(17,8) ,
24044	 => std_logic_vector(to_unsigned(25,8) ,
24045	 => std_logic_vector(to_unsigned(19,8) ,
24046	 => std_logic_vector(to_unsigned(6,8) ,
24047	 => std_logic_vector(to_unsigned(5,8) ,
24048	 => std_logic_vector(to_unsigned(4,8) ,
24049	 => std_logic_vector(to_unsigned(2,8) ,
24050	 => std_logic_vector(to_unsigned(29,8) ,
24051	 => std_logic_vector(to_unsigned(171,8) ,
24052	 => std_logic_vector(to_unsigned(170,8) ,
24053	 => std_logic_vector(to_unsigned(157,8) ,
24054	 => std_logic_vector(to_unsigned(154,8) ,
24055	 => std_logic_vector(to_unsigned(164,8) ,
24056	 => std_logic_vector(to_unsigned(125,8) ,
24057	 => std_logic_vector(to_unsigned(10,8) ,
24058	 => std_logic_vector(to_unsigned(3,8) ,
24059	 => std_logic_vector(to_unsigned(4,8) ,
24060	 => std_logic_vector(to_unsigned(5,8) ,
24061	 => std_logic_vector(to_unsigned(14,8) ,
24062	 => std_logic_vector(to_unsigned(7,8) ,
24063	 => std_logic_vector(to_unsigned(4,8) ,
24064	 => std_logic_vector(to_unsigned(3,8) ,
24065	 => std_logic_vector(to_unsigned(4,8) ,
24066	 => std_logic_vector(to_unsigned(3,8) ,
24067	 => std_logic_vector(to_unsigned(1,8) ,
24068	 => std_logic_vector(to_unsigned(2,8) ,
24069	 => std_logic_vector(to_unsigned(4,8) ,
24070	 => std_logic_vector(to_unsigned(4,8) ,
24071	 => std_logic_vector(to_unsigned(11,8) ,
24072	 => std_logic_vector(to_unsigned(6,8) ,
24073	 => std_logic_vector(to_unsigned(1,8) ,
24074	 => std_logic_vector(to_unsigned(43,8) ,
24075	 => std_logic_vector(to_unsigned(112,8) ,
24076	 => std_logic_vector(to_unsigned(7,8) ,
24077	 => std_logic_vector(to_unsigned(8,8) ,
24078	 => std_logic_vector(to_unsigned(44,8) ,
24079	 => std_logic_vector(to_unsigned(41,8) ,
24080	 => std_logic_vector(to_unsigned(8,8) ,
24081	 => std_logic_vector(to_unsigned(3,8) ,
24082	 => std_logic_vector(to_unsigned(5,8) ,
24083	 => std_logic_vector(to_unsigned(17,8) ,
24084	 => std_logic_vector(to_unsigned(27,8) ,
24085	 => std_logic_vector(to_unsigned(27,8) ,
24086	 => std_logic_vector(to_unsigned(25,8) ,
24087	 => std_logic_vector(to_unsigned(64,8) ,
24088	 => std_logic_vector(to_unsigned(118,8) ,
24089	 => std_logic_vector(to_unsigned(108,8) ,
24090	 => std_logic_vector(to_unsigned(130,8) ,
24091	 => std_logic_vector(to_unsigned(138,8) ,
24092	 => std_logic_vector(to_unsigned(152,8) ,
24093	 => std_logic_vector(to_unsigned(166,8) ,
24094	 => std_logic_vector(to_unsigned(164,8) ,
24095	 => std_logic_vector(to_unsigned(161,8) ,
24096	 => std_logic_vector(to_unsigned(161,8) ,
24097	 => std_logic_vector(to_unsigned(163,8) ,
24098	 => std_logic_vector(to_unsigned(170,8) ,
24099	 => std_logic_vector(to_unsigned(163,8) ,
24100	 => std_logic_vector(to_unsigned(161,8) ,
24101	 => std_logic_vector(to_unsigned(166,8) ,
24102	 => std_logic_vector(to_unsigned(144,8) ,
24103	 => std_logic_vector(to_unsigned(99,8) ,
24104	 => std_logic_vector(to_unsigned(136,8) ,
24105	 => std_logic_vector(to_unsigned(144,8) ,
24106	 => std_logic_vector(to_unsigned(133,8) ,
24107	 => std_logic_vector(to_unsigned(146,8) ,
24108	 => std_logic_vector(to_unsigned(147,8) ,
24109	 => std_logic_vector(to_unsigned(127,8) ,
24110	 => std_logic_vector(to_unsigned(146,8) ,
24111	 => std_logic_vector(to_unsigned(159,8) ,
24112	 => std_logic_vector(to_unsigned(156,8) ,
24113	 => std_logic_vector(to_unsigned(147,8) ,
24114	 => std_logic_vector(to_unsigned(115,8) ,
24115	 => std_logic_vector(to_unsigned(12,8) ,
24116	 => std_logic_vector(to_unsigned(2,8) ,
24117	 => std_logic_vector(to_unsigned(24,8) ,
24118	 => std_logic_vector(to_unsigned(6,8) ,
24119	 => std_logic_vector(to_unsigned(2,8) ,
24120	 => std_logic_vector(to_unsigned(6,8) ,
24121	 => std_logic_vector(to_unsigned(6,8) ,
24122	 => std_logic_vector(to_unsigned(3,8) ,
24123	 => std_logic_vector(to_unsigned(4,8) ,
24124	 => std_logic_vector(to_unsigned(4,8) ,
24125	 => std_logic_vector(to_unsigned(16,8) ,
24126	 => std_logic_vector(to_unsigned(14,8) ,
24127	 => std_logic_vector(to_unsigned(6,8) ,
24128	 => std_logic_vector(to_unsigned(11,8) ,
24129	 => std_logic_vector(to_unsigned(13,8) ,
24130	 => std_logic_vector(to_unsigned(22,8) ,
24131	 => std_logic_vector(to_unsigned(90,8) ,
24132	 => std_logic_vector(to_unsigned(161,8) ,
24133	 => std_logic_vector(to_unsigned(161,8) ,
24134	 => std_logic_vector(to_unsigned(157,8) ,
24135	 => std_logic_vector(to_unsigned(156,8) ,
24136	 => std_logic_vector(to_unsigned(154,8) ,
24137	 => std_logic_vector(to_unsigned(156,8) ,
24138	 => std_logic_vector(to_unsigned(149,8) ,
24139	 => std_logic_vector(to_unsigned(136,8) ,
24140	 => std_logic_vector(to_unsigned(142,8) ,
24141	 => std_logic_vector(to_unsigned(144,8) ,
24142	 => std_logic_vector(to_unsigned(134,8) ,
24143	 => std_logic_vector(to_unsigned(45,8) ,
24144	 => std_logic_vector(to_unsigned(4,8) ,
24145	 => std_logic_vector(to_unsigned(8,8) ,
24146	 => std_logic_vector(to_unsigned(6,8) ,
24147	 => std_logic_vector(to_unsigned(3,8) ,
24148	 => std_logic_vector(to_unsigned(24,8) ,
24149	 => std_logic_vector(to_unsigned(35,8) ,
24150	 => std_logic_vector(to_unsigned(6,8) ,
24151	 => std_logic_vector(to_unsigned(7,8) ,
24152	 => std_logic_vector(to_unsigned(15,8) ,
24153	 => std_logic_vector(to_unsigned(22,8) ,
24154	 => std_logic_vector(to_unsigned(22,8) ,
24155	 => std_logic_vector(to_unsigned(44,8) ,
24156	 => std_logic_vector(to_unsigned(88,8) ,
24157	 => std_logic_vector(to_unsigned(107,8) ,
24158	 => std_logic_vector(to_unsigned(125,8) ,
24159	 => std_logic_vector(to_unsigned(152,8) ,
24160	 => std_logic_vector(to_unsigned(141,8) ,
24161	 => std_logic_vector(to_unsigned(128,8) ,
24162	 => std_logic_vector(to_unsigned(130,8) ,
24163	 => std_logic_vector(to_unsigned(111,8) ,
24164	 => std_logic_vector(to_unsigned(27,8) ,
24165	 => std_logic_vector(to_unsigned(7,8) ,
24166	 => std_logic_vector(to_unsigned(13,8) ,
24167	 => std_logic_vector(to_unsigned(12,8) ,
24168	 => std_logic_vector(to_unsigned(9,8) ,
24169	 => std_logic_vector(to_unsigned(8,8) ,
24170	 => std_logic_vector(to_unsigned(5,8) ,
24171	 => std_logic_vector(to_unsigned(3,8) ,
24172	 => std_logic_vector(to_unsigned(4,8) ,
24173	 => std_logic_vector(to_unsigned(7,8) ,
24174	 => std_logic_vector(to_unsigned(13,8) ,
24175	 => std_logic_vector(to_unsigned(9,8) ,
24176	 => std_logic_vector(to_unsigned(15,8) ,
24177	 => std_logic_vector(to_unsigned(27,8) ,
24178	 => std_logic_vector(to_unsigned(27,8) ,
24179	 => std_logic_vector(to_unsigned(38,8) ,
24180	 => std_logic_vector(to_unsigned(27,8) ,
24181	 => std_logic_vector(to_unsigned(12,8) ,
24182	 => std_logic_vector(to_unsigned(13,8) ,
24183	 => std_logic_vector(to_unsigned(18,8) ,
24184	 => std_logic_vector(to_unsigned(29,8) ,
24185	 => std_logic_vector(to_unsigned(29,8) ,
24186	 => std_logic_vector(to_unsigned(20,8) ,
24187	 => std_logic_vector(to_unsigned(41,8) ,
24188	 => std_logic_vector(to_unsigned(96,8) ,
24189	 => std_logic_vector(to_unsigned(124,8) ,
24190	 => std_logic_vector(to_unsigned(119,8) ,
24191	 => std_logic_vector(to_unsigned(112,8) ,
24192	 => std_logic_vector(to_unsigned(109,8) ,
24193	 => std_logic_vector(to_unsigned(112,8) ,
24194	 => std_logic_vector(to_unsigned(23,8) ,
24195	 => std_logic_vector(to_unsigned(2,8) ,
24196	 => std_logic_vector(to_unsigned(3,8) ,
24197	 => std_logic_vector(to_unsigned(5,8) ,
24198	 => std_logic_vector(to_unsigned(6,8) ,
24199	 => std_logic_vector(to_unsigned(17,8) ,
24200	 => std_logic_vector(to_unsigned(29,8) ,
24201	 => std_logic_vector(to_unsigned(16,8) ,
24202	 => std_logic_vector(to_unsigned(18,8) ,
24203	 => std_logic_vector(to_unsigned(13,8) ,
24204	 => std_logic_vector(to_unsigned(3,8) ,
24205	 => std_logic_vector(to_unsigned(23,8) ,
24206	 => std_logic_vector(to_unsigned(133,8) ,
24207	 => std_logic_vector(to_unsigned(146,8) ,
24208	 => std_logic_vector(to_unsigned(130,8) ,
24209	 => std_logic_vector(to_unsigned(131,8) ,
24210	 => std_logic_vector(to_unsigned(133,8) ,
24211	 => std_logic_vector(to_unsigned(131,8) ,
24212	 => std_logic_vector(to_unsigned(134,8) ,
24213	 => std_logic_vector(to_unsigned(138,8) ,
24214	 => std_logic_vector(to_unsigned(139,8) ,
24215	 => std_logic_vector(to_unsigned(138,8) ,
24216	 => std_logic_vector(to_unsigned(139,8) ,
24217	 => std_logic_vector(to_unsigned(142,8) ,
24218	 => std_logic_vector(to_unsigned(144,8) ,
24219	 => std_logic_vector(to_unsigned(141,8) ,
24220	 => std_logic_vector(to_unsigned(138,8) ,
24221	 => std_logic_vector(to_unsigned(131,8) ,
24222	 => std_logic_vector(to_unsigned(138,8) ,
24223	 => std_logic_vector(to_unsigned(119,8) ,
24224	 => std_logic_vector(to_unsigned(43,8) ,
24225	 => std_logic_vector(to_unsigned(30,8) ,
24226	 => std_logic_vector(to_unsigned(15,8) ,
24227	 => std_logic_vector(to_unsigned(13,8) ,
24228	 => std_logic_vector(to_unsigned(17,8) ,
24229	 => std_logic_vector(to_unsigned(10,8) ,
24230	 => std_logic_vector(to_unsigned(8,8) ,
24231	 => std_logic_vector(to_unsigned(7,8) ,
24232	 => std_logic_vector(to_unsigned(5,8) ,
24233	 => std_logic_vector(to_unsigned(23,8) ,
24234	 => std_logic_vector(to_unsigned(136,8) ,
24235	 => std_logic_vector(to_unsigned(161,8) ,
24236	 => std_logic_vector(to_unsigned(147,8) ,
24237	 => std_logic_vector(to_unsigned(146,8) ,
24238	 => std_logic_vector(to_unsigned(144,8) ,
24239	 => std_logic_vector(to_unsigned(142,8) ,
24240	 => std_logic_vector(to_unsigned(138,8) ,
24241	 => std_logic_vector(to_unsigned(125,8) ,
24242	 => std_logic_vector(to_unsigned(65,8) ,
24243	 => std_logic_vector(to_unsigned(40,8) ,
24244	 => std_logic_vector(to_unsigned(29,8) ,
24245	 => std_logic_vector(to_unsigned(18,8) ,
24246	 => std_logic_vector(to_unsigned(15,8) ,
24247	 => std_logic_vector(to_unsigned(16,8) ,
24248	 => std_logic_vector(to_unsigned(27,8) ,
24249	 => std_logic_vector(to_unsigned(42,8) ,
24250	 => std_logic_vector(to_unsigned(18,8) ,
24251	 => std_logic_vector(to_unsigned(1,8) ,
24252	 => std_logic_vector(to_unsigned(0,8) ,
24253	 => std_logic_vector(to_unsigned(0,8) ,
24254	 => std_logic_vector(to_unsigned(3,8) ,
24255	 => std_logic_vector(to_unsigned(6,8) ,
24256	 => std_logic_vector(to_unsigned(5,8) ,
24257	 => std_logic_vector(to_unsigned(9,8) ,
24258	 => std_logic_vector(to_unsigned(93,8) ,
24259	 => std_logic_vector(to_unsigned(186,8) ,
24260	 => std_logic_vector(to_unsigned(159,8) ,
24261	 => std_logic_vector(to_unsigned(166,8) ,
24262	 => std_logic_vector(to_unsigned(164,8) ,
24263	 => std_logic_vector(to_unsigned(166,8) ,
24264	 => std_logic_vector(to_unsigned(166,8) ,
24265	 => std_logic_vector(to_unsigned(166,8) ,
24266	 => std_logic_vector(to_unsigned(166,8) ,
24267	 => std_logic_vector(to_unsigned(164,8) ,
24268	 => std_logic_vector(to_unsigned(164,8) ,
24269	 => std_logic_vector(to_unsigned(159,8) ,
24270	 => std_logic_vector(to_unsigned(164,8) ,
24271	 => std_logic_vector(to_unsigned(157,8) ,
24272	 => std_logic_vector(to_unsigned(156,8) ,
24273	 => std_logic_vector(to_unsigned(151,8) ,
24274	 => std_logic_vector(to_unsigned(151,8) ,
24275	 => std_logic_vector(to_unsigned(163,8) ,
24276	 => std_logic_vector(to_unsigned(141,8) ,
24277	 => std_logic_vector(to_unsigned(77,8) ,
24278	 => std_logic_vector(to_unsigned(4,8) ,
24279	 => std_logic_vector(to_unsigned(3,8) ,
24280	 => std_logic_vector(to_unsigned(5,8) ,
24281	 => std_logic_vector(to_unsigned(14,8) ,
24282	 => std_logic_vector(to_unsigned(23,8) ,
24283	 => std_logic_vector(to_unsigned(12,8) ,
24284	 => std_logic_vector(to_unsigned(9,8) ,
24285	 => std_logic_vector(to_unsigned(25,8) ,
24286	 => std_logic_vector(to_unsigned(6,8) ,
24287	 => std_logic_vector(to_unsigned(26,8) ,
24288	 => std_logic_vector(to_unsigned(144,8) ,
24289	 => std_logic_vector(to_unsigned(74,8) ,
24290	 => std_logic_vector(to_unsigned(99,8) ,
24291	 => std_logic_vector(to_unsigned(119,8) ,
24292	 => std_logic_vector(to_unsigned(114,8) ,
24293	 => std_logic_vector(to_unsigned(111,8) ,
24294	 => std_logic_vector(to_unsigned(103,8) ,
24295	 => std_logic_vector(to_unsigned(104,8) ,
24296	 => std_logic_vector(to_unsigned(105,8) ,
24297	 => std_logic_vector(to_unsigned(105,8) ,
24298	 => std_logic_vector(to_unsigned(107,8) ,
24299	 => std_logic_vector(to_unsigned(91,8) ,
24300	 => std_logic_vector(to_unsigned(96,8) ,
24301	 => std_logic_vector(to_unsigned(104,8) ,
24302	 => std_logic_vector(to_unsigned(101,8) ,
24303	 => std_logic_vector(to_unsigned(108,8) ,
24304	 => std_logic_vector(to_unsigned(114,8) ,
24305	 => std_logic_vector(to_unsigned(104,8) ,
24306	 => std_logic_vector(to_unsigned(104,8) ,
24307	 => std_logic_vector(to_unsigned(109,8) ,
24308	 => std_logic_vector(to_unsigned(105,8) ,
24309	 => std_logic_vector(to_unsigned(104,8) ,
24310	 => std_logic_vector(to_unsigned(109,8) ,
24311	 => std_logic_vector(to_unsigned(146,8) ,
24312	 => std_logic_vector(to_unsigned(170,8) ,
24313	 => std_logic_vector(to_unsigned(161,8) ,
24314	 => std_logic_vector(to_unsigned(133,8) ,
24315	 => std_logic_vector(to_unsigned(124,8) ,
24316	 => std_logic_vector(to_unsigned(124,8) ,
24317	 => std_logic_vector(to_unsigned(114,8) ,
24318	 => std_logic_vector(to_unsigned(112,8) ,
24319	 => std_logic_vector(to_unsigned(115,8) ,
24320	 => std_logic_vector(to_unsigned(112,8) ,
24321	 => std_logic_vector(to_unsigned(163,8) ,
24322	 => std_logic_vector(to_unsigned(164,8) ,
24323	 => std_logic_vector(to_unsigned(164,8) ,
24324	 => std_logic_vector(to_unsigned(161,8) ,
24325	 => std_logic_vector(to_unsigned(161,8) ,
24326	 => std_logic_vector(to_unsigned(164,8) ,
24327	 => std_logic_vector(to_unsigned(103,8) ,
24328	 => std_logic_vector(to_unsigned(69,8) ,
24329	 => std_logic_vector(to_unsigned(71,8) ,
24330	 => std_logic_vector(to_unsigned(51,8) ,
24331	 => std_logic_vector(to_unsigned(35,8) ,
24332	 => std_logic_vector(to_unsigned(26,8) ,
24333	 => std_logic_vector(to_unsigned(7,8) ,
24334	 => std_logic_vector(to_unsigned(1,8) ,
24335	 => std_logic_vector(to_unsigned(4,8) ,
24336	 => std_logic_vector(to_unsigned(3,8) ,
24337	 => std_logic_vector(to_unsigned(39,8) ,
24338	 => std_logic_vector(to_unsigned(41,8) ,
24339	 => std_logic_vector(to_unsigned(11,8) ,
24340	 => std_logic_vector(to_unsigned(53,8) ,
24341	 => std_logic_vector(to_unsigned(84,8) ,
24342	 => std_logic_vector(to_unsigned(36,8) ,
24343	 => std_logic_vector(to_unsigned(81,8) ,
24344	 => std_logic_vector(to_unsigned(171,8) ,
24345	 => std_logic_vector(to_unsigned(112,8) ,
24346	 => std_logic_vector(to_unsigned(10,8) ,
24347	 => std_logic_vector(to_unsigned(2,8) ,
24348	 => std_logic_vector(to_unsigned(2,8) ,
24349	 => std_logic_vector(to_unsigned(1,8) ,
24350	 => std_logic_vector(to_unsigned(3,8) ,
24351	 => std_logic_vector(to_unsigned(7,8) ,
24352	 => std_logic_vector(to_unsigned(8,8) ,
24353	 => std_logic_vector(to_unsigned(3,8) ,
24354	 => std_logic_vector(to_unsigned(1,8) ,
24355	 => std_logic_vector(to_unsigned(9,8) ,
24356	 => std_logic_vector(to_unsigned(63,8) ,
24357	 => std_logic_vector(to_unsigned(22,8) ,
24358	 => std_logic_vector(to_unsigned(2,8) ,
24359	 => std_logic_vector(to_unsigned(2,8) ,
24360	 => std_logic_vector(to_unsigned(1,8) ,
24361	 => std_logic_vector(to_unsigned(15,8) ,
24362	 => std_logic_vector(to_unsigned(41,8) ,
24363	 => std_logic_vector(to_unsigned(35,8) ,
24364	 => std_logic_vector(to_unsigned(42,8) ,
24365	 => std_logic_vector(to_unsigned(39,8) ,
24366	 => std_logic_vector(to_unsigned(17,8) ,
24367	 => std_logic_vector(to_unsigned(5,8) ,
24368	 => std_logic_vector(to_unsigned(0,8) ,
24369	 => std_logic_vector(to_unsigned(0,8) ,
24370	 => std_logic_vector(to_unsigned(31,8) ,
24371	 => std_logic_vector(to_unsigned(183,8) ,
24372	 => std_logic_vector(to_unsigned(163,8) ,
24373	 => std_logic_vector(to_unsigned(156,8) ,
24374	 => std_logic_vector(to_unsigned(151,8) ,
24375	 => std_logic_vector(to_unsigned(170,8) ,
24376	 => std_logic_vector(to_unsigned(138,8) ,
24377	 => std_logic_vector(to_unsigned(18,8) ,
24378	 => std_logic_vector(to_unsigned(5,8) ,
24379	 => std_logic_vector(to_unsigned(6,8) ,
24380	 => std_logic_vector(to_unsigned(5,8) ,
24381	 => std_logic_vector(to_unsigned(9,8) ,
24382	 => std_logic_vector(to_unsigned(7,8) ,
24383	 => std_logic_vector(to_unsigned(7,8) ,
24384	 => std_logic_vector(to_unsigned(5,8) ,
24385	 => std_logic_vector(to_unsigned(4,8) ,
24386	 => std_logic_vector(to_unsigned(4,8) ,
24387	 => std_logic_vector(to_unsigned(2,8) ,
24388	 => std_logic_vector(to_unsigned(3,8) ,
24389	 => std_logic_vector(to_unsigned(4,8) ,
24390	 => std_logic_vector(to_unsigned(4,8) ,
24391	 => std_logic_vector(to_unsigned(9,8) ,
24392	 => std_logic_vector(to_unsigned(7,8) ,
24393	 => std_logic_vector(to_unsigned(1,8) ,
24394	 => std_logic_vector(to_unsigned(14,8) ,
24395	 => std_logic_vector(to_unsigned(82,8) ,
24396	 => std_logic_vector(to_unsigned(37,8) ,
24397	 => std_logic_vector(to_unsigned(15,8) ,
24398	 => std_logic_vector(to_unsigned(103,8) ,
24399	 => std_logic_vector(to_unsigned(184,8) ,
24400	 => std_logic_vector(to_unsigned(136,8) ,
24401	 => std_logic_vector(to_unsigned(30,8) ,
24402	 => std_logic_vector(to_unsigned(2,8) ,
24403	 => std_logic_vector(to_unsigned(13,8) ,
24404	 => std_logic_vector(to_unsigned(37,8) ,
24405	 => std_logic_vector(to_unsigned(24,8) ,
24406	 => std_logic_vector(to_unsigned(17,8) ,
24407	 => std_logic_vector(to_unsigned(25,8) ,
24408	 => std_logic_vector(to_unsigned(81,8) ,
24409	 => std_logic_vector(to_unsigned(92,8) ,
24410	 => std_logic_vector(to_unsigned(121,8) ,
24411	 => std_logic_vector(to_unsigned(147,8) ,
24412	 => std_logic_vector(to_unsigned(156,8) ,
24413	 => std_logic_vector(to_unsigned(161,8) ,
24414	 => std_logic_vector(to_unsigned(164,8) ,
24415	 => std_logic_vector(to_unsigned(166,8) ,
24416	 => std_logic_vector(to_unsigned(164,8) ,
24417	 => std_logic_vector(to_unsigned(161,8) ,
24418	 => std_logic_vector(to_unsigned(168,8) ,
24419	 => std_logic_vector(to_unsigned(163,8) ,
24420	 => std_logic_vector(to_unsigned(161,8) ,
24421	 => std_logic_vector(to_unsigned(168,8) ,
24422	 => std_logic_vector(to_unsigned(109,8) ,
24423	 => std_logic_vector(to_unsigned(77,8) ,
24424	 => std_logic_vector(to_unsigned(147,8) ,
24425	 => std_logic_vector(to_unsigned(133,8) ,
24426	 => std_logic_vector(to_unsigned(124,8) ,
24427	 => std_logic_vector(to_unsigned(154,8) ,
24428	 => std_logic_vector(to_unsigned(157,8) ,
24429	 => std_logic_vector(to_unsigned(118,8) ,
24430	 => std_logic_vector(to_unsigned(115,8) ,
24431	 => std_logic_vector(to_unsigned(133,8) ,
24432	 => std_logic_vector(to_unsigned(131,8) ,
24433	 => std_logic_vector(to_unsigned(97,8) ,
24434	 => std_logic_vector(to_unsigned(45,8) ,
24435	 => std_logic_vector(to_unsigned(3,8) ,
24436	 => std_logic_vector(to_unsigned(6,8) ,
24437	 => std_logic_vector(to_unsigned(28,8) ,
24438	 => std_logic_vector(to_unsigned(1,8) ,
24439	 => std_logic_vector(to_unsigned(1,8) ,
24440	 => std_logic_vector(to_unsigned(5,8) ,
24441	 => std_logic_vector(to_unsigned(13,8) ,
24442	 => std_logic_vector(to_unsigned(19,8) ,
24443	 => std_logic_vector(to_unsigned(15,8) ,
24444	 => std_logic_vector(to_unsigned(9,8) ,
24445	 => std_logic_vector(to_unsigned(23,8) ,
24446	 => std_logic_vector(to_unsigned(16,8) ,
24447	 => std_logic_vector(to_unsigned(3,8) ,
24448	 => std_logic_vector(to_unsigned(6,8) ,
24449	 => std_logic_vector(to_unsigned(8,8) ,
24450	 => std_logic_vector(to_unsigned(22,8) ,
24451	 => std_logic_vector(to_unsigned(93,8) ,
24452	 => std_logic_vector(to_unsigned(130,8) ,
24453	 => std_logic_vector(to_unsigned(154,8) ,
24454	 => std_logic_vector(to_unsigned(166,8) ,
24455	 => std_logic_vector(to_unsigned(154,8) ,
24456	 => std_logic_vector(to_unsigned(146,8) ,
24457	 => std_logic_vector(to_unsigned(152,8) ,
24458	 => std_logic_vector(to_unsigned(147,8) ,
24459	 => std_logic_vector(to_unsigned(142,8) ,
24460	 => std_logic_vector(to_unsigned(139,8) ,
24461	 => std_logic_vector(to_unsigned(86,8) ,
24462	 => std_logic_vector(to_unsigned(45,8) ,
24463	 => std_logic_vector(to_unsigned(11,8) ,
24464	 => std_logic_vector(to_unsigned(4,8) ,
24465	 => std_logic_vector(to_unsigned(4,8) ,
24466	 => std_logic_vector(to_unsigned(11,8) ,
24467	 => std_logic_vector(to_unsigned(6,8) ,
24468	 => std_logic_vector(to_unsigned(17,8) ,
24469	 => std_logic_vector(to_unsigned(41,8) ,
24470	 => std_logic_vector(to_unsigned(8,8) ,
24471	 => std_logic_vector(to_unsigned(6,8) ,
24472	 => std_logic_vector(to_unsigned(17,8) ,
24473	 => std_logic_vector(to_unsigned(25,8) ,
24474	 => std_logic_vector(to_unsigned(12,8) ,
24475	 => std_logic_vector(to_unsigned(21,8) ,
24476	 => std_logic_vector(to_unsigned(45,8) ,
24477	 => std_logic_vector(to_unsigned(69,8) ,
24478	 => std_logic_vector(to_unsigned(109,8) ,
24479	 => std_logic_vector(to_unsigned(142,8) ,
24480	 => std_logic_vector(to_unsigned(149,8) ,
24481	 => std_logic_vector(to_unsigned(136,8) ,
24482	 => std_logic_vector(to_unsigned(151,8) ,
24483	 => std_logic_vector(to_unsigned(59,8) ,
24484	 => std_logic_vector(to_unsigned(8,8) ,
24485	 => std_logic_vector(to_unsigned(10,8) ,
24486	 => std_logic_vector(to_unsigned(17,8) ,
24487	 => std_logic_vector(to_unsigned(18,8) ,
24488	 => std_logic_vector(to_unsigned(10,8) ,
24489	 => std_logic_vector(to_unsigned(7,8) ,
24490	 => std_logic_vector(to_unsigned(8,8) ,
24491	 => std_logic_vector(to_unsigned(5,8) ,
24492	 => std_logic_vector(to_unsigned(5,8) ,
24493	 => std_logic_vector(to_unsigned(3,8) ,
24494	 => std_logic_vector(to_unsigned(6,8) ,
24495	 => std_logic_vector(to_unsigned(14,8) ,
24496	 => std_logic_vector(to_unsigned(23,8) ,
24497	 => std_logic_vector(to_unsigned(36,8) ,
24498	 => std_logic_vector(to_unsigned(35,8) ,
24499	 => std_logic_vector(to_unsigned(35,8) ,
24500	 => std_logic_vector(to_unsigned(29,8) ,
24501	 => std_logic_vector(to_unsigned(15,8) ,
24502	 => std_logic_vector(to_unsigned(11,8) ,
24503	 => std_logic_vector(to_unsigned(10,8) ,
24504	 => std_logic_vector(to_unsigned(13,8) ,
24505	 => std_logic_vector(to_unsigned(21,8) ,
24506	 => std_logic_vector(to_unsigned(18,8) ,
24507	 => std_logic_vector(to_unsigned(24,8) ,
24508	 => std_logic_vector(to_unsigned(69,8) ,
24509	 => std_logic_vector(to_unsigned(125,8) ,
24510	 => std_logic_vector(to_unsigned(116,8) ,
24511	 => std_logic_vector(to_unsigned(116,8) ,
24512	 => std_logic_vector(to_unsigned(114,8) ,
24513	 => std_logic_vector(to_unsigned(136,8) ,
24514	 => std_logic_vector(to_unsigned(57,8) ,
24515	 => std_logic_vector(to_unsigned(8,8) ,
24516	 => std_logic_vector(to_unsigned(6,8) ,
24517	 => std_logic_vector(to_unsigned(7,8) ,
24518	 => std_logic_vector(to_unsigned(8,8) ,
24519	 => std_logic_vector(to_unsigned(6,8) ,
24520	 => std_logic_vector(to_unsigned(5,8) ,
24521	 => std_logic_vector(to_unsigned(1,8) ,
24522	 => std_logic_vector(to_unsigned(6,8) ,
24523	 => std_logic_vector(to_unsigned(7,8) ,
24524	 => std_logic_vector(to_unsigned(3,8) ,
24525	 => std_logic_vector(to_unsigned(49,8) ,
24526	 => std_logic_vector(to_unsigned(157,8) ,
24527	 => std_logic_vector(to_unsigned(157,8) ,
24528	 => std_logic_vector(to_unsigned(149,8) ,
24529	 => std_logic_vector(to_unsigned(139,8) ,
24530	 => std_logic_vector(to_unsigned(133,8) ,
24531	 => std_logic_vector(to_unsigned(131,8) ,
24532	 => std_logic_vector(to_unsigned(138,8) ,
24533	 => std_logic_vector(to_unsigned(139,8) ,
24534	 => std_logic_vector(to_unsigned(139,8) ,
24535	 => std_logic_vector(to_unsigned(141,8) ,
24536	 => std_logic_vector(to_unsigned(139,8) ,
24537	 => std_logic_vector(to_unsigned(141,8) ,
24538	 => std_logic_vector(to_unsigned(139,8) ,
24539	 => std_logic_vector(to_unsigned(136,8) ,
24540	 => std_logic_vector(to_unsigned(136,8) ,
24541	 => std_logic_vector(to_unsigned(133,8) ,
24542	 => std_logic_vector(to_unsigned(157,8) ,
24543	 => std_logic_vector(to_unsigned(82,8) ,
24544	 => std_logic_vector(to_unsigned(25,8) ,
24545	 => std_logic_vector(to_unsigned(14,8) ,
24546	 => std_logic_vector(to_unsigned(4,8) ,
24547	 => std_logic_vector(to_unsigned(8,8) ,
24548	 => std_logic_vector(to_unsigned(7,8) ,
24549	 => std_logic_vector(to_unsigned(7,8) ,
24550	 => std_logic_vector(to_unsigned(8,8) ,
24551	 => std_logic_vector(to_unsigned(8,8) ,
24552	 => std_logic_vector(to_unsigned(2,8) ,
24553	 => std_logic_vector(to_unsigned(12,8) ,
24554	 => std_logic_vector(to_unsigned(131,8) ,
24555	 => std_logic_vector(to_unsigned(164,8) ,
24556	 => std_logic_vector(to_unsigned(156,8) ,
24557	 => std_logic_vector(to_unsigned(154,8) ,
24558	 => std_logic_vector(to_unsigned(146,8) ,
24559	 => std_logic_vector(to_unsigned(147,8) ,
24560	 => std_logic_vector(to_unsigned(139,8) ,
24561	 => std_logic_vector(to_unsigned(118,8) ,
24562	 => std_logic_vector(to_unsigned(107,8) ,
24563	 => std_logic_vector(to_unsigned(101,8) ,
24564	 => std_logic_vector(to_unsigned(108,8) ,
24565	 => std_logic_vector(to_unsigned(122,8) ,
24566	 => std_logic_vector(to_unsigned(124,8) ,
24567	 => std_logic_vector(to_unsigned(127,8) ,
24568	 => std_logic_vector(to_unsigned(105,8) ,
24569	 => std_logic_vector(to_unsigned(32,8) ,
24570	 => std_logic_vector(to_unsigned(5,8) ,
24571	 => std_logic_vector(to_unsigned(1,8) ,
24572	 => std_logic_vector(to_unsigned(1,8) ,
24573	 => std_logic_vector(to_unsigned(1,8) ,
24574	 => std_logic_vector(to_unsigned(8,8) ,
24575	 => std_logic_vector(to_unsigned(10,8) ,
24576	 => std_logic_vector(to_unsigned(4,8) ,
24577	 => std_logic_vector(to_unsigned(5,8) ,
24578	 => std_logic_vector(to_unsigned(47,8) ,
24579	 => std_logic_vector(to_unsigned(177,8) ,
24580	 => std_logic_vector(to_unsigned(164,8) ,
24581	 => std_logic_vector(to_unsigned(163,8) ,
24582	 => std_logic_vector(to_unsigned(166,8) ,
24583	 => std_logic_vector(to_unsigned(163,8) ,
24584	 => std_logic_vector(to_unsigned(164,8) ,
24585	 => std_logic_vector(to_unsigned(170,8) ,
24586	 => std_logic_vector(to_unsigned(168,8) ,
24587	 => std_logic_vector(to_unsigned(164,8) ,
24588	 => std_logic_vector(to_unsigned(164,8) ,
24589	 => std_logic_vector(to_unsigned(163,8) ,
24590	 => std_logic_vector(to_unsigned(157,8) ,
24591	 => std_logic_vector(to_unsigned(157,8) ,
24592	 => std_logic_vector(to_unsigned(157,8) ,
24593	 => std_logic_vector(to_unsigned(163,8) ,
24594	 => std_logic_vector(to_unsigned(164,8) ,
24595	 => std_logic_vector(to_unsigned(64,8) ,
24596	 => std_logic_vector(to_unsigned(12,8) ,
24597	 => std_logic_vector(to_unsigned(9,8) ,
24598	 => std_logic_vector(to_unsigned(2,8) ,
24599	 => std_logic_vector(to_unsigned(5,8) ,
24600	 => std_logic_vector(to_unsigned(9,8) ,
24601	 => std_logic_vector(to_unsigned(21,8) ,
24602	 => std_logic_vector(to_unsigned(21,8) ,
24603	 => std_logic_vector(to_unsigned(6,8) ,
24604	 => std_logic_vector(to_unsigned(12,8) ,
24605	 => std_logic_vector(to_unsigned(25,8) ,
24606	 => std_logic_vector(to_unsigned(4,8) ,
24607	 => std_logic_vector(to_unsigned(29,8) ,
24608	 => std_logic_vector(to_unsigned(131,8) ,
24609	 => std_logic_vector(to_unsigned(10,8) ,
24610	 => std_logic_vector(to_unsigned(5,8) ,
24611	 => std_logic_vector(to_unsigned(24,8) ,
24612	 => std_logic_vector(to_unsigned(111,8) ,
24613	 => std_logic_vector(to_unsigned(142,8) ,
24614	 => std_logic_vector(to_unsigned(109,8) ,
24615	 => std_logic_vector(to_unsigned(111,8) ,
24616	 => std_logic_vector(to_unsigned(115,8) ,
24617	 => std_logic_vector(to_unsigned(114,8) ,
24618	 => std_logic_vector(to_unsigned(114,8) ,
24619	 => std_logic_vector(to_unsigned(97,8) ,
24620	 => std_logic_vector(to_unsigned(97,8) ,
24621	 => std_logic_vector(to_unsigned(99,8) ,
24622	 => std_logic_vector(to_unsigned(87,8) ,
24623	 => std_logic_vector(to_unsigned(91,8) ,
24624	 => std_logic_vector(to_unsigned(100,8) ,
24625	 => std_logic_vector(to_unsigned(101,8) ,
24626	 => std_logic_vector(to_unsigned(105,8) ,
24627	 => std_logic_vector(to_unsigned(115,8) ,
24628	 => std_logic_vector(to_unsigned(114,8) ,
24629	 => std_logic_vector(to_unsigned(114,8) ,
24630	 => std_logic_vector(to_unsigned(108,8) ,
24631	 => std_logic_vector(to_unsigned(130,8) ,
24632	 => std_logic_vector(to_unsigned(168,8) ,
24633	 => std_logic_vector(to_unsigned(170,8) ,
24634	 => std_logic_vector(to_unsigned(149,8) ,
24635	 => std_logic_vector(to_unsigned(131,8) ,
24636	 => std_logic_vector(to_unsigned(133,8) ,
24637	 => std_logic_vector(to_unsigned(114,8) ,
24638	 => std_logic_vector(to_unsigned(105,8) ,
24639	 => std_logic_vector(to_unsigned(114,8) ,
24640	 => std_logic_vector(to_unsigned(114,8) ,
24641	 => std_logic_vector(to_unsigned(157,8) ,
24642	 => std_logic_vector(to_unsigned(161,8) ,
24643	 => std_logic_vector(to_unsigned(161,8) ,
24644	 => std_logic_vector(to_unsigned(156,8) ,
24645	 => std_logic_vector(to_unsigned(159,8) ,
24646	 => std_logic_vector(to_unsigned(156,8) ,
24647	 => std_logic_vector(to_unsigned(91,8) ,
24648	 => std_logic_vector(to_unsigned(77,8) ,
24649	 => std_logic_vector(to_unsigned(99,8) ,
24650	 => std_logic_vector(to_unsigned(99,8) ,
24651	 => std_logic_vector(to_unsigned(51,8) ,
24652	 => std_logic_vector(to_unsigned(18,8) ,
24653	 => std_logic_vector(to_unsigned(10,8) ,
24654	 => std_logic_vector(to_unsigned(3,8) ,
24655	 => std_logic_vector(to_unsigned(1,8) ,
24656	 => std_logic_vector(to_unsigned(1,8) ,
24657	 => std_logic_vector(to_unsigned(10,8) ,
24658	 => std_logic_vector(to_unsigned(71,8) ,
24659	 => std_logic_vector(to_unsigned(22,8) ,
24660	 => std_logic_vector(to_unsigned(26,8) ,
24661	 => std_logic_vector(to_unsigned(101,8) ,
24662	 => std_logic_vector(to_unsigned(2,8) ,
24663	 => std_logic_vector(to_unsigned(2,8) ,
24664	 => std_logic_vector(to_unsigned(105,8) ,
24665	 => std_logic_vector(to_unsigned(192,8) ,
24666	 => std_logic_vector(to_unsigned(118,8) ,
24667	 => std_logic_vector(to_unsigned(15,8) ,
24668	 => std_logic_vector(to_unsigned(0,8) ,
24669	 => std_logic_vector(to_unsigned(1,8) ,
24670	 => std_logic_vector(to_unsigned(5,8) ,
24671	 => std_logic_vector(to_unsigned(7,8) ,
24672	 => std_logic_vector(to_unsigned(12,8) ,
24673	 => std_logic_vector(to_unsigned(5,8) ,
24674	 => std_logic_vector(to_unsigned(1,8) ,
24675	 => std_logic_vector(to_unsigned(1,8) ,
24676	 => std_logic_vector(to_unsigned(3,8) ,
24677	 => std_logic_vector(to_unsigned(2,8) ,
24678	 => std_logic_vector(to_unsigned(2,8) ,
24679	 => std_logic_vector(to_unsigned(2,8) ,
24680	 => std_logic_vector(to_unsigned(2,8) ,
24681	 => std_logic_vector(to_unsigned(66,8) ,
24682	 => std_logic_vector(to_unsigned(154,8) ,
24683	 => std_logic_vector(to_unsigned(105,8) ,
24684	 => std_logic_vector(to_unsigned(88,8) ,
24685	 => std_logic_vector(to_unsigned(71,8) ,
24686	 => std_logic_vector(to_unsigned(41,8) ,
24687	 => std_logic_vector(to_unsigned(10,8) ,
24688	 => std_logic_vector(to_unsigned(1,8) ,
24689	 => std_logic_vector(to_unsigned(0,8) ,
24690	 => std_logic_vector(to_unsigned(61,8) ,
24691	 => std_logic_vector(to_unsigned(188,8) ,
24692	 => std_logic_vector(to_unsigned(163,8) ,
24693	 => std_logic_vector(to_unsigned(161,8) ,
24694	 => std_logic_vector(to_unsigned(154,8) ,
24695	 => std_logic_vector(to_unsigned(163,8) ,
24696	 => std_logic_vector(to_unsigned(142,8) ,
24697	 => std_logic_vector(to_unsigned(27,8) ,
24698	 => std_logic_vector(to_unsigned(7,8) ,
24699	 => std_logic_vector(to_unsigned(8,8) ,
24700	 => std_logic_vector(to_unsigned(4,8) ,
24701	 => std_logic_vector(to_unsigned(1,8) ,
24702	 => std_logic_vector(to_unsigned(2,8) ,
24703	 => std_logic_vector(to_unsigned(5,8) ,
24704	 => std_logic_vector(to_unsigned(4,8) ,
24705	 => std_logic_vector(to_unsigned(4,8) ,
24706	 => std_logic_vector(to_unsigned(4,8) ,
24707	 => std_logic_vector(to_unsigned(3,8) ,
24708	 => std_logic_vector(to_unsigned(3,8) ,
24709	 => std_logic_vector(to_unsigned(3,8) ,
24710	 => std_logic_vector(to_unsigned(3,8) ,
24711	 => std_logic_vector(to_unsigned(6,8) ,
24712	 => std_logic_vector(to_unsigned(9,8) ,
24713	 => std_logic_vector(to_unsigned(3,8) ,
24714	 => std_logic_vector(to_unsigned(5,8) ,
24715	 => std_logic_vector(to_unsigned(53,8) ,
24716	 => std_logic_vector(to_unsigned(60,8) ,
24717	 => std_logic_vector(to_unsigned(51,8) ,
24718	 => std_logic_vector(to_unsigned(144,8) ,
24719	 => std_logic_vector(to_unsigned(177,8) ,
24720	 => std_logic_vector(to_unsigned(184,8) ,
24721	 => std_logic_vector(to_unsigned(175,8) ,
24722	 => std_logic_vector(to_unsigned(29,8) ,
24723	 => std_logic_vector(to_unsigned(13,8) ,
24724	 => std_logic_vector(to_unsigned(46,8) ,
24725	 => std_logic_vector(to_unsigned(36,8) ,
24726	 => std_logic_vector(to_unsigned(20,8) ,
24727	 => std_logic_vector(to_unsigned(23,8) ,
24728	 => std_logic_vector(to_unsigned(97,8) ,
24729	 => std_logic_vector(to_unsigned(130,8) ,
24730	 => std_logic_vector(to_unsigned(133,8) ,
24731	 => std_logic_vector(to_unsigned(142,8) ,
24732	 => std_logic_vector(to_unsigned(152,8) ,
24733	 => std_logic_vector(to_unsigned(161,8) ,
24734	 => std_logic_vector(to_unsigned(163,8) ,
24735	 => std_logic_vector(to_unsigned(159,8) ,
24736	 => std_logic_vector(to_unsigned(163,8) ,
24737	 => std_logic_vector(to_unsigned(159,8) ,
24738	 => std_logic_vector(to_unsigned(163,8) ,
24739	 => std_logic_vector(to_unsigned(163,8) ,
24740	 => std_logic_vector(to_unsigned(161,8) ,
24741	 => std_logic_vector(to_unsigned(173,8) ,
24742	 => std_logic_vector(to_unsigned(82,8) ,
24743	 => std_logic_vector(to_unsigned(82,8) ,
24744	 => std_logic_vector(to_unsigned(136,8) ,
24745	 => std_logic_vector(to_unsigned(91,8) ,
24746	 => std_logic_vector(to_unsigned(104,8) ,
24747	 => std_logic_vector(to_unsigned(144,8) ,
24748	 => std_logic_vector(to_unsigned(161,8) ,
24749	 => std_logic_vector(to_unsigned(116,8) ,
24750	 => std_logic_vector(to_unsigned(74,8) ,
24751	 => std_logic_vector(to_unsigned(104,8) ,
24752	 => std_logic_vector(to_unsigned(133,8) ,
24753	 => std_logic_vector(to_unsigned(99,8) ,
24754	 => std_logic_vector(to_unsigned(13,8) ,
24755	 => std_logic_vector(to_unsigned(0,8) ,
24756	 => std_logic_vector(to_unsigned(26,8) ,
24757	 => std_logic_vector(to_unsigned(23,8) ,
24758	 => std_logic_vector(to_unsigned(0,8) ,
24759	 => std_logic_vector(to_unsigned(1,8) ,
24760	 => std_logic_vector(to_unsigned(3,8) ,
24761	 => std_logic_vector(to_unsigned(5,8) ,
24762	 => std_logic_vector(to_unsigned(10,8) ,
24763	 => std_logic_vector(to_unsigned(3,8) ,
24764	 => std_logic_vector(to_unsigned(3,8) ,
24765	 => std_logic_vector(to_unsigned(14,8) ,
24766	 => std_logic_vector(to_unsigned(15,8) ,
24767	 => std_logic_vector(to_unsigned(8,8) ,
24768	 => std_logic_vector(to_unsigned(6,8) ,
24769	 => std_logic_vector(to_unsigned(5,8) ,
24770	 => std_logic_vector(to_unsigned(27,8) ,
24771	 => std_logic_vector(to_unsigned(92,8) ,
24772	 => std_logic_vector(to_unsigned(109,8) ,
24773	 => std_logic_vector(to_unsigned(131,8) ,
24774	 => std_logic_vector(to_unsigned(152,8) ,
24775	 => std_logic_vector(to_unsigned(161,8) ,
24776	 => std_logic_vector(to_unsigned(154,8) ,
24777	 => std_logic_vector(to_unsigned(152,8) ,
24778	 => std_logic_vector(to_unsigned(147,8) ,
24779	 => std_logic_vector(to_unsigned(136,8) ,
24780	 => std_logic_vector(to_unsigned(81,8) ,
24781	 => std_logic_vector(to_unsigned(44,8) ,
24782	 => std_logic_vector(to_unsigned(33,8) ,
24783	 => std_logic_vector(to_unsigned(10,8) ,
24784	 => std_logic_vector(to_unsigned(6,8) ,
24785	 => std_logic_vector(to_unsigned(1,8) ,
24786	 => std_logic_vector(to_unsigned(7,8) ,
24787	 => std_logic_vector(to_unsigned(17,8) ,
24788	 => std_logic_vector(to_unsigned(9,8) ,
24789	 => std_logic_vector(to_unsigned(6,8) ,
24790	 => std_logic_vector(to_unsigned(10,8) ,
24791	 => std_logic_vector(to_unsigned(7,8) ,
24792	 => std_logic_vector(to_unsigned(15,8) ,
24793	 => std_logic_vector(to_unsigned(41,8) ,
24794	 => std_logic_vector(to_unsigned(16,8) ,
24795	 => std_logic_vector(to_unsigned(22,8) ,
24796	 => std_logic_vector(to_unsigned(37,8) ,
24797	 => std_logic_vector(to_unsigned(49,8) ,
24798	 => std_logic_vector(to_unsigned(69,8) ,
24799	 => std_logic_vector(to_unsigned(85,8) ,
24800	 => std_logic_vector(to_unsigned(101,8) ,
24801	 => std_logic_vector(to_unsigned(125,8) ,
24802	 => std_logic_vector(to_unsigned(142,8) ,
24803	 => std_logic_vector(to_unsigned(27,8) ,
24804	 => std_logic_vector(to_unsigned(7,8) ,
24805	 => std_logic_vector(to_unsigned(16,8) ,
24806	 => std_logic_vector(to_unsigned(19,8) ,
24807	 => std_logic_vector(to_unsigned(22,8) ,
24808	 => std_logic_vector(to_unsigned(12,8) ,
24809	 => std_logic_vector(to_unsigned(8,8) ,
24810	 => std_logic_vector(to_unsigned(8,8) ,
24811	 => std_logic_vector(to_unsigned(10,8) ,
24812	 => std_logic_vector(to_unsigned(11,8) ,
24813	 => std_logic_vector(to_unsigned(17,8) ,
24814	 => std_logic_vector(to_unsigned(9,8) ,
24815	 => std_logic_vector(to_unsigned(33,8) ,
24816	 => std_logic_vector(to_unsigned(38,8) ,
24817	 => std_logic_vector(to_unsigned(39,8) ,
24818	 => std_logic_vector(to_unsigned(32,8) ,
24819	 => std_logic_vector(to_unsigned(29,8) ,
24820	 => std_logic_vector(to_unsigned(26,8) ,
24821	 => std_logic_vector(to_unsigned(16,8) ,
24822	 => std_logic_vector(to_unsigned(10,8) ,
24823	 => std_logic_vector(to_unsigned(9,8) ,
24824	 => std_logic_vector(to_unsigned(10,8) ,
24825	 => std_logic_vector(to_unsigned(14,8) ,
24826	 => std_logic_vector(to_unsigned(14,8) ,
24827	 => std_logic_vector(to_unsigned(19,8) ,
24828	 => std_logic_vector(to_unsigned(36,8) ,
24829	 => std_logic_vector(to_unsigned(104,8) ,
24830	 => std_logic_vector(to_unsigned(127,8) ,
24831	 => std_logic_vector(to_unsigned(125,8) ,
24832	 => std_logic_vector(to_unsigned(125,8) ,
24833	 => std_logic_vector(to_unsigned(99,8) ,
24834	 => std_logic_vector(to_unsigned(62,8) ,
24835	 => std_logic_vector(to_unsigned(25,8) ,
24836	 => std_logic_vector(to_unsigned(8,8) ,
24837	 => std_logic_vector(to_unsigned(8,8) ,
24838	 => std_logic_vector(to_unsigned(17,8) ,
24839	 => std_logic_vector(to_unsigned(12,8) ,
24840	 => std_logic_vector(to_unsigned(6,8) ,
24841	 => std_logic_vector(to_unsigned(7,8) ,
24842	 => std_logic_vector(to_unsigned(18,8) ,
24843	 => std_logic_vector(to_unsigned(38,8) ,
24844	 => std_logic_vector(to_unsigned(26,8) ,
24845	 => std_logic_vector(to_unsigned(71,8) ,
24846	 => std_logic_vector(to_unsigned(149,8) ,
24847	 => std_logic_vector(to_unsigned(156,8) ,
24848	 => std_logic_vector(to_unsigned(159,8) ,
24849	 => std_logic_vector(to_unsigned(156,8) ,
24850	 => std_logic_vector(to_unsigned(147,8) ,
24851	 => std_logic_vector(to_unsigned(139,8) ,
24852	 => std_logic_vector(to_unsigned(138,8) ,
24853	 => std_logic_vector(to_unsigned(138,8) ,
24854	 => std_logic_vector(to_unsigned(136,8) ,
24855	 => std_logic_vector(to_unsigned(138,8) ,
24856	 => std_logic_vector(to_unsigned(138,8) ,
24857	 => std_logic_vector(to_unsigned(138,8) ,
24858	 => std_logic_vector(to_unsigned(138,8) ,
24859	 => std_logic_vector(to_unsigned(133,8) ,
24860	 => std_logic_vector(to_unsigned(136,8) ,
24861	 => std_logic_vector(to_unsigned(125,8) ,
24862	 => std_logic_vector(to_unsigned(72,8) ,
24863	 => std_logic_vector(to_unsigned(32,8) ,
24864	 => std_logic_vector(to_unsigned(8,8) ,
24865	 => std_logic_vector(to_unsigned(2,8) ,
24866	 => std_logic_vector(to_unsigned(4,8) ,
24867	 => std_logic_vector(to_unsigned(6,8) ,
24868	 => std_logic_vector(to_unsigned(6,8) ,
24869	 => std_logic_vector(to_unsigned(4,8) ,
24870	 => std_logic_vector(to_unsigned(6,8) ,
24871	 => std_logic_vector(to_unsigned(5,8) ,
24872	 => std_logic_vector(to_unsigned(3,8) ,
24873	 => std_logic_vector(to_unsigned(9,8) ,
24874	 => std_logic_vector(to_unsigned(73,8) ,
24875	 => std_logic_vector(to_unsigned(163,8) ,
24876	 => std_logic_vector(to_unsigned(159,8) ,
24877	 => std_logic_vector(to_unsigned(152,8) ,
24878	 => std_logic_vector(to_unsigned(144,8) ,
24879	 => std_logic_vector(to_unsigned(142,8) ,
24880	 => std_logic_vector(to_unsigned(144,8) ,
24881	 => std_logic_vector(to_unsigned(133,8) ,
24882	 => std_logic_vector(to_unsigned(131,8) ,
24883	 => std_logic_vector(to_unsigned(142,8) ,
24884	 => std_logic_vector(to_unsigned(79,8) ,
24885	 => std_logic_vector(to_unsigned(56,8) ,
24886	 => std_logic_vector(to_unsigned(51,8) ,
24887	 => std_logic_vector(to_unsigned(22,8) ,
24888	 => std_logic_vector(to_unsigned(5,8) ,
24889	 => std_logic_vector(to_unsigned(4,8) ,
24890	 => std_logic_vector(to_unsigned(9,8) ,
24891	 => std_logic_vector(to_unsigned(11,8) ,
24892	 => std_logic_vector(to_unsigned(6,8) ,
24893	 => std_logic_vector(to_unsigned(9,8) ,
24894	 => std_logic_vector(to_unsigned(4,8) ,
24895	 => std_logic_vector(to_unsigned(7,8) ,
24896	 => std_logic_vector(to_unsigned(6,8) ,
24897	 => std_logic_vector(to_unsigned(4,8) ,
24898	 => std_logic_vector(to_unsigned(19,8) ,
24899	 => std_logic_vector(to_unsigned(141,8) ,
24900	 => std_logic_vector(to_unsigned(177,8) ,
24901	 => std_logic_vector(to_unsigned(163,8) ,
24902	 => std_logic_vector(to_unsigned(159,8) ,
24903	 => std_logic_vector(to_unsigned(161,8) ,
24904	 => std_logic_vector(to_unsigned(168,8) ,
24905	 => std_logic_vector(to_unsigned(164,8) ,
24906	 => std_logic_vector(to_unsigned(168,8) ,
24907	 => std_logic_vector(to_unsigned(164,8) ,
24908	 => std_logic_vector(to_unsigned(166,8) ,
24909	 => std_logic_vector(to_unsigned(157,8) ,
24910	 => std_logic_vector(to_unsigned(161,8) ,
24911	 => std_logic_vector(to_unsigned(163,8) ,
24912	 => std_logic_vector(to_unsigned(157,8) ,
24913	 => std_logic_vector(to_unsigned(163,8) ,
24914	 => std_logic_vector(to_unsigned(74,8) ,
24915	 => std_logic_vector(to_unsigned(3,8) ,
24916	 => std_logic_vector(to_unsigned(18,8) ,
24917	 => std_logic_vector(to_unsigned(10,8) ,
24918	 => std_logic_vector(to_unsigned(1,8) ,
24919	 => std_logic_vector(to_unsigned(6,8) ,
24920	 => std_logic_vector(to_unsigned(5,8) ,
24921	 => std_logic_vector(to_unsigned(5,8) ,
24922	 => std_logic_vector(to_unsigned(6,8) ,
24923	 => std_logic_vector(to_unsigned(11,8) ,
24924	 => std_logic_vector(to_unsigned(24,8) ,
24925	 => std_logic_vector(to_unsigned(25,8) ,
24926	 => std_logic_vector(to_unsigned(3,8) ,
24927	 => std_logic_vector(to_unsigned(33,8) ,
24928	 => std_logic_vector(to_unsigned(138,8) ,
24929	 => std_logic_vector(to_unsigned(25,8) ,
24930	 => std_logic_vector(to_unsigned(2,8) ,
24931	 => std_logic_vector(to_unsigned(13,8) ,
24932	 => std_logic_vector(to_unsigned(142,8) ,
24933	 => std_logic_vector(to_unsigned(168,8) ,
24934	 => std_logic_vector(to_unsigned(142,8) ,
24935	 => std_logic_vector(to_unsigned(121,8) ,
24936	 => std_logic_vector(to_unsigned(127,8) ,
24937	 => std_logic_vector(to_unsigned(133,8) ,
24938	 => std_logic_vector(to_unsigned(119,8) ,
24939	 => std_logic_vector(to_unsigned(104,8) ,
24940	 => std_logic_vector(to_unsigned(92,8) ,
24941	 => std_logic_vector(to_unsigned(92,8) ,
24942	 => std_logic_vector(to_unsigned(88,8) ,
24943	 => std_logic_vector(to_unsigned(84,8) ,
24944	 => std_logic_vector(to_unsigned(90,8) ,
24945	 => std_logic_vector(to_unsigned(92,8) ,
24946	 => std_logic_vector(to_unsigned(100,8) ,
24947	 => std_logic_vector(to_unsigned(109,8) ,
24948	 => std_logic_vector(to_unsigned(114,8) ,
24949	 => std_logic_vector(to_unsigned(115,8) ,
24950	 => std_logic_vector(to_unsigned(111,8) ,
24951	 => std_logic_vector(to_unsigned(116,8) ,
24952	 => std_logic_vector(to_unsigned(154,8) ,
24953	 => std_logic_vector(to_unsigned(170,8) ,
24954	 => std_logic_vector(to_unsigned(168,8) ,
24955	 => std_logic_vector(to_unsigned(147,8) ,
24956	 => std_logic_vector(to_unsigned(122,8) ,
24957	 => std_logic_vector(to_unsigned(121,8) ,
24958	 => std_logic_vector(to_unsigned(115,8) ,
24959	 => std_logic_vector(to_unsigned(115,8) ,
24960	 => std_logic_vector(to_unsigned(111,8) ,
24961	 => std_logic_vector(to_unsigned(163,8) ,
24962	 => std_logic_vector(to_unsigned(163,8) ,
24963	 => std_logic_vector(to_unsigned(163,8) ,
24964	 => std_logic_vector(to_unsigned(154,8) ,
24965	 => std_logic_vector(to_unsigned(159,8) ,
24966	 => std_logic_vector(to_unsigned(154,8) ,
24967	 => std_logic_vector(to_unsigned(101,8) ,
24968	 => std_logic_vector(to_unsigned(99,8) ,
24969	 => std_logic_vector(to_unsigned(90,8) ,
24970	 => std_logic_vector(to_unsigned(85,8) ,
24971	 => std_logic_vector(to_unsigned(74,8) ,
24972	 => std_logic_vector(to_unsigned(45,8) ,
24973	 => std_logic_vector(to_unsigned(13,8) ,
24974	 => std_logic_vector(to_unsigned(2,8) ,
24975	 => std_logic_vector(to_unsigned(0,8) ,
24976	 => std_logic_vector(to_unsigned(4,8) ,
24977	 => std_logic_vector(to_unsigned(13,8) ,
24978	 => std_logic_vector(to_unsigned(12,8) ,
24979	 => std_logic_vector(to_unsigned(1,8) ,
24980	 => std_logic_vector(to_unsigned(15,8) ,
24981	 => std_logic_vector(to_unsigned(151,8) ,
24982	 => std_logic_vector(to_unsigned(67,8) ,
24983	 => std_logic_vector(to_unsigned(52,8) ,
24984	 => std_logic_vector(to_unsigned(147,8) ,
24985	 => std_logic_vector(to_unsigned(151,8) ,
24986	 => std_logic_vector(to_unsigned(152,8) ,
24987	 => std_logic_vector(to_unsigned(86,8) ,
24988	 => std_logic_vector(to_unsigned(7,8) ,
24989	 => std_logic_vector(to_unsigned(0,8) ,
24990	 => std_logic_vector(to_unsigned(3,8) ,
24991	 => std_logic_vector(to_unsigned(8,8) ,
24992	 => std_logic_vector(to_unsigned(7,8) ,
24993	 => std_logic_vector(to_unsigned(6,8) ,
24994	 => std_logic_vector(to_unsigned(2,8) ,
24995	 => std_logic_vector(to_unsigned(1,8) ,
24996	 => std_logic_vector(to_unsigned(1,8) ,
24997	 => std_logic_vector(to_unsigned(1,8) ,
24998	 => std_logic_vector(to_unsigned(3,8) ,
24999	 => std_logic_vector(to_unsigned(2,8) ,
25000	 => std_logic_vector(to_unsigned(6,8) ,
25001	 => std_logic_vector(to_unsigned(133,8) ,
25002	 => std_logic_vector(to_unsigned(168,8) ,
25003	 => std_logic_vector(to_unsigned(141,8) ,
25004	 => std_logic_vector(to_unsigned(122,8) ,
25005	 => std_logic_vector(to_unsigned(93,8) ,
25006	 => std_logic_vector(to_unsigned(39,8) ,
25007	 => std_logic_vector(to_unsigned(5,8) ,
25008	 => std_logic_vector(to_unsigned(0,8) ,
25009	 => std_logic_vector(to_unsigned(1,8) ,
25010	 => std_logic_vector(to_unsigned(92,8) ,
25011	 => std_logic_vector(to_unsigned(188,8) ,
25012	 => std_logic_vector(to_unsigned(157,8) ,
25013	 => std_logic_vector(to_unsigned(156,8) ,
25014	 => std_logic_vector(to_unsigned(154,8) ,
25015	 => std_logic_vector(to_unsigned(146,8) ,
25016	 => std_logic_vector(to_unsigned(111,8) ,
25017	 => std_logic_vector(to_unsigned(26,8) ,
25018	 => std_logic_vector(to_unsigned(9,8) ,
25019	 => std_logic_vector(to_unsigned(8,8) ,
25020	 => std_logic_vector(to_unsigned(4,8) ,
25021	 => std_logic_vector(to_unsigned(8,8) ,
25022	 => std_logic_vector(to_unsigned(3,8) ,
25023	 => std_logic_vector(to_unsigned(3,8) ,
25024	 => std_logic_vector(to_unsigned(5,8) ,
25025	 => std_logic_vector(to_unsigned(4,8) ,
25026	 => std_logic_vector(to_unsigned(4,8) ,
25027	 => std_logic_vector(to_unsigned(3,8) ,
25028	 => std_logic_vector(to_unsigned(3,8) ,
25029	 => std_logic_vector(to_unsigned(3,8) ,
25030	 => std_logic_vector(to_unsigned(4,8) ,
25031	 => std_logic_vector(to_unsigned(6,8) ,
25032	 => std_logic_vector(to_unsigned(7,8) ,
25033	 => std_logic_vector(to_unsigned(5,8) ,
25034	 => std_logic_vector(to_unsigned(1,8) ,
25035	 => std_logic_vector(to_unsigned(28,8) ,
25036	 => std_logic_vector(to_unsigned(82,8) ,
25037	 => std_logic_vector(to_unsigned(46,8) ,
25038	 => std_logic_vector(to_unsigned(69,8) ,
25039	 => std_logic_vector(to_unsigned(156,8) ,
25040	 => std_logic_vector(to_unsigned(161,8) ,
25041	 => std_logic_vector(to_unsigned(170,8) ,
25042	 => std_logic_vector(to_unsigned(30,8) ,
25043	 => std_logic_vector(to_unsigned(13,8) ,
25044	 => std_logic_vector(to_unsigned(44,8) ,
25045	 => std_logic_vector(to_unsigned(23,8) ,
25046	 => std_logic_vector(to_unsigned(12,8) ,
25047	 => std_logic_vector(to_unsigned(41,8) ,
25048	 => std_logic_vector(to_unsigned(116,8) ,
25049	 => std_logic_vector(to_unsigned(138,8) ,
25050	 => std_logic_vector(to_unsigned(138,8) ,
25051	 => std_logic_vector(to_unsigned(134,8) ,
25052	 => std_logic_vector(to_unsigned(157,8) ,
25053	 => std_logic_vector(to_unsigned(161,8) ,
25054	 => std_logic_vector(to_unsigned(157,8) ,
25055	 => std_logic_vector(to_unsigned(138,8) ,
25056	 => std_logic_vector(to_unsigned(147,8) ,
25057	 => std_logic_vector(to_unsigned(164,8) ,
25058	 => std_logic_vector(to_unsigned(157,8) ,
25059	 => std_logic_vector(to_unsigned(161,8) ,
25060	 => std_logic_vector(to_unsigned(163,8) ,
25061	 => std_logic_vector(to_unsigned(159,8) ,
25062	 => std_logic_vector(to_unsigned(57,8) ,
25063	 => std_logic_vector(to_unsigned(72,8) ,
25064	 => std_logic_vector(to_unsigned(128,8) ,
25065	 => std_logic_vector(to_unsigned(74,8) ,
25066	 => std_logic_vector(to_unsigned(97,8) ,
25067	 => std_logic_vector(to_unsigned(133,8) ,
25068	 => std_logic_vector(to_unsigned(154,8) ,
25069	 => std_logic_vector(to_unsigned(108,8) ,
25070	 => std_logic_vector(to_unsigned(88,8) ,
25071	 => std_logic_vector(to_unsigned(121,8) ,
25072	 => std_logic_vector(to_unsigned(112,8) ,
25073	 => std_logic_vector(to_unsigned(90,8) ,
25074	 => std_logic_vector(to_unsigned(12,8) ,
25075	 => std_logic_vector(to_unsigned(2,8) ,
25076	 => std_logic_vector(to_unsigned(73,8) ,
25077	 => std_logic_vector(to_unsigned(24,8) ,
25078	 => std_logic_vector(to_unsigned(1,8) ,
25079	 => std_logic_vector(to_unsigned(0,8) ,
25080	 => std_logic_vector(to_unsigned(2,8) ,
25081	 => std_logic_vector(to_unsigned(3,8) ,
25082	 => std_logic_vector(to_unsigned(2,8) ,
25083	 => std_logic_vector(to_unsigned(4,8) ,
25084	 => std_logic_vector(to_unsigned(4,8) ,
25085	 => std_logic_vector(to_unsigned(4,8) ,
25086	 => std_logic_vector(to_unsigned(12,8) ,
25087	 => std_logic_vector(to_unsigned(11,8) ,
25088	 => std_logic_vector(to_unsigned(4,8) ,
25089	 => std_logic_vector(to_unsigned(6,8) ,
25090	 => std_logic_vector(to_unsigned(38,8) ,
25091	 => std_logic_vector(to_unsigned(74,8) ,
25092	 => std_logic_vector(to_unsigned(124,8) ,
25093	 => std_logic_vector(to_unsigned(136,8) ,
25094	 => std_logic_vector(to_unsigned(139,8) ,
25095	 => std_logic_vector(to_unsigned(159,8) ,
25096	 => std_logic_vector(to_unsigned(157,8) ,
25097	 => std_logic_vector(to_unsigned(157,8) ,
25098	 => std_logic_vector(to_unsigned(144,8) ,
25099	 => std_logic_vector(to_unsigned(92,8) ,
25100	 => std_logic_vector(to_unsigned(38,8) ,
25101	 => std_logic_vector(to_unsigned(35,8) ,
25102	 => std_logic_vector(to_unsigned(25,8) ,
25103	 => std_logic_vector(to_unsigned(23,8) ,
25104	 => std_logic_vector(to_unsigned(18,8) ,
25105	 => std_logic_vector(to_unsigned(2,8) ,
25106	 => std_logic_vector(to_unsigned(3,8) ,
25107	 => std_logic_vector(to_unsigned(12,8) ,
25108	 => std_logic_vector(to_unsigned(6,8) ,
25109	 => std_logic_vector(to_unsigned(8,8) ,
25110	 => std_logic_vector(to_unsigned(17,8) ,
25111	 => std_logic_vector(to_unsigned(7,8) ,
25112	 => std_logic_vector(to_unsigned(28,8) ,
25113	 => std_logic_vector(to_unsigned(51,8) ,
25114	 => std_logic_vector(to_unsigned(21,8) ,
25115	 => std_logic_vector(to_unsigned(27,8) ,
25116	 => std_logic_vector(to_unsigned(49,8) ,
25117	 => std_logic_vector(to_unsigned(48,8) ,
25118	 => std_logic_vector(to_unsigned(44,8) ,
25119	 => std_logic_vector(to_unsigned(39,8) ,
25120	 => std_logic_vector(to_unsigned(36,8) ,
25121	 => std_logic_vector(to_unsigned(56,8) ,
25122	 => std_logic_vector(to_unsigned(111,8) ,
25123	 => std_logic_vector(to_unsigned(24,8) ,
25124	 => std_logic_vector(to_unsigned(13,8) ,
25125	 => std_logic_vector(to_unsigned(27,8) ,
25126	 => std_logic_vector(to_unsigned(24,8) ,
25127	 => std_logic_vector(to_unsigned(29,8) ,
25128	 => std_logic_vector(to_unsigned(19,8) ,
25129	 => std_logic_vector(to_unsigned(13,8) ,
25130	 => std_logic_vector(to_unsigned(9,8) ,
25131	 => std_logic_vector(to_unsigned(12,8) ,
25132	 => std_logic_vector(to_unsigned(14,8) ,
25133	 => std_logic_vector(to_unsigned(27,8) ,
25134	 => std_logic_vector(to_unsigned(18,8) ,
25135	 => std_logic_vector(to_unsigned(27,8) ,
25136	 => std_logic_vector(to_unsigned(39,8) ,
25137	 => std_logic_vector(to_unsigned(29,8) ,
25138	 => std_logic_vector(to_unsigned(26,8) ,
25139	 => std_logic_vector(to_unsigned(26,8) ,
25140	 => std_logic_vector(to_unsigned(25,8) ,
25141	 => std_logic_vector(to_unsigned(19,8) ,
25142	 => std_logic_vector(to_unsigned(13,8) ,
25143	 => std_logic_vector(to_unsigned(11,8) ,
25144	 => std_logic_vector(to_unsigned(8,8) ,
25145	 => std_logic_vector(to_unsigned(10,8) ,
25146	 => std_logic_vector(to_unsigned(14,8) ,
25147	 => std_logic_vector(to_unsigned(15,8) ,
25148	 => std_logic_vector(to_unsigned(26,8) ,
25149	 => std_logic_vector(to_unsigned(104,8) ,
25150	 => std_logic_vector(to_unsigned(149,8) ,
25151	 => std_logic_vector(to_unsigned(128,8) ,
25152	 => std_logic_vector(to_unsigned(116,8) ,
25153	 => std_logic_vector(to_unsigned(51,8) ,
25154	 => std_logic_vector(to_unsigned(62,8) ,
25155	 => std_logic_vector(to_unsigned(44,8) ,
25156	 => std_logic_vector(to_unsigned(7,8) ,
25157	 => std_logic_vector(to_unsigned(7,8) ,
25158	 => std_logic_vector(to_unsigned(13,8) ,
25159	 => std_logic_vector(to_unsigned(42,8) ,
25160	 => std_logic_vector(to_unsigned(44,8) ,
25161	 => std_logic_vector(to_unsigned(19,8) ,
25162	 => std_logic_vector(to_unsigned(24,8) ,
25163	 => std_logic_vector(to_unsigned(45,8) ,
25164	 => std_logic_vector(to_unsigned(13,8) ,
25165	 => std_logic_vector(to_unsigned(48,8) ,
25166	 => std_logic_vector(to_unsigned(163,8) ,
25167	 => std_logic_vector(to_unsigned(152,8) ,
25168	 => std_logic_vector(to_unsigned(156,8) ,
25169	 => std_logic_vector(to_unsigned(157,8) ,
25170	 => std_logic_vector(to_unsigned(159,8) ,
25171	 => std_logic_vector(to_unsigned(154,8) ,
25172	 => std_logic_vector(to_unsigned(138,8) ,
25173	 => std_logic_vector(to_unsigned(134,8) ,
25174	 => std_logic_vector(to_unsigned(138,8) ,
25175	 => std_logic_vector(to_unsigned(136,8) ,
25176	 => std_logic_vector(to_unsigned(136,8) ,
25177	 => std_logic_vector(to_unsigned(136,8) ,
25178	 => std_logic_vector(to_unsigned(133,8) ,
25179	 => std_logic_vector(to_unsigned(133,8) ,
25180	 => std_logic_vector(to_unsigned(138,8) ,
25181	 => std_logic_vector(to_unsigned(72,8) ,
25182	 => std_logic_vector(to_unsigned(20,8) ,
25183	 => std_logic_vector(to_unsigned(14,8) ,
25184	 => std_logic_vector(to_unsigned(13,8) ,
25185	 => std_logic_vector(to_unsigned(6,8) ,
25186	 => std_logic_vector(to_unsigned(6,8) ,
25187	 => std_logic_vector(to_unsigned(9,8) ,
25188	 => std_logic_vector(to_unsigned(8,8) ,
25189	 => std_logic_vector(to_unsigned(4,8) ,
25190	 => std_logic_vector(to_unsigned(4,8) ,
25191	 => std_logic_vector(to_unsigned(3,8) ,
25192	 => std_logic_vector(to_unsigned(6,8) ,
25193	 => std_logic_vector(to_unsigned(10,8) ,
25194	 => std_logic_vector(to_unsigned(20,8) ,
25195	 => std_logic_vector(to_unsigned(67,8) ,
25196	 => std_logic_vector(to_unsigned(138,8) ,
25197	 => std_logic_vector(to_unsigned(161,8) ,
25198	 => std_logic_vector(to_unsigned(156,8) ,
25199	 => std_logic_vector(to_unsigned(151,8) ,
25200	 => std_logic_vector(to_unsigned(142,8) ,
25201	 => std_logic_vector(to_unsigned(136,8) ,
25202	 => std_logic_vector(to_unsigned(154,8) ,
25203	 => std_logic_vector(to_unsigned(108,8) ,
25204	 => std_logic_vector(to_unsigned(4,8) ,
25205	 => std_logic_vector(to_unsigned(0,8) ,
25206	 => std_logic_vector(to_unsigned(1,8) ,
25207	 => std_logic_vector(to_unsigned(1,8) ,
25208	 => std_logic_vector(to_unsigned(5,8) ,
25209	 => std_logic_vector(to_unsigned(17,8) ,
25210	 => std_logic_vector(to_unsigned(16,8) ,
25211	 => std_logic_vector(to_unsigned(13,8) ,
25212	 => std_logic_vector(to_unsigned(10,8) ,
25213	 => std_logic_vector(to_unsigned(15,8) ,
25214	 => std_logic_vector(to_unsigned(19,8) ,
25215	 => std_logic_vector(to_unsigned(8,8) ,
25216	 => std_logic_vector(to_unsigned(7,8) ,
25217	 => std_logic_vector(to_unsigned(6,8) ,
25218	 => std_logic_vector(to_unsigned(16,8) ,
25219	 => std_logic_vector(to_unsigned(108,8) ,
25220	 => std_logic_vector(to_unsigned(171,8) ,
25221	 => std_logic_vector(to_unsigned(177,8) ,
25222	 => std_logic_vector(to_unsigned(183,8) ,
25223	 => std_logic_vector(to_unsigned(170,8) ,
25224	 => std_logic_vector(to_unsigned(164,8) ,
25225	 => std_logic_vector(to_unsigned(164,8) ,
25226	 => std_logic_vector(to_unsigned(163,8) ,
25227	 => std_logic_vector(to_unsigned(170,8) ,
25228	 => std_logic_vector(to_unsigned(168,8) ,
25229	 => std_logic_vector(to_unsigned(161,8) ,
25230	 => std_logic_vector(to_unsigned(166,8) ,
25231	 => std_logic_vector(to_unsigned(166,8) ,
25232	 => std_logic_vector(to_unsigned(133,8) ,
25233	 => std_logic_vector(to_unsigned(91,8) ,
25234	 => std_logic_vector(to_unsigned(30,8) ,
25235	 => std_logic_vector(to_unsigned(20,8) ,
25236	 => std_logic_vector(to_unsigned(62,8) ,
25237	 => std_logic_vector(to_unsigned(12,8) ,
25238	 => std_logic_vector(to_unsigned(1,8) ,
25239	 => std_logic_vector(to_unsigned(5,8) ,
25240	 => std_logic_vector(to_unsigned(6,8) ,
25241	 => std_logic_vector(to_unsigned(8,8) ,
25242	 => std_logic_vector(to_unsigned(14,8) ,
25243	 => std_logic_vector(to_unsigned(18,8) ,
25244	 => std_logic_vector(to_unsigned(19,8) ,
25245	 => std_logic_vector(to_unsigned(20,8) ,
25246	 => std_logic_vector(to_unsigned(4,8) ,
25247	 => std_logic_vector(to_unsigned(56,8) ,
25248	 => std_logic_vector(to_unsigned(133,8) ,
25249	 => std_logic_vector(to_unsigned(23,8) ,
25250	 => std_logic_vector(to_unsigned(7,8) ,
25251	 => std_logic_vector(to_unsigned(52,8) ,
25252	 => std_logic_vector(to_unsigned(121,8) ,
25253	 => std_logic_vector(to_unsigned(133,8) ,
25254	 => std_logic_vector(to_unsigned(161,8) ,
25255	 => std_logic_vector(to_unsigned(154,8) ,
25256	 => std_logic_vector(to_unsigned(141,8) ,
25257	 => std_logic_vector(to_unsigned(128,8) ,
25258	 => std_logic_vector(to_unsigned(116,8) ,
25259	 => std_logic_vector(to_unsigned(109,8) ,
25260	 => std_logic_vector(to_unsigned(100,8) ,
25261	 => std_logic_vector(to_unsigned(97,8) ,
25262	 => std_logic_vector(to_unsigned(95,8) ,
25263	 => std_logic_vector(to_unsigned(90,8) ,
25264	 => std_logic_vector(to_unsigned(93,8) ,
25265	 => std_logic_vector(to_unsigned(97,8) ,
25266	 => std_logic_vector(to_unsigned(103,8) ,
25267	 => std_logic_vector(to_unsigned(108,8) ,
25268	 => std_logic_vector(to_unsigned(105,8) ,
25269	 => std_logic_vector(to_unsigned(112,8) ,
25270	 => std_logic_vector(to_unsigned(127,8) ,
25271	 => std_logic_vector(to_unsigned(118,8) ,
25272	 => std_logic_vector(to_unsigned(134,8) ,
25273	 => std_logic_vector(to_unsigned(164,8) ,
25274	 => std_logic_vector(to_unsigned(168,8) ,
25275	 => std_logic_vector(to_unsigned(163,8) ,
25276	 => std_logic_vector(to_unsigned(139,8) ,
25277	 => std_logic_vector(to_unsigned(125,8) ,
25278	 => std_logic_vector(to_unsigned(125,8) ,
25279	 => std_logic_vector(to_unsigned(115,8) ,
25280	 => std_logic_vector(to_unsigned(109,8) ,
25281	 => std_logic_vector(to_unsigned(161,8) ,
25282	 => std_logic_vector(to_unsigned(163,8) ,
25283	 => std_logic_vector(to_unsigned(161,8) ,
25284	 => std_logic_vector(to_unsigned(157,8) ,
25285	 => std_logic_vector(to_unsigned(163,8) ,
25286	 => std_logic_vector(to_unsigned(156,8) ,
25287	 => std_logic_vector(to_unsigned(90,8) ,
25288	 => std_logic_vector(to_unsigned(56,8) ,
25289	 => std_logic_vector(to_unsigned(43,8) ,
25290	 => std_logic_vector(to_unsigned(34,8) ,
25291	 => std_logic_vector(to_unsigned(23,8) ,
25292	 => std_logic_vector(to_unsigned(19,8) ,
25293	 => std_logic_vector(to_unsigned(12,8) ,
25294	 => std_logic_vector(to_unsigned(4,8) ,
25295	 => std_logic_vector(to_unsigned(12,8) ,
25296	 => std_logic_vector(to_unsigned(54,8) ,
25297	 => std_logic_vector(to_unsigned(60,8) ,
25298	 => std_logic_vector(to_unsigned(14,8) ,
25299	 => std_logic_vector(to_unsigned(1,8) ,
25300	 => std_logic_vector(to_unsigned(1,8) ,
25301	 => std_logic_vector(to_unsigned(72,8) ,
25302	 => std_logic_vector(to_unsigned(171,8) ,
25303	 => std_logic_vector(to_unsigned(154,8) ,
25304	 => std_logic_vector(to_unsigned(136,8) ,
25305	 => std_logic_vector(to_unsigned(121,8) ,
25306	 => std_logic_vector(to_unsigned(114,8) ,
25307	 => std_logic_vector(to_unsigned(146,8) ,
25308	 => std_logic_vector(to_unsigned(121,8) ,
25309	 => std_logic_vector(to_unsigned(27,8) ,
25310	 => std_logic_vector(to_unsigned(2,8) ,
25311	 => std_logic_vector(to_unsigned(2,8) ,
25312	 => std_logic_vector(to_unsigned(4,8) ,
25313	 => std_logic_vector(to_unsigned(6,8) ,
25314	 => std_logic_vector(to_unsigned(2,8) ,
25315	 => std_logic_vector(to_unsigned(1,8) ,
25316	 => std_logic_vector(to_unsigned(2,8) ,
25317	 => std_logic_vector(to_unsigned(2,8) ,
25318	 => std_logic_vector(to_unsigned(3,8) ,
25319	 => std_logic_vector(to_unsigned(2,8) ,
25320	 => std_logic_vector(to_unsigned(11,8) ,
25321	 => std_logic_vector(to_unsigned(141,8) ,
25322	 => std_logic_vector(to_unsigned(152,8) ,
25323	 => std_logic_vector(to_unsigned(146,8) ,
25324	 => std_logic_vector(to_unsigned(133,8) ,
25325	 => std_logic_vector(to_unsigned(82,8) ,
25326	 => std_logic_vector(to_unsigned(33,8) ,
25327	 => std_logic_vector(to_unsigned(3,8) ,
25328	 => std_logic_vector(to_unsigned(0,8) ,
25329	 => std_logic_vector(to_unsigned(1,8) ,
25330	 => std_logic_vector(to_unsigned(108,8) ,
25331	 => std_logic_vector(to_unsigned(186,8) ,
25332	 => std_logic_vector(to_unsigned(157,8) ,
25333	 => std_logic_vector(to_unsigned(151,8) ,
25334	 => std_logic_vector(to_unsigned(149,8) ,
25335	 => std_logic_vector(to_unsigned(152,8) ,
25336	 => std_logic_vector(to_unsigned(96,8) ,
25337	 => std_logic_vector(to_unsigned(17,8) ,
25338	 => std_logic_vector(to_unsigned(10,8) ,
25339	 => std_logic_vector(to_unsigned(13,8) ,
25340	 => std_logic_vector(to_unsigned(5,8) ,
25341	 => std_logic_vector(to_unsigned(6,8) ,
25342	 => std_logic_vector(to_unsigned(9,8) ,
25343	 => std_logic_vector(to_unsigned(4,8) ,
25344	 => std_logic_vector(to_unsigned(4,8) ,
25345	 => std_logic_vector(to_unsigned(5,8) ,
25346	 => std_logic_vector(to_unsigned(4,8) ,
25347	 => std_logic_vector(to_unsigned(4,8) ,
25348	 => std_logic_vector(to_unsigned(4,8) ,
25349	 => std_logic_vector(to_unsigned(4,8) ,
25350	 => std_logic_vector(to_unsigned(6,8) ,
25351	 => std_logic_vector(to_unsigned(6,8) ,
25352	 => std_logic_vector(to_unsigned(7,8) ,
25353	 => std_logic_vector(to_unsigned(9,8) ,
25354	 => std_logic_vector(to_unsigned(2,8) ,
25355	 => std_logic_vector(to_unsigned(7,8) ,
25356	 => std_logic_vector(to_unsigned(80,8) ,
25357	 => std_logic_vector(to_unsigned(67,8) ,
25358	 => std_logic_vector(to_unsigned(70,8) ,
25359	 => std_logic_vector(to_unsigned(142,8) ,
25360	 => std_logic_vector(to_unsigned(179,8) ,
25361	 => std_logic_vector(to_unsigned(141,8) ,
25362	 => std_logic_vector(to_unsigned(14,8) ,
25363	 => std_logic_vector(to_unsigned(19,8) ,
25364	 => std_logic_vector(to_unsigned(40,8) ,
25365	 => std_logic_vector(to_unsigned(13,8) ,
25366	 => std_logic_vector(to_unsigned(6,8) ,
25367	 => std_logic_vector(to_unsigned(57,8) ,
25368	 => std_logic_vector(to_unsigned(133,8) ,
25369	 => std_logic_vector(to_unsigned(139,8) ,
25370	 => std_logic_vector(to_unsigned(141,8) ,
25371	 => std_logic_vector(to_unsigned(114,8) ,
25372	 => std_logic_vector(to_unsigned(121,8) ,
25373	 => std_logic_vector(to_unsigned(154,8) ,
25374	 => std_logic_vector(to_unsigned(163,8) ,
25375	 => std_logic_vector(to_unsigned(154,8) ,
25376	 => std_logic_vector(to_unsigned(154,8) ,
25377	 => std_logic_vector(to_unsigned(164,8) ,
25378	 => std_logic_vector(to_unsigned(154,8) ,
25379	 => std_logic_vector(to_unsigned(144,8) ,
25380	 => std_logic_vector(to_unsigned(151,8) ,
25381	 => std_logic_vector(to_unsigned(147,8) ,
25382	 => std_logic_vector(to_unsigned(25,8) ,
25383	 => std_logic_vector(to_unsigned(44,8) ,
25384	 => std_logic_vector(to_unsigned(107,8) ,
25385	 => std_logic_vector(to_unsigned(88,8) ,
25386	 => std_logic_vector(to_unsigned(108,8) ,
25387	 => std_logic_vector(to_unsigned(125,8) ,
25388	 => std_logic_vector(to_unsigned(152,8) ,
25389	 => std_logic_vector(to_unsigned(115,8) ,
25390	 => std_logic_vector(to_unsigned(72,8) ,
25391	 => std_logic_vector(to_unsigned(95,8) ,
25392	 => std_logic_vector(to_unsigned(81,8) ,
25393	 => std_logic_vector(to_unsigned(88,8) ,
25394	 => std_logic_vector(to_unsigned(11,8) ,
25395	 => std_logic_vector(to_unsigned(7,8) ,
25396	 => std_logic_vector(to_unsigned(69,8) ,
25397	 => std_logic_vector(to_unsigned(18,8) ,
25398	 => std_logic_vector(to_unsigned(7,8) ,
25399	 => std_logic_vector(to_unsigned(1,8) ,
25400	 => std_logic_vector(to_unsigned(1,8) ,
25401	 => std_logic_vector(to_unsigned(2,8) ,
25402	 => std_logic_vector(to_unsigned(1,8) ,
25403	 => std_logic_vector(to_unsigned(5,8) ,
25404	 => std_logic_vector(to_unsigned(7,8) ,
25405	 => std_logic_vector(to_unsigned(5,8) ,
25406	 => std_logic_vector(to_unsigned(17,8) ,
25407	 => std_logic_vector(to_unsigned(11,8) ,
25408	 => std_logic_vector(to_unsigned(2,8) ,
25409	 => std_logic_vector(to_unsigned(6,8) ,
25410	 => std_logic_vector(to_unsigned(32,8) ,
25411	 => std_logic_vector(to_unsigned(81,8) ,
25412	 => std_logic_vector(to_unsigned(144,8) ,
25413	 => std_logic_vector(to_unsigned(147,8) ,
25414	 => std_logic_vector(to_unsigned(139,8) ,
25415	 => std_logic_vector(to_unsigned(154,8) ,
25416	 => std_logic_vector(to_unsigned(154,8) ,
25417	 => std_logic_vector(to_unsigned(161,8) ,
25418	 => std_logic_vector(to_unsigned(124,8) ,
25419	 => std_logic_vector(to_unsigned(53,8) ,
25420	 => std_logic_vector(to_unsigned(22,8) ,
25421	 => std_logic_vector(to_unsigned(7,8) ,
25422	 => std_logic_vector(to_unsigned(4,8) ,
25423	 => std_logic_vector(to_unsigned(9,8) ,
25424	 => std_logic_vector(to_unsigned(18,8) ,
25425	 => std_logic_vector(to_unsigned(11,8) ,
25426	 => std_logic_vector(to_unsigned(6,8) ,
25427	 => std_logic_vector(to_unsigned(9,8) ,
25428	 => std_logic_vector(to_unsigned(10,8) ,
25429	 => std_logic_vector(to_unsigned(13,8) ,
25430	 => std_logic_vector(to_unsigned(14,8) ,
25431	 => std_logic_vector(to_unsigned(7,8) ,
25432	 => std_logic_vector(to_unsigned(24,8) ,
25433	 => std_logic_vector(to_unsigned(57,8) ,
25434	 => std_logic_vector(to_unsigned(33,8) ,
25435	 => std_logic_vector(to_unsigned(32,8) ,
25436	 => std_logic_vector(to_unsigned(51,8) ,
25437	 => std_logic_vector(to_unsigned(37,8) ,
25438	 => std_logic_vector(to_unsigned(33,8) ,
25439	 => std_logic_vector(to_unsigned(33,8) ,
25440	 => std_logic_vector(to_unsigned(38,8) ,
25441	 => std_logic_vector(to_unsigned(41,8) ,
25442	 => std_logic_vector(to_unsigned(61,8) ,
25443	 => std_logic_vector(to_unsigned(25,8) ,
25444	 => std_logic_vector(to_unsigned(16,8) ,
25445	 => std_logic_vector(to_unsigned(33,8) ,
25446	 => std_logic_vector(to_unsigned(30,8) ,
25447	 => std_logic_vector(to_unsigned(30,8) ,
25448	 => std_logic_vector(to_unsigned(25,8) ,
25449	 => std_logic_vector(to_unsigned(22,8) ,
25450	 => std_logic_vector(to_unsigned(13,8) ,
25451	 => std_logic_vector(to_unsigned(12,8) ,
25452	 => std_logic_vector(to_unsigned(17,8) ,
25453	 => std_logic_vector(to_unsigned(17,8) ,
25454	 => std_logic_vector(to_unsigned(13,8) ,
25455	 => std_logic_vector(to_unsigned(17,8) ,
25456	 => std_logic_vector(to_unsigned(25,8) ,
25457	 => std_logic_vector(to_unsigned(25,8) ,
25458	 => std_logic_vector(to_unsigned(29,8) ,
25459	 => std_logic_vector(to_unsigned(27,8) ,
25460	 => std_logic_vector(to_unsigned(23,8) ,
25461	 => std_logic_vector(to_unsigned(17,8) ,
25462	 => std_logic_vector(to_unsigned(13,8) ,
25463	 => std_logic_vector(to_unsigned(10,8) ,
25464	 => std_logic_vector(to_unsigned(8,8) ,
25465	 => std_logic_vector(to_unsigned(9,8) ,
25466	 => std_logic_vector(to_unsigned(12,8) ,
25467	 => std_logic_vector(to_unsigned(9,8) ,
25468	 => std_logic_vector(to_unsigned(48,8) ,
25469	 => std_logic_vector(to_unsigned(127,8) ,
25470	 => std_logic_vector(to_unsigned(125,8) ,
25471	 => std_logic_vector(to_unsigned(124,8) ,
25472	 => std_logic_vector(to_unsigned(103,8) ,
25473	 => std_logic_vector(to_unsigned(30,8) ,
25474	 => std_logic_vector(to_unsigned(67,8) ,
25475	 => std_logic_vector(to_unsigned(55,8) ,
25476	 => std_logic_vector(to_unsigned(2,8) ,
25477	 => std_logic_vector(to_unsigned(5,8) ,
25478	 => std_logic_vector(to_unsigned(9,8) ,
25479	 => std_logic_vector(to_unsigned(17,8) ,
25480	 => std_logic_vector(to_unsigned(14,8) ,
25481	 => std_logic_vector(to_unsigned(8,8) ,
25482	 => std_logic_vector(to_unsigned(27,8) ,
25483	 => std_logic_vector(to_unsigned(42,8) ,
25484	 => std_logic_vector(to_unsigned(11,8) ,
25485	 => std_logic_vector(to_unsigned(71,8) ,
25486	 => std_logic_vector(to_unsigned(173,8) ,
25487	 => std_logic_vector(to_unsigned(147,8) ,
25488	 => std_logic_vector(to_unsigned(154,8) ,
25489	 => std_logic_vector(to_unsigned(154,8) ,
25490	 => std_logic_vector(to_unsigned(157,8) ,
25491	 => std_logic_vector(to_unsigned(161,8) ,
25492	 => std_logic_vector(to_unsigned(147,8) ,
25493	 => std_logic_vector(to_unsigned(136,8) ,
25494	 => std_logic_vector(to_unsigned(141,8) ,
25495	 => std_logic_vector(to_unsigned(142,8) ,
25496	 => std_logic_vector(to_unsigned(138,8) ,
25497	 => std_logic_vector(to_unsigned(133,8) ,
25498	 => std_logic_vector(to_unsigned(133,8) ,
25499	 => std_logic_vector(to_unsigned(142,8) ,
25500	 => std_logic_vector(to_unsigned(111,8) ,
25501	 => std_logic_vector(to_unsigned(25,8) ,
25502	 => std_logic_vector(to_unsigned(11,8) ,
25503	 => std_logic_vector(to_unsigned(9,8) ,
25504	 => std_logic_vector(to_unsigned(11,8) ,
25505	 => std_logic_vector(to_unsigned(8,8) ,
25506	 => std_logic_vector(to_unsigned(7,8) ,
25507	 => std_logic_vector(to_unsigned(10,8) ,
25508	 => std_logic_vector(to_unsigned(6,8) ,
25509	 => std_logic_vector(to_unsigned(3,8) ,
25510	 => std_logic_vector(to_unsigned(4,8) ,
25511	 => std_logic_vector(to_unsigned(5,8) ,
25512	 => std_logic_vector(to_unsigned(7,8) ,
25513	 => std_logic_vector(to_unsigned(12,8) ,
25514	 => std_logic_vector(to_unsigned(9,8) ,
25515	 => std_logic_vector(to_unsigned(27,8) ,
25516	 => std_logic_vector(to_unsigned(127,8) ,
25517	 => std_logic_vector(to_unsigned(173,8) ,
25518	 => std_logic_vector(to_unsigned(138,8) ,
25519	 => std_logic_vector(to_unsigned(133,8) ,
25520	 => std_logic_vector(to_unsigned(151,8) ,
25521	 => std_logic_vector(to_unsigned(136,8) ,
25522	 => std_logic_vector(to_unsigned(152,8) ,
25523	 => std_logic_vector(to_unsigned(112,8) ,
25524	 => std_logic_vector(to_unsigned(24,8) ,
25525	 => std_logic_vector(to_unsigned(8,8) ,
25526	 => std_logic_vector(to_unsigned(4,8) ,
25527	 => std_logic_vector(to_unsigned(5,8) ,
25528	 => std_logic_vector(to_unsigned(7,8) ,
25529	 => std_logic_vector(to_unsigned(10,8) ,
25530	 => std_logic_vector(to_unsigned(9,8) ,
25531	 => std_logic_vector(to_unsigned(10,8) ,
25532	 => std_logic_vector(to_unsigned(10,8) ,
25533	 => std_logic_vector(to_unsigned(6,8) ,
25534	 => std_logic_vector(to_unsigned(11,8) ,
25535	 => std_logic_vector(to_unsigned(11,8) ,
25536	 => std_logic_vector(to_unsigned(9,8) ,
25537	 => std_logic_vector(to_unsigned(6,8) ,
25538	 => std_logic_vector(to_unsigned(12,8) ,
25539	 => std_logic_vector(to_unsigned(73,8) ,
25540	 => std_logic_vector(to_unsigned(97,8) ,
25541	 => std_logic_vector(to_unsigned(76,8) ,
25542	 => std_logic_vector(to_unsigned(100,8) ,
25543	 => std_logic_vector(to_unsigned(151,8) ,
25544	 => std_logic_vector(to_unsigned(171,8) ,
25545	 => std_logic_vector(to_unsigned(159,8) ,
25546	 => std_logic_vector(to_unsigned(168,8) ,
25547	 => std_logic_vector(to_unsigned(171,8) ,
25548	 => std_logic_vector(to_unsigned(163,8) ,
25549	 => std_logic_vector(to_unsigned(166,8) ,
25550	 => std_logic_vector(to_unsigned(149,8) ,
25551	 => std_logic_vector(to_unsigned(125,8) ,
25552	 => std_logic_vector(to_unsigned(78,8) ,
25553	 => std_logic_vector(to_unsigned(58,8) ,
25554	 => std_logic_vector(to_unsigned(70,8) ,
25555	 => std_logic_vector(to_unsigned(70,8) ,
25556	 => std_logic_vector(to_unsigned(73,8) ,
25557	 => std_logic_vector(to_unsigned(27,8) ,
25558	 => std_logic_vector(to_unsigned(1,8) ,
25559	 => std_logic_vector(to_unsigned(3,8) ,
25560	 => std_logic_vector(to_unsigned(6,8) ,
25561	 => std_logic_vector(to_unsigned(8,8) ,
25562	 => std_logic_vector(to_unsigned(10,8) ,
25563	 => std_logic_vector(to_unsigned(12,8) ,
25564	 => std_logic_vector(to_unsigned(16,8) ,
25565	 => std_logic_vector(to_unsigned(9,8) ,
25566	 => std_logic_vector(to_unsigned(16,8) ,
25567	 => std_logic_vector(to_unsigned(112,8) ,
25568	 => std_logic_vector(to_unsigned(114,8) ,
25569	 => std_logic_vector(to_unsigned(11,8) ,
25570	 => std_logic_vector(to_unsigned(5,8) ,
25571	 => std_logic_vector(to_unsigned(60,8) ,
25572	 => std_logic_vector(to_unsigned(97,8) ,
25573	 => std_logic_vector(to_unsigned(104,8) ,
25574	 => std_logic_vector(to_unsigned(105,8) ,
25575	 => std_logic_vector(to_unsigned(142,8) ,
25576	 => std_logic_vector(to_unsigned(164,8) ,
25577	 => std_logic_vector(to_unsigned(147,8) ,
25578	 => std_logic_vector(to_unsigned(124,8) ,
25579	 => std_logic_vector(to_unsigned(111,8) ,
25580	 => std_logic_vector(to_unsigned(103,8) ,
25581	 => std_logic_vector(to_unsigned(101,8) ,
25582	 => std_logic_vector(to_unsigned(100,8) ,
25583	 => std_logic_vector(to_unsigned(92,8) ,
25584	 => std_logic_vector(to_unsigned(93,8) ,
25585	 => std_logic_vector(to_unsigned(100,8) ,
25586	 => std_logic_vector(to_unsigned(105,8) ,
25587	 => std_logic_vector(to_unsigned(112,8) ,
25588	 => std_logic_vector(to_unsigned(109,8) ,
25589	 => std_logic_vector(to_unsigned(118,8) ,
25590	 => std_logic_vector(to_unsigned(130,8) ,
25591	 => std_logic_vector(to_unsigned(127,8) ,
25592	 => std_logic_vector(to_unsigned(127,8) ,
25593	 => std_logic_vector(to_unsigned(142,8) ,
25594	 => std_logic_vector(to_unsigned(163,8) ,
25595	 => std_logic_vector(to_unsigned(171,8) ,
25596	 => std_logic_vector(to_unsigned(166,8) ,
25597	 => std_logic_vector(to_unsigned(142,8) ,
25598	 => std_logic_vector(to_unsigned(128,8) ,
25599	 => std_logic_vector(to_unsigned(115,8) ,
25600	 => std_logic_vector(to_unsigned(112,8) ,
25601	 => std_logic_vector(to_unsigned(161,8) ,
25602	 => std_logic_vector(to_unsigned(161,8) ,
25603	 => std_logic_vector(to_unsigned(157,8) ,
25604	 => std_logic_vector(to_unsigned(152,8) ,
25605	 => std_logic_vector(to_unsigned(159,8) ,
25606	 => std_logic_vector(to_unsigned(147,8) ,
25607	 => std_logic_vector(to_unsigned(38,8) ,
25608	 => std_logic_vector(to_unsigned(11,8) ,
25609	 => std_logic_vector(to_unsigned(25,8) ,
25610	 => std_logic_vector(to_unsigned(18,8) ,
25611	 => std_logic_vector(to_unsigned(10,8) ,
25612	 => std_logic_vector(to_unsigned(8,8) ,
25613	 => std_logic_vector(to_unsigned(6,8) ,
25614	 => std_logic_vector(to_unsigned(53,8) ,
25615	 => std_logic_vector(to_unsigned(107,8) ,
25616	 => std_logic_vector(to_unsigned(74,8) ,
25617	 => std_logic_vector(to_unsigned(63,8) ,
25618	 => std_logic_vector(to_unsigned(35,8) ,
25619	 => std_logic_vector(to_unsigned(2,8) ,
25620	 => std_logic_vector(to_unsigned(0,8) ,
25621	 => std_logic_vector(to_unsigned(15,8) ,
25622	 => std_logic_vector(to_unsigned(67,8) ,
25623	 => std_logic_vector(to_unsigned(30,8) ,
25624	 => std_logic_vector(to_unsigned(28,8) ,
25625	 => std_logic_vector(to_unsigned(31,8) ,
25626	 => std_logic_vector(to_unsigned(38,8) ,
25627	 => std_logic_vector(to_unsigned(69,8) ,
25628	 => std_logic_vector(to_unsigned(139,8) ,
25629	 => std_logic_vector(to_unsigned(161,8) ,
25630	 => std_logic_vector(to_unsigned(66,8) ,
25631	 => std_logic_vector(to_unsigned(19,8) ,
25632	 => std_logic_vector(to_unsigned(9,8) ,
25633	 => std_logic_vector(to_unsigned(3,8) ,
25634	 => std_logic_vector(to_unsigned(1,8) ,
25635	 => std_logic_vector(to_unsigned(0,8) ,
25636	 => std_logic_vector(to_unsigned(2,8) ,
25637	 => std_logic_vector(to_unsigned(3,8) ,
25638	 => std_logic_vector(to_unsigned(4,8) ,
25639	 => std_logic_vector(to_unsigned(2,8) ,
25640	 => std_logic_vector(to_unsigned(6,8) ,
25641	 => std_logic_vector(to_unsigned(109,8) ,
25642	 => std_logic_vector(to_unsigned(163,8) ,
25643	 => std_logic_vector(to_unsigned(139,8) ,
25644	 => std_logic_vector(to_unsigned(114,8) ,
25645	 => std_logic_vector(to_unsigned(50,8) ,
25646	 => std_logic_vector(to_unsigned(16,8) ,
25647	 => std_logic_vector(to_unsigned(2,8) ,
25648	 => std_logic_vector(to_unsigned(0,8) ,
25649	 => std_logic_vector(to_unsigned(4,8) ,
25650	 => std_logic_vector(to_unsigned(125,8) ,
25651	 => std_logic_vector(to_unsigned(173,8) ,
25652	 => std_logic_vector(to_unsigned(161,8) ,
25653	 => std_logic_vector(to_unsigned(161,8) ,
25654	 => std_logic_vector(to_unsigned(154,8) ,
25655	 => std_logic_vector(to_unsigned(164,8) ,
25656	 => std_logic_vector(to_unsigned(142,8) ,
25657	 => std_logic_vector(to_unsigned(22,8) ,
25658	 => std_logic_vector(to_unsigned(7,8) ,
25659	 => std_logic_vector(to_unsigned(18,8) ,
25660	 => std_logic_vector(to_unsigned(10,8) ,
25661	 => std_logic_vector(to_unsigned(3,8) ,
25662	 => std_logic_vector(to_unsigned(8,8) ,
25663	 => std_logic_vector(to_unsigned(9,8) ,
25664	 => std_logic_vector(to_unsigned(3,8) ,
25665	 => std_logic_vector(to_unsigned(4,8) ,
25666	 => std_logic_vector(to_unsigned(5,8) ,
25667	 => std_logic_vector(to_unsigned(4,8) ,
25668	 => std_logic_vector(to_unsigned(4,8) ,
25669	 => std_logic_vector(to_unsigned(3,8) ,
25670	 => std_logic_vector(to_unsigned(5,8) ,
25671	 => std_logic_vector(to_unsigned(5,8) ,
25672	 => std_logic_vector(to_unsigned(5,8) ,
25673	 => std_logic_vector(to_unsigned(9,8) ,
25674	 => std_logic_vector(to_unsigned(4,8) ,
25675	 => std_logic_vector(to_unsigned(0,8) ,
25676	 => std_logic_vector(to_unsigned(18,8) ,
25677	 => std_logic_vector(to_unsigned(78,8) ,
25678	 => std_logic_vector(to_unsigned(116,8) ,
25679	 => std_logic_vector(to_unsigned(146,8) ,
25680	 => std_logic_vector(to_unsigned(175,8) ,
25681	 => std_logic_vector(to_unsigned(130,8) ,
25682	 => std_logic_vector(to_unsigned(7,8) ,
25683	 => std_logic_vector(to_unsigned(18,8) ,
25684	 => std_logic_vector(to_unsigned(37,8) ,
25685	 => std_logic_vector(to_unsigned(12,8) ,
25686	 => std_logic_vector(to_unsigned(4,8) ,
25687	 => std_logic_vector(to_unsigned(81,8) ,
25688	 => std_logic_vector(to_unsigned(163,8) ,
25689	 => std_logic_vector(to_unsigned(116,8) ,
25690	 => std_logic_vector(to_unsigned(127,8) ,
25691	 => std_logic_vector(to_unsigned(97,8) ,
25692	 => std_logic_vector(to_unsigned(77,8) ,
25693	 => std_logic_vector(to_unsigned(144,8) ,
25694	 => std_logic_vector(to_unsigned(166,8) ,
25695	 => std_logic_vector(to_unsigned(163,8) ,
25696	 => std_logic_vector(to_unsigned(161,8) ,
25697	 => std_logic_vector(to_unsigned(157,8) ,
25698	 => std_logic_vector(to_unsigned(163,8) ,
25699	 => std_logic_vector(to_unsigned(149,8) ,
25700	 => std_logic_vector(to_unsigned(152,8) ,
25701	 => std_logic_vector(to_unsigned(141,8) ,
25702	 => std_logic_vector(to_unsigned(40,8) ,
25703	 => std_logic_vector(to_unsigned(55,8) ,
25704	 => std_logic_vector(to_unsigned(87,8) ,
25705	 => std_logic_vector(to_unsigned(92,8) ,
25706	 => std_logic_vector(to_unsigned(101,8) ,
25707	 => std_logic_vector(to_unsigned(133,8) ,
25708	 => std_logic_vector(to_unsigned(149,8) ,
25709	 => std_logic_vector(to_unsigned(91,8) ,
25710	 => std_logic_vector(to_unsigned(30,8) ,
25711	 => std_logic_vector(to_unsigned(52,8) ,
25712	 => std_logic_vector(to_unsigned(68,8) ,
25713	 => std_logic_vector(to_unsigned(58,8) ,
25714	 => std_logic_vector(to_unsigned(4,8) ,
25715	 => std_logic_vector(to_unsigned(2,8) ,
25716	 => std_logic_vector(to_unsigned(4,8) ,
25717	 => std_logic_vector(to_unsigned(19,8) ,
25718	 => std_logic_vector(to_unsigned(35,8) ,
25719	 => std_logic_vector(to_unsigned(8,8) ,
25720	 => std_logic_vector(to_unsigned(1,8) ,
25721	 => std_logic_vector(to_unsigned(1,8) ,
25722	 => std_logic_vector(to_unsigned(1,8) ,
25723	 => std_logic_vector(to_unsigned(0,8) ,
25724	 => std_logic_vector(to_unsigned(2,8) ,
25725	 => std_logic_vector(to_unsigned(13,8) ,
25726	 => std_logic_vector(to_unsigned(24,8) ,
25727	 => std_logic_vector(to_unsigned(3,8) ,
25728	 => std_logic_vector(to_unsigned(2,8) ,
25729	 => std_logic_vector(to_unsigned(10,8) ,
25730	 => std_logic_vector(to_unsigned(35,8) ,
25731	 => std_logic_vector(to_unsigned(99,8) ,
25732	 => std_logic_vector(to_unsigned(136,8) ,
25733	 => std_logic_vector(to_unsigned(141,8) ,
25734	 => std_logic_vector(to_unsigned(136,8) ,
25735	 => std_logic_vector(to_unsigned(147,8) ,
25736	 => std_logic_vector(to_unsigned(156,8) ,
25737	 => std_logic_vector(to_unsigned(154,8) ,
25738	 => std_logic_vector(to_unsigned(87,8) ,
25739	 => std_logic_vector(to_unsigned(32,8) ,
25740	 => std_logic_vector(to_unsigned(22,8) ,
25741	 => std_logic_vector(to_unsigned(9,8) ,
25742	 => std_logic_vector(to_unsigned(6,8) ,
25743	 => std_logic_vector(to_unsigned(1,8) ,
25744	 => std_logic_vector(to_unsigned(3,8) ,
25745	 => std_logic_vector(to_unsigned(15,8) ,
25746	 => std_logic_vector(to_unsigned(16,8) ,
25747	 => std_logic_vector(to_unsigned(10,8) ,
25748	 => std_logic_vector(to_unsigned(12,8) ,
25749	 => std_logic_vector(to_unsigned(10,8) ,
25750	 => std_logic_vector(to_unsigned(25,8) ,
25751	 => std_logic_vector(to_unsigned(13,8) ,
25752	 => std_logic_vector(to_unsigned(2,8) ,
25753	 => std_logic_vector(to_unsigned(32,8) ,
25754	 => std_logic_vector(to_unsigned(43,8) ,
25755	 => std_logic_vector(to_unsigned(34,8) ,
25756	 => std_logic_vector(to_unsigned(30,8) ,
25757	 => std_logic_vector(to_unsigned(20,8) ,
25758	 => std_logic_vector(to_unsigned(30,8) ,
25759	 => std_logic_vector(to_unsigned(32,8) ,
25760	 => std_logic_vector(to_unsigned(30,8) ,
25761	 => std_logic_vector(to_unsigned(41,8) ,
25762	 => std_logic_vector(to_unsigned(41,8) ,
25763	 => std_logic_vector(to_unsigned(22,8) ,
25764	 => std_logic_vector(to_unsigned(16,8) ,
25765	 => std_logic_vector(to_unsigned(32,8) ,
25766	 => std_logic_vector(to_unsigned(21,8) ,
25767	 => std_logic_vector(to_unsigned(19,8) ,
25768	 => std_logic_vector(to_unsigned(25,8) ,
25769	 => std_logic_vector(to_unsigned(25,8) ,
25770	 => std_logic_vector(to_unsigned(17,8) ,
25771	 => std_logic_vector(to_unsigned(12,8) ,
25772	 => std_logic_vector(to_unsigned(21,8) ,
25773	 => std_logic_vector(to_unsigned(32,8) ,
25774	 => std_logic_vector(to_unsigned(19,8) ,
25775	 => std_logic_vector(to_unsigned(17,8) ,
25776	 => std_logic_vector(to_unsigned(21,8) ,
25777	 => std_logic_vector(to_unsigned(23,8) ,
25778	 => std_logic_vector(to_unsigned(34,8) ,
25779	 => std_logic_vector(to_unsigned(33,8) ,
25780	 => std_logic_vector(to_unsigned(26,8) ,
25781	 => std_logic_vector(to_unsigned(17,8) ,
25782	 => std_logic_vector(to_unsigned(8,8) ,
25783	 => std_logic_vector(to_unsigned(6,8) ,
25784	 => std_logic_vector(to_unsigned(9,8) ,
25785	 => std_logic_vector(to_unsigned(10,8) ,
25786	 => std_logic_vector(to_unsigned(7,8) ,
25787	 => std_logic_vector(to_unsigned(9,8) ,
25788	 => std_logic_vector(to_unsigned(91,8) ,
25789	 => std_logic_vector(to_unsigned(101,8) ,
25790	 => std_logic_vector(to_unsigned(96,8) ,
25791	 => std_logic_vector(to_unsigned(105,8) ,
25792	 => std_logic_vector(to_unsigned(109,8) ,
25793	 => std_logic_vector(to_unsigned(76,8) ,
25794	 => std_logic_vector(to_unsigned(107,8) ,
25795	 => std_logic_vector(to_unsigned(81,8) ,
25796	 => std_logic_vector(to_unsigned(4,8) ,
25797	 => std_logic_vector(to_unsigned(3,8) ,
25798	 => std_logic_vector(to_unsigned(6,8) ,
25799	 => std_logic_vector(to_unsigned(5,8) ,
25800	 => std_logic_vector(to_unsigned(6,8) ,
25801	 => std_logic_vector(to_unsigned(8,8) ,
25802	 => std_logic_vector(to_unsigned(4,8) ,
25803	 => std_logic_vector(to_unsigned(7,8) ,
25804	 => std_logic_vector(to_unsigned(45,8) ,
25805	 => std_logic_vector(to_unsigned(151,8) ,
25806	 => std_logic_vector(to_unsigned(154,8) ,
25807	 => std_logic_vector(to_unsigned(133,8) ,
25808	 => std_logic_vector(to_unsigned(146,8) ,
25809	 => std_logic_vector(to_unsigned(152,8) ,
25810	 => std_logic_vector(to_unsigned(152,8) ,
25811	 => std_logic_vector(to_unsigned(159,8) ,
25812	 => std_logic_vector(to_unsigned(157,8) ,
25813	 => std_logic_vector(to_unsigned(139,8) ,
25814	 => std_logic_vector(to_unsigned(144,8) ,
25815	 => std_logic_vector(to_unsigned(151,8) ,
25816	 => std_logic_vector(to_unsigned(144,8) ,
25817	 => std_logic_vector(to_unsigned(141,8) ,
25818	 => std_logic_vector(to_unsigned(139,8) ,
25819	 => std_logic_vector(to_unsigned(156,8) ,
25820	 => std_logic_vector(to_unsigned(73,8) ,
25821	 => std_logic_vector(to_unsigned(9,8) ,
25822	 => std_logic_vector(to_unsigned(6,8) ,
25823	 => std_logic_vector(to_unsigned(7,8) ,
25824	 => std_logic_vector(to_unsigned(8,8) ,
25825	 => std_logic_vector(to_unsigned(45,8) ,
25826	 => std_logic_vector(to_unsigned(20,8) ,
25827	 => std_logic_vector(to_unsigned(3,8) ,
25828	 => std_logic_vector(to_unsigned(3,8) ,
25829	 => std_logic_vector(to_unsigned(3,8) ,
25830	 => std_logic_vector(to_unsigned(6,8) ,
25831	 => std_logic_vector(to_unsigned(7,8) ,
25832	 => std_logic_vector(to_unsigned(8,8) ,
25833	 => std_logic_vector(to_unsigned(12,8) ,
25834	 => std_logic_vector(to_unsigned(8,8) ,
25835	 => std_logic_vector(to_unsigned(34,8) ,
25836	 => std_logic_vector(to_unsigned(164,8) ,
25837	 => std_logic_vector(to_unsigned(163,8) ,
25838	 => std_logic_vector(to_unsigned(66,8) ,
25839	 => std_logic_vector(to_unsigned(79,8) ,
25840	 => std_logic_vector(to_unsigned(136,8) ,
25841	 => std_logic_vector(to_unsigned(142,8) ,
25842	 => std_logic_vector(to_unsigned(141,8) ,
25843	 => std_logic_vector(to_unsigned(157,8) ,
25844	 => std_logic_vector(to_unsigned(142,8) ,
25845	 => std_logic_vector(to_unsigned(32,8) ,
25846	 => std_logic_vector(to_unsigned(2,8) ,
25847	 => std_logic_vector(to_unsigned(5,8) ,
25848	 => std_logic_vector(to_unsigned(7,8) ,
25849	 => std_logic_vector(to_unsigned(8,8) ,
25850	 => std_logic_vector(to_unsigned(8,8) ,
25851	 => std_logic_vector(to_unsigned(15,8) ,
25852	 => std_logic_vector(to_unsigned(12,8) ,
25853	 => std_logic_vector(to_unsigned(4,8) ,
25854	 => std_logic_vector(to_unsigned(6,8) ,
25855	 => std_logic_vector(to_unsigned(11,8) ,
25856	 => std_logic_vector(to_unsigned(9,8) ,
25857	 => std_logic_vector(to_unsigned(6,8) ,
25858	 => std_logic_vector(to_unsigned(10,8) ,
25859	 => std_logic_vector(to_unsigned(51,8) ,
25860	 => std_logic_vector(to_unsigned(43,8) ,
25861	 => std_logic_vector(to_unsigned(10,8) ,
25862	 => std_logic_vector(to_unsigned(10,8) ,
25863	 => std_logic_vector(to_unsigned(68,8) ,
25864	 => std_logic_vector(to_unsigned(170,8) ,
25865	 => std_logic_vector(to_unsigned(170,8) ,
25866	 => std_logic_vector(to_unsigned(171,8) ,
25867	 => std_logic_vector(to_unsigned(163,8) ,
25868	 => std_logic_vector(to_unsigned(170,8) ,
25869	 => std_logic_vector(to_unsigned(170,8) ,
25870	 => std_logic_vector(to_unsigned(104,8) ,
25871	 => std_logic_vector(to_unsigned(68,8) ,
25872	 => std_logic_vector(to_unsigned(64,8) ,
25873	 => std_logic_vector(to_unsigned(107,8) ,
25874	 => std_logic_vector(to_unsigned(144,8) ,
25875	 => std_logic_vector(to_unsigned(97,8) ,
25876	 => std_logic_vector(to_unsigned(35,8) ,
25877	 => std_logic_vector(to_unsigned(24,8) ,
25878	 => std_logic_vector(to_unsigned(12,8) ,
25879	 => std_logic_vector(to_unsigned(2,8) ,
25880	 => std_logic_vector(to_unsigned(4,8) ,
25881	 => std_logic_vector(to_unsigned(3,8) ,
25882	 => std_logic_vector(to_unsigned(5,8) ,
25883	 => std_logic_vector(to_unsigned(9,8) ,
25884	 => std_logic_vector(to_unsigned(9,8) ,
25885	 => std_logic_vector(to_unsigned(12,8) ,
25886	 => std_logic_vector(to_unsigned(58,8) ,
25887	 => std_logic_vector(to_unsigned(144,8) ,
25888	 => std_logic_vector(to_unsigned(118,8) ,
25889	 => std_logic_vector(to_unsigned(12,8) ,
25890	 => std_logic_vector(to_unsigned(2,8) ,
25891	 => std_logic_vector(to_unsigned(57,8) ,
25892	 => std_logic_vector(to_unsigned(105,8) ,
25893	 => std_logic_vector(to_unsigned(90,8) ,
25894	 => std_logic_vector(to_unsigned(70,8) ,
25895	 => std_logic_vector(to_unsigned(119,8) ,
25896	 => std_logic_vector(to_unsigned(159,8) ,
25897	 => std_logic_vector(to_unsigned(149,8) ,
25898	 => std_logic_vector(to_unsigned(131,8) ,
25899	 => std_logic_vector(to_unsigned(114,8) ,
25900	 => std_logic_vector(to_unsigned(101,8) ,
25901	 => std_logic_vector(to_unsigned(103,8) ,
25902	 => std_logic_vector(to_unsigned(104,8) ,
25903	 => std_logic_vector(to_unsigned(96,8) ,
25904	 => std_logic_vector(to_unsigned(96,8) ,
25905	 => std_logic_vector(to_unsigned(96,8) ,
25906	 => std_logic_vector(to_unsigned(104,8) ,
25907	 => std_logic_vector(to_unsigned(116,8) ,
25908	 => std_logic_vector(to_unsigned(105,8) ,
25909	 => std_logic_vector(to_unsigned(121,8) ,
25910	 => std_logic_vector(to_unsigned(131,8) ,
25911	 => std_logic_vector(to_unsigned(133,8) ,
25912	 => std_logic_vector(to_unsigned(128,8) ,
25913	 => std_logic_vector(to_unsigned(128,8) ,
25914	 => std_logic_vector(to_unsigned(157,8) ,
25915	 => std_logic_vector(to_unsigned(170,8) ,
25916	 => std_logic_vector(to_unsigned(168,8) ,
25917	 => std_logic_vector(to_unsigned(164,8) ,
25918	 => std_logic_vector(to_unsigned(136,8) ,
25919	 => std_logic_vector(to_unsigned(121,8) ,
25920	 => std_logic_vector(to_unsigned(116,8) ,
25921	 => std_logic_vector(to_unsigned(159,8) ,
25922	 => std_logic_vector(to_unsigned(157,8) ,
25923	 => std_logic_vector(to_unsigned(161,8) ,
25924	 => std_logic_vector(to_unsigned(156,8) ,
25925	 => std_logic_vector(to_unsigned(163,8) ,
25926	 => std_logic_vector(to_unsigned(146,8) ,
25927	 => std_logic_vector(to_unsigned(22,8) ,
25928	 => std_logic_vector(to_unsigned(7,8) ,
25929	 => std_logic_vector(to_unsigned(29,8) ,
25930	 => std_logic_vector(to_unsigned(37,8) ,
25931	 => std_logic_vector(to_unsigned(61,8) ,
25932	 => std_logic_vector(to_unsigned(53,8) ,
25933	 => std_logic_vector(to_unsigned(48,8) ,
25934	 => std_logic_vector(to_unsigned(87,8) ,
25935	 => std_logic_vector(to_unsigned(105,8) ,
25936	 => std_logic_vector(to_unsigned(40,8) ,
25937	 => std_logic_vector(to_unsigned(9,8) ,
25938	 => std_logic_vector(to_unsigned(5,8) ,
25939	 => std_logic_vector(to_unsigned(0,8) ,
25940	 => std_logic_vector(to_unsigned(1,8) ,
25941	 => std_logic_vector(to_unsigned(2,8) ,
25942	 => std_logic_vector(to_unsigned(8,8) ,
25943	 => std_logic_vector(to_unsigned(7,8) ,
25944	 => std_logic_vector(to_unsigned(4,8) ,
25945	 => std_logic_vector(to_unsigned(4,8) ,
25946	 => std_logic_vector(to_unsigned(3,8) ,
25947	 => std_logic_vector(to_unsigned(5,8) ,
25948	 => std_logic_vector(to_unsigned(35,8) ,
25949	 => std_logic_vector(to_unsigned(107,8) ,
25950	 => std_logic_vector(to_unsigned(161,8) ,
25951	 => std_logic_vector(to_unsigned(151,8) ,
25952	 => std_logic_vector(to_unsigned(103,8) ,
25953	 => std_logic_vector(to_unsigned(38,8) ,
25954	 => std_logic_vector(to_unsigned(6,8) ,
25955	 => std_logic_vector(to_unsigned(1,8) ,
25956	 => std_logic_vector(to_unsigned(0,8) ,
25957	 => std_logic_vector(to_unsigned(0,8) ,
25958	 => std_logic_vector(to_unsigned(2,8) ,
25959	 => std_logic_vector(to_unsigned(1,8) ,
25960	 => std_logic_vector(to_unsigned(5,8) ,
25961	 => std_logic_vector(to_unsigned(111,8) ,
25962	 => std_logic_vector(to_unsigned(147,8) ,
25963	 => std_logic_vector(to_unsigned(124,8) ,
25964	 => std_logic_vector(to_unsigned(85,8) ,
25965	 => std_logic_vector(to_unsigned(26,8) ,
25966	 => std_logic_vector(to_unsigned(4,8) ,
25967	 => std_logic_vector(to_unsigned(1,8) ,
25968	 => std_logic_vector(to_unsigned(0,8) ,
25969	 => std_logic_vector(to_unsigned(14,8) ,
25970	 => std_logic_vector(to_unsigned(161,8) ,
25971	 => std_logic_vector(to_unsigned(170,8) ,
25972	 => std_logic_vector(to_unsigned(157,8) ,
25973	 => std_logic_vector(to_unsigned(161,8) ,
25974	 => std_logic_vector(to_unsigned(161,8) ,
25975	 => std_logic_vector(to_unsigned(163,8) ,
25976	 => std_logic_vector(to_unsigned(163,8) ,
25977	 => std_logic_vector(to_unsigned(41,8) ,
25978	 => std_logic_vector(to_unsigned(5,8) ,
25979	 => std_logic_vector(to_unsigned(17,8) ,
25980	 => std_logic_vector(to_unsigned(11,8) ,
25981	 => std_logic_vector(to_unsigned(6,8) ,
25982	 => std_logic_vector(to_unsigned(4,8) ,
25983	 => std_logic_vector(to_unsigned(9,8) ,
25984	 => std_logic_vector(to_unsigned(9,8) ,
25985	 => std_logic_vector(to_unsigned(4,8) ,
25986	 => std_logic_vector(to_unsigned(4,8) ,
25987	 => std_logic_vector(to_unsigned(5,8) ,
25988	 => std_logic_vector(to_unsigned(3,8) ,
25989	 => std_logic_vector(to_unsigned(4,8) ,
25990	 => std_logic_vector(to_unsigned(4,8) ,
25991	 => std_logic_vector(to_unsigned(4,8) ,
25992	 => std_logic_vector(to_unsigned(4,8) ,
25993	 => std_logic_vector(to_unsigned(8,8) ,
25994	 => std_logic_vector(to_unsigned(5,8) ,
25995	 => std_logic_vector(to_unsigned(1,8) ,
25996	 => std_logic_vector(to_unsigned(2,8) ,
25997	 => std_logic_vector(to_unsigned(57,8) ,
25998	 => std_logic_vector(to_unsigned(144,8) ,
25999	 => std_logic_vector(to_unsigned(142,8) ,
26000	 => std_logic_vector(to_unsigned(171,8) ,
26001	 => std_logic_vector(to_unsigned(131,8) ,
26002	 => std_logic_vector(to_unsigned(26,8) ,
26003	 => std_logic_vector(to_unsigned(41,8) ,
26004	 => std_logic_vector(to_unsigned(32,8) ,
26005	 => std_logic_vector(to_unsigned(3,8) ,
26006	 => std_logic_vector(to_unsigned(10,8) ,
26007	 => std_logic_vector(to_unsigned(141,8) ,
26008	 => std_logic_vector(to_unsigned(175,8) ,
26009	 => std_logic_vector(to_unsigned(107,8) ,
26010	 => std_logic_vector(to_unsigned(86,8) ,
26011	 => std_logic_vector(to_unsigned(121,8) ,
26012	 => std_logic_vector(to_unsigned(100,8) ,
26013	 => std_logic_vector(to_unsigned(128,8) ,
26014	 => std_logic_vector(to_unsigned(164,8) ,
26015	 => std_logic_vector(to_unsigned(161,8) ,
26016	 => std_logic_vector(to_unsigned(157,8) ,
26017	 => std_logic_vector(to_unsigned(152,8) ,
26018	 => std_logic_vector(to_unsigned(152,8) ,
26019	 => std_logic_vector(to_unsigned(147,8) ,
26020	 => std_logic_vector(to_unsigned(159,8) ,
26021	 => std_logic_vector(to_unsigned(128,8) ,
26022	 => std_logic_vector(to_unsigned(68,8) ,
26023	 => std_logic_vector(to_unsigned(76,8) ,
26024	 => std_logic_vector(to_unsigned(99,8) ,
26025	 => std_logic_vector(to_unsigned(76,8) ,
26026	 => std_logic_vector(to_unsigned(79,8) ,
26027	 => std_logic_vector(to_unsigned(114,8) ,
26028	 => std_logic_vector(to_unsigned(111,8) ,
26029	 => std_logic_vector(to_unsigned(61,8) ,
26030	 => std_logic_vector(to_unsigned(18,8) ,
26031	 => std_logic_vector(to_unsigned(29,8) ,
26032	 => std_logic_vector(to_unsigned(45,8) ,
26033	 => std_logic_vector(to_unsigned(16,8) ,
26034	 => std_logic_vector(to_unsigned(2,8) ,
26035	 => std_logic_vector(to_unsigned(2,8) ,
26036	 => std_logic_vector(to_unsigned(0,8) ,
26037	 => std_logic_vector(to_unsigned(6,8) ,
26038	 => std_logic_vector(to_unsigned(53,8) ,
26039	 => std_logic_vector(to_unsigned(26,8) ,
26040	 => std_logic_vector(to_unsigned(3,8) ,
26041	 => std_logic_vector(to_unsigned(1,8) ,
26042	 => std_logic_vector(to_unsigned(0,8) ,
26043	 => std_logic_vector(to_unsigned(4,8) ,
26044	 => std_logic_vector(to_unsigned(12,8) ,
26045	 => std_logic_vector(to_unsigned(12,8) ,
26046	 => std_logic_vector(to_unsigned(11,8) ,
26047	 => std_logic_vector(to_unsigned(2,8) ,
26048	 => std_logic_vector(to_unsigned(4,8) ,
26049	 => std_logic_vector(to_unsigned(15,8) ,
26050	 => std_logic_vector(to_unsigned(51,8) ,
26051	 => std_logic_vector(to_unsigned(119,8) ,
26052	 => std_logic_vector(to_unsigned(122,8) ,
26053	 => std_logic_vector(to_unsigned(115,8) ,
26054	 => std_logic_vector(to_unsigned(90,8) ,
26055	 => std_logic_vector(to_unsigned(97,8) ,
26056	 => std_logic_vector(to_unsigned(157,8) ,
26057	 => std_logic_vector(to_unsigned(139,8) ,
26058	 => std_logic_vector(to_unsigned(49,8) ,
26059	 => std_logic_vector(to_unsigned(26,8) ,
26060	 => std_logic_vector(to_unsigned(27,8) ,
26061	 => std_logic_vector(to_unsigned(20,8) ,
26062	 => std_logic_vector(to_unsigned(15,8) ,
26063	 => std_logic_vector(to_unsigned(5,8) ,
26064	 => std_logic_vector(to_unsigned(3,8) ,
26065	 => std_logic_vector(to_unsigned(6,8) ,
26066	 => std_logic_vector(to_unsigned(18,8) ,
26067	 => std_logic_vector(to_unsigned(13,8) ,
26068	 => std_logic_vector(to_unsigned(8,8) ,
26069	 => std_logic_vector(to_unsigned(28,8) ,
26070	 => std_logic_vector(to_unsigned(38,8) ,
26071	 => std_logic_vector(to_unsigned(13,8) ,
26072	 => std_logic_vector(to_unsigned(4,8) ,
26073	 => std_logic_vector(to_unsigned(5,8) ,
26074	 => std_logic_vector(to_unsigned(13,8) ,
26075	 => std_logic_vector(to_unsigned(17,8) ,
26076	 => std_logic_vector(to_unsigned(24,8) ,
26077	 => std_logic_vector(to_unsigned(30,8) ,
26078	 => std_logic_vector(to_unsigned(30,8) ,
26079	 => std_logic_vector(to_unsigned(35,8) ,
26080	 => std_logic_vector(to_unsigned(39,8) ,
26081	 => std_logic_vector(to_unsigned(44,8) ,
26082	 => std_logic_vector(to_unsigned(37,8) ,
26083	 => std_logic_vector(to_unsigned(17,8) ,
26084	 => std_logic_vector(to_unsigned(17,8) ,
26085	 => std_logic_vector(to_unsigned(37,8) ,
26086	 => std_logic_vector(to_unsigned(13,8) ,
26087	 => std_logic_vector(to_unsigned(5,8) ,
26088	 => std_logic_vector(to_unsigned(17,8) ,
26089	 => std_logic_vector(to_unsigned(24,8) ,
26090	 => std_logic_vector(to_unsigned(22,8) ,
26091	 => std_logic_vector(to_unsigned(14,8) ,
26092	 => std_logic_vector(to_unsigned(18,8) ,
26093	 => std_logic_vector(to_unsigned(25,8) ,
26094	 => std_logic_vector(to_unsigned(19,8) ,
26095	 => std_logic_vector(to_unsigned(21,8) ,
26096	 => std_logic_vector(to_unsigned(27,8) ,
26097	 => std_logic_vector(to_unsigned(27,8) ,
26098	 => std_logic_vector(to_unsigned(35,8) ,
26099	 => std_logic_vector(to_unsigned(35,8) ,
26100	 => std_logic_vector(to_unsigned(29,8) ,
26101	 => std_logic_vector(to_unsigned(17,8) ,
26102	 => std_logic_vector(to_unsigned(5,8) ,
26103	 => std_logic_vector(to_unsigned(2,8) ,
26104	 => std_logic_vector(to_unsigned(8,8) ,
26105	 => std_logic_vector(to_unsigned(15,8) ,
26106	 => std_logic_vector(to_unsigned(7,8) ,
26107	 => std_logic_vector(to_unsigned(21,8) ,
26108	 => std_logic_vector(to_unsigned(109,8) ,
26109	 => std_logic_vector(to_unsigned(97,8) ,
26110	 => std_logic_vector(to_unsigned(116,8) ,
26111	 => std_logic_vector(to_unsigned(130,8) ,
26112	 => std_logic_vector(to_unsigned(127,8) ,
26113	 => std_logic_vector(to_unsigned(125,8) ,
26114	 => std_logic_vector(to_unsigned(136,8) ,
26115	 => std_logic_vector(to_unsigned(101,8) ,
26116	 => std_logic_vector(to_unsigned(13,8) ,
26117	 => std_logic_vector(to_unsigned(2,8) ,
26118	 => std_logic_vector(to_unsigned(6,8) ,
26119	 => std_logic_vector(to_unsigned(6,8) ,
26120	 => std_logic_vector(to_unsigned(11,8) ,
26121	 => std_logic_vector(to_unsigned(16,8) ,
26122	 => std_logic_vector(to_unsigned(13,8) ,
26123	 => std_logic_vector(to_unsigned(17,8) ,
26124	 => std_logic_vector(to_unsigned(86,8) ,
26125	 => std_logic_vector(to_unsigned(159,8) ,
26126	 => std_logic_vector(to_unsigned(142,8) ,
26127	 => std_logic_vector(to_unsigned(141,8) ,
26128	 => std_logic_vector(to_unsigned(159,8) ,
26129	 => std_logic_vector(to_unsigned(151,8) ,
26130	 => std_logic_vector(to_unsigned(142,8) ,
26131	 => std_logic_vector(to_unsigned(154,8) ,
26132	 => std_logic_vector(to_unsigned(157,8) ,
26133	 => std_logic_vector(to_unsigned(142,8) ,
26134	 => std_logic_vector(to_unsigned(141,8) ,
26135	 => std_logic_vector(to_unsigned(146,8) ,
26136	 => std_logic_vector(to_unsigned(144,8) ,
26137	 => std_logic_vector(to_unsigned(142,8) ,
26138	 => std_logic_vector(to_unsigned(146,8) ,
26139	 => std_logic_vector(to_unsigned(136,8) ,
26140	 => std_logic_vector(to_unsigned(30,8) ,
26141	 => std_logic_vector(to_unsigned(7,8) ,
26142	 => std_logic_vector(to_unsigned(8,8) ,
26143	 => std_logic_vector(to_unsigned(5,8) ,
26144	 => std_logic_vector(to_unsigned(14,8) ,
26145	 => std_logic_vector(to_unsigned(97,8) ,
26146	 => std_logic_vector(to_unsigned(25,8) ,
26147	 => std_logic_vector(to_unsigned(5,8) ,
26148	 => std_logic_vector(to_unsigned(5,8) ,
26149	 => std_logic_vector(to_unsigned(4,8) ,
26150	 => std_logic_vector(to_unsigned(6,8) ,
26151	 => std_logic_vector(to_unsigned(6,8) ,
26152	 => std_logic_vector(to_unsigned(10,8) ,
26153	 => std_logic_vector(to_unsigned(10,8) ,
26154	 => std_logic_vector(to_unsigned(14,8) ,
26155	 => std_logic_vector(to_unsigned(91,8) ,
26156	 => std_logic_vector(to_unsigned(188,8) ,
26157	 => std_logic_vector(to_unsigned(88,8) ,
26158	 => std_logic_vector(to_unsigned(32,8) ,
26159	 => std_logic_vector(to_unsigned(59,8) ,
26160	 => std_logic_vector(to_unsigned(96,8) ,
26161	 => std_logic_vector(to_unsigned(130,8) ,
26162	 => std_logic_vector(to_unsigned(147,8) ,
26163	 => std_logic_vector(to_unsigned(86,8) ,
26164	 => std_logic_vector(to_unsigned(30,8) ,
26165	 => std_logic_vector(to_unsigned(11,8) ,
26166	 => std_logic_vector(to_unsigned(3,8) ,
26167	 => std_logic_vector(to_unsigned(3,8) ,
26168	 => std_logic_vector(to_unsigned(5,8) ,
26169	 => std_logic_vector(to_unsigned(8,8) ,
26170	 => std_logic_vector(to_unsigned(10,8) ,
26171	 => std_logic_vector(to_unsigned(10,8) ,
26172	 => std_logic_vector(to_unsigned(6,8) ,
26173	 => std_logic_vector(to_unsigned(7,8) ,
26174	 => std_logic_vector(to_unsigned(8,8) ,
26175	 => std_logic_vector(to_unsigned(9,8) ,
26176	 => std_logic_vector(to_unsigned(12,8) ,
26177	 => std_logic_vector(to_unsigned(8,8) ,
26178	 => std_logic_vector(to_unsigned(7,8) ,
26179	 => std_logic_vector(to_unsigned(29,8) ,
26180	 => std_logic_vector(to_unsigned(25,8) ,
26181	 => std_logic_vector(to_unsigned(8,8) ,
26182	 => std_logic_vector(to_unsigned(9,8) ,
26183	 => std_logic_vector(to_unsigned(61,8) ,
26184	 => std_logic_vector(to_unsigned(124,8) ,
26185	 => std_logic_vector(to_unsigned(136,8) ,
26186	 => std_logic_vector(to_unsigned(168,8) ,
26187	 => std_logic_vector(to_unsigned(168,8) ,
26188	 => std_logic_vector(to_unsigned(173,8) ,
26189	 => std_logic_vector(to_unsigned(152,8) ,
26190	 => std_logic_vector(to_unsigned(85,8) ,
26191	 => std_logic_vector(to_unsigned(62,8) ,
26192	 => std_logic_vector(to_unsigned(99,8) ,
26193	 => std_logic_vector(to_unsigned(124,8) ,
26194	 => std_logic_vector(to_unsigned(99,8) ,
26195	 => std_logic_vector(to_unsigned(41,8) ,
26196	 => std_logic_vector(to_unsigned(1,8) ,
26197	 => std_logic_vector(to_unsigned(2,8) ,
26198	 => std_logic_vector(to_unsigned(18,8) ,
26199	 => std_logic_vector(to_unsigned(11,8) ,
26200	 => std_logic_vector(to_unsigned(3,8) ,
26201	 => std_logic_vector(to_unsigned(3,8) ,
26202	 => std_logic_vector(to_unsigned(2,8) ,
26203	 => std_logic_vector(to_unsigned(6,8) ,
26204	 => std_logic_vector(to_unsigned(37,8) ,
26205	 => std_logic_vector(to_unsigned(22,8) ,
26206	 => std_logic_vector(to_unsigned(7,8) ,
26207	 => std_logic_vector(to_unsigned(115,8) ,
26208	 => std_logic_vector(to_unsigned(146,8) ,
26209	 => std_logic_vector(to_unsigned(15,8) ,
26210	 => std_logic_vector(to_unsigned(5,8) ,
26211	 => std_logic_vector(to_unsigned(51,8) ,
26212	 => std_logic_vector(to_unsigned(81,8) ,
26213	 => std_logic_vector(to_unsigned(81,8) ,
26214	 => std_logic_vector(to_unsigned(111,8) ,
26215	 => std_logic_vector(to_unsigned(138,8) ,
26216	 => std_logic_vector(to_unsigned(125,8) ,
26217	 => std_logic_vector(to_unsigned(93,8) ,
26218	 => std_logic_vector(to_unsigned(100,8) ,
26219	 => std_logic_vector(to_unsigned(119,8) ,
26220	 => std_logic_vector(to_unsigned(99,8) ,
26221	 => std_logic_vector(to_unsigned(101,8) ,
26222	 => std_logic_vector(to_unsigned(109,8) ,
26223	 => std_logic_vector(to_unsigned(103,8) ,
26224	 => std_logic_vector(to_unsigned(103,8) ,
26225	 => std_logic_vector(to_unsigned(95,8) ,
26226	 => std_logic_vector(to_unsigned(116,8) ,
26227	 => std_logic_vector(to_unsigned(130,8) ,
26228	 => std_logic_vector(to_unsigned(109,8) ,
26229	 => std_logic_vector(to_unsigned(115,8) ,
26230	 => std_logic_vector(to_unsigned(138,8) ,
26231	 => std_logic_vector(to_unsigned(136,8) ,
26232	 => std_logic_vector(to_unsigned(131,8) ,
26233	 => std_logic_vector(to_unsigned(127,8) ,
26234	 => std_logic_vector(to_unsigned(144,8) ,
26235	 => std_logic_vector(to_unsigned(170,8) ,
26236	 => std_logic_vector(to_unsigned(164,8) ,
26237	 => std_logic_vector(to_unsigned(164,8) ,
26238	 => std_logic_vector(to_unsigned(144,8) ,
26239	 => std_logic_vector(to_unsigned(119,8) ,
26240	 => std_logic_vector(to_unsigned(109,8) ,
26241	 => std_logic_vector(to_unsigned(164,8) ,
26242	 => std_logic_vector(to_unsigned(159,8) ,
26243	 => std_logic_vector(to_unsigned(159,8) ,
26244	 => std_logic_vector(to_unsigned(159,8) ,
26245	 => std_logic_vector(to_unsigned(166,8) ,
26246	 => std_logic_vector(to_unsigned(156,8) ,
26247	 => std_logic_vector(to_unsigned(28,8) ,
26248	 => std_logic_vector(to_unsigned(15,8) ,
26249	 => std_logic_vector(to_unsigned(22,8) ,
26250	 => std_logic_vector(to_unsigned(49,8) ,
26251	 => std_logic_vector(to_unsigned(66,8) ,
26252	 => std_logic_vector(to_unsigned(60,8) ,
26253	 => std_logic_vector(to_unsigned(56,8) ,
26254	 => std_logic_vector(to_unsigned(14,8) ,
26255	 => std_logic_vector(to_unsigned(11,8) ,
26256	 => std_logic_vector(to_unsigned(15,8) ,
26257	 => std_logic_vector(to_unsigned(3,8) ,
26258	 => std_logic_vector(to_unsigned(0,8) ,
26259	 => std_logic_vector(to_unsigned(0,8) ,
26260	 => std_logic_vector(to_unsigned(2,8) ,
26261	 => std_logic_vector(to_unsigned(4,8) ,
26262	 => std_logic_vector(to_unsigned(3,8) ,
26263	 => std_logic_vector(to_unsigned(4,8) ,
26264	 => std_logic_vector(to_unsigned(4,8) ,
26265	 => std_logic_vector(to_unsigned(3,8) ,
26266	 => std_logic_vector(to_unsigned(3,8) ,
26267	 => std_logic_vector(to_unsigned(1,8) ,
26268	 => std_logic_vector(to_unsigned(2,8) ,
26269	 => std_logic_vector(to_unsigned(18,8) ,
26270	 => std_logic_vector(to_unsigned(81,8) ,
26271	 => std_logic_vector(to_unsigned(142,8) ,
26272	 => std_logic_vector(to_unsigned(164,8) ,
26273	 => std_logic_vector(to_unsigned(144,8) ,
26274	 => std_logic_vector(to_unsigned(101,8) ,
26275	 => std_logic_vector(to_unsigned(49,8) ,
26276	 => std_logic_vector(to_unsigned(23,8) ,
26277	 => std_logic_vector(to_unsigned(10,8) ,
26278	 => std_logic_vector(to_unsigned(3,8) ,
26279	 => std_logic_vector(to_unsigned(1,8) ,
26280	 => std_logic_vector(to_unsigned(31,8) ,
26281	 => std_logic_vector(to_unsigned(142,8) ,
26282	 => std_logic_vector(to_unsigned(122,8) ,
26283	 => std_logic_vector(to_unsigned(107,8) ,
26284	 => std_logic_vector(to_unsigned(41,8) ,
26285	 => std_logic_vector(to_unsigned(5,8) ,
26286	 => std_logic_vector(to_unsigned(1,8) ,
26287	 => std_logic_vector(to_unsigned(1,8) ,
26288	 => std_logic_vector(to_unsigned(0,8) ,
26289	 => std_logic_vector(to_unsigned(25,8) ,
26290	 => std_logic_vector(to_unsigned(183,8) ,
26291	 => std_logic_vector(to_unsigned(177,8) ,
26292	 => std_logic_vector(to_unsigned(179,8) ,
26293	 => std_logic_vector(to_unsigned(175,8) ,
26294	 => std_logic_vector(to_unsigned(161,8) ,
26295	 => std_logic_vector(to_unsigned(173,8) ,
26296	 => std_logic_vector(to_unsigned(166,8) ,
26297	 => std_logic_vector(to_unsigned(43,8) ,
26298	 => std_logic_vector(to_unsigned(5,8) ,
26299	 => std_logic_vector(to_unsigned(16,8) ,
26300	 => std_logic_vector(to_unsigned(13,8) ,
26301	 => std_logic_vector(to_unsigned(11,8) ,
26302	 => std_logic_vector(to_unsigned(6,8) ,
26303	 => std_logic_vector(to_unsigned(6,8) ,
26304	 => std_logic_vector(to_unsigned(8,8) ,
26305	 => std_logic_vector(to_unsigned(7,8) ,
26306	 => std_logic_vector(to_unsigned(7,8) ,
26307	 => std_logic_vector(to_unsigned(7,8) ,
26308	 => std_logic_vector(to_unsigned(4,8) ,
26309	 => std_logic_vector(to_unsigned(3,8) ,
26310	 => std_logic_vector(to_unsigned(4,8) ,
26311	 => std_logic_vector(to_unsigned(4,8) ,
26312	 => std_logic_vector(to_unsigned(6,8) ,
26313	 => std_logic_vector(to_unsigned(6,8) ,
26314	 => std_logic_vector(to_unsigned(3,8) ,
26315	 => std_logic_vector(to_unsigned(2,8) ,
26316	 => std_logic_vector(to_unsigned(2,8) ,
26317	 => std_logic_vector(to_unsigned(8,8) ,
26318	 => std_logic_vector(to_unsigned(74,8) ,
26319	 => std_logic_vector(to_unsigned(156,8) ,
26320	 => std_logic_vector(to_unsigned(168,8) ,
26321	 => std_logic_vector(to_unsigned(130,8) ,
26322	 => std_logic_vector(to_unsigned(104,8) ,
26323	 => std_logic_vector(to_unsigned(119,8) ,
26324	 => std_logic_vector(to_unsigned(88,8) ,
26325	 => std_logic_vector(to_unsigned(19,8) ,
26326	 => std_logic_vector(to_unsigned(39,8) ,
26327	 => std_logic_vector(to_unsigned(192,8) ,
26328	 => std_logic_vector(to_unsigned(166,8) ,
26329	 => std_logic_vector(to_unsigned(130,8) ,
26330	 => std_logic_vector(to_unsigned(85,8) ,
26331	 => std_logic_vector(to_unsigned(121,8) ,
26332	 => std_logic_vector(to_unsigned(131,8) ,
26333	 => std_logic_vector(to_unsigned(144,8) ,
26334	 => std_logic_vector(to_unsigned(161,8) ,
26335	 => std_logic_vector(to_unsigned(161,8) ,
26336	 => std_logic_vector(to_unsigned(149,8) ,
26337	 => std_logic_vector(to_unsigned(121,8) ,
26338	 => std_logic_vector(to_unsigned(104,8) ,
26339	 => std_logic_vector(to_unsigned(118,8) ,
26340	 => std_logic_vector(to_unsigned(161,8) ,
26341	 => std_logic_vector(to_unsigned(128,8) ,
26342	 => std_logic_vector(to_unsigned(53,8) ,
26343	 => std_logic_vector(to_unsigned(99,8) ,
26344	 => std_logic_vector(to_unsigned(118,8) ,
26345	 => std_logic_vector(to_unsigned(85,8) ,
26346	 => std_logic_vector(to_unsigned(62,8) ,
26347	 => std_logic_vector(to_unsigned(44,8) ,
26348	 => std_logic_vector(to_unsigned(103,8) ,
26349	 => std_logic_vector(to_unsigned(43,8) ,
26350	 => std_logic_vector(to_unsigned(7,8) ,
26351	 => std_logic_vector(to_unsigned(23,8) ,
26352	 => std_logic_vector(to_unsigned(53,8) ,
26353	 => std_logic_vector(to_unsigned(24,8) ,
26354	 => std_logic_vector(to_unsigned(2,8) ,
26355	 => std_logic_vector(to_unsigned(0,8) ,
26356	 => std_logic_vector(to_unsigned(1,8) ,
26357	 => std_logic_vector(to_unsigned(0,8) ,
26358	 => std_logic_vector(to_unsigned(5,8) ,
26359	 => std_logic_vector(to_unsigned(29,8) ,
26360	 => std_logic_vector(to_unsigned(10,8) ,
26361	 => std_logic_vector(to_unsigned(0,8) ,
26362	 => std_logic_vector(to_unsigned(3,8) ,
26363	 => std_logic_vector(to_unsigned(11,8) ,
26364	 => std_logic_vector(to_unsigned(20,8) ,
26365	 => std_logic_vector(to_unsigned(9,8) ,
26366	 => std_logic_vector(to_unsigned(2,8) ,
26367	 => std_logic_vector(to_unsigned(2,8) ,
26368	 => std_logic_vector(to_unsigned(8,8) ,
26369	 => std_logic_vector(to_unsigned(24,8) ,
26370	 => std_logic_vector(to_unsigned(51,8) ,
26371	 => std_logic_vector(to_unsigned(121,8) ,
26372	 => std_logic_vector(to_unsigned(99,8) ,
26373	 => std_logic_vector(to_unsigned(81,8) ,
26374	 => std_logic_vector(to_unsigned(70,8) ,
26375	 => std_logic_vector(to_unsigned(60,8) ,
26376	 => std_logic_vector(to_unsigned(142,8) ,
26377	 => std_logic_vector(to_unsigned(122,8) ,
26378	 => std_logic_vector(to_unsigned(45,8) ,
26379	 => std_logic_vector(to_unsigned(19,8) ,
26380	 => std_logic_vector(to_unsigned(20,8) ,
26381	 => std_logic_vector(to_unsigned(18,8) ,
26382	 => std_logic_vector(to_unsigned(22,8) ,
26383	 => std_logic_vector(to_unsigned(12,8) ,
26384	 => std_logic_vector(to_unsigned(17,8) ,
26385	 => std_logic_vector(to_unsigned(17,8) ,
26386	 => std_logic_vector(to_unsigned(19,8) ,
26387	 => std_logic_vector(to_unsigned(18,8) ,
26388	 => std_logic_vector(to_unsigned(26,8) ,
26389	 => std_logic_vector(to_unsigned(35,8) ,
26390	 => std_logic_vector(to_unsigned(5,8) ,
26391	 => std_logic_vector(to_unsigned(7,8) ,
26392	 => std_logic_vector(to_unsigned(14,8) ,
26393	 => std_logic_vector(to_unsigned(10,8) ,
26394	 => std_logic_vector(to_unsigned(13,8) ,
26395	 => std_logic_vector(to_unsigned(17,8) ,
26396	 => std_logic_vector(to_unsigned(25,8) ,
26397	 => std_logic_vector(to_unsigned(32,8) ,
26398	 => std_logic_vector(to_unsigned(19,8) ,
26399	 => std_logic_vector(to_unsigned(30,8) ,
26400	 => std_logic_vector(to_unsigned(39,8) ,
26401	 => std_logic_vector(to_unsigned(46,8) ,
26402	 => std_logic_vector(to_unsigned(32,8) ,
26403	 => std_logic_vector(to_unsigned(17,8) ,
26404	 => std_logic_vector(to_unsigned(18,8) ,
26405	 => std_logic_vector(to_unsigned(48,8) ,
26406	 => std_logic_vector(to_unsigned(25,8) ,
26407	 => std_logic_vector(to_unsigned(3,8) ,
26408	 => std_logic_vector(to_unsigned(10,8) ,
26409	 => std_logic_vector(to_unsigned(30,8) ,
26410	 => std_logic_vector(to_unsigned(24,8) ,
26411	 => std_logic_vector(to_unsigned(22,8) ,
26412	 => std_logic_vector(to_unsigned(20,8) ,
26413	 => std_logic_vector(to_unsigned(14,8) ,
26414	 => std_logic_vector(to_unsigned(8,8) ,
26415	 => std_logic_vector(to_unsigned(14,8) ,
26416	 => std_logic_vector(to_unsigned(30,8) ,
26417	 => std_logic_vector(to_unsigned(31,8) ,
26418	 => std_logic_vector(to_unsigned(30,8) ,
26419	 => std_logic_vector(to_unsigned(37,8) ,
26420	 => std_logic_vector(to_unsigned(27,8) ,
26421	 => std_logic_vector(to_unsigned(16,8) ,
26422	 => std_logic_vector(to_unsigned(6,8) ,
26423	 => std_logic_vector(to_unsigned(2,8) ,
26424	 => std_logic_vector(to_unsigned(13,8) ,
26425	 => std_logic_vector(to_unsigned(23,8) ,
26426	 => std_logic_vector(to_unsigned(12,8) ,
26427	 => std_logic_vector(to_unsigned(48,8) ,
26428	 => std_logic_vector(to_unsigned(88,8) ,
26429	 => std_logic_vector(to_unsigned(65,8) ,
26430	 => std_logic_vector(to_unsigned(96,8) ,
26431	 => std_logic_vector(to_unsigned(119,8) ,
26432	 => std_logic_vector(to_unsigned(141,8) ,
26433	 => std_logic_vector(to_unsigned(131,8) ,
26434	 => std_logic_vector(to_unsigned(125,8) ,
26435	 => std_logic_vector(to_unsigned(118,8) ,
26436	 => std_logic_vector(to_unsigned(62,8) ,
26437	 => std_logic_vector(to_unsigned(6,8) ,
26438	 => std_logic_vector(to_unsigned(6,8) ,
26439	 => std_logic_vector(to_unsigned(7,8) ,
26440	 => std_logic_vector(to_unsigned(7,8) ,
26441	 => std_logic_vector(to_unsigned(21,8) ,
26442	 => std_logic_vector(to_unsigned(42,8) ,
26443	 => std_logic_vector(to_unsigned(21,8) ,
26444	 => std_logic_vector(to_unsigned(28,8) ,
26445	 => std_logic_vector(to_unsigned(142,8) ,
26446	 => std_logic_vector(to_unsigned(141,8) ,
26447	 => std_logic_vector(to_unsigned(138,8) ,
26448	 => std_logic_vector(to_unsigned(96,8) ,
26449	 => std_logic_vector(to_unsigned(79,8) ,
26450	 => std_logic_vector(to_unsigned(146,8) ,
26451	 => std_logic_vector(to_unsigned(149,8) ,
26452	 => std_logic_vector(to_unsigned(154,8) ,
26453	 => std_logic_vector(to_unsigned(147,8) ,
26454	 => std_logic_vector(to_unsigned(134,8) ,
26455	 => std_logic_vector(to_unsigned(134,8) ,
26456	 => std_logic_vector(to_unsigned(142,8) ,
26457	 => std_logic_vector(to_unsigned(139,8) ,
26458	 => std_logic_vector(to_unsigned(152,8) ,
26459	 => std_logic_vector(to_unsigned(87,8) ,
26460	 => std_logic_vector(to_unsigned(9,8) ,
26461	 => std_logic_vector(to_unsigned(9,8) ,
26462	 => std_logic_vector(to_unsigned(12,8) ,
26463	 => std_logic_vector(to_unsigned(7,8) ,
26464	 => std_logic_vector(to_unsigned(38,8) ,
26465	 => std_logic_vector(to_unsigned(116,8) ,
26466	 => std_logic_vector(to_unsigned(15,8) ,
26467	 => std_logic_vector(to_unsigned(9,8) ,
26468	 => std_logic_vector(to_unsigned(7,8) ,
26469	 => std_logic_vector(to_unsigned(4,8) ,
26470	 => std_logic_vector(to_unsigned(6,8) ,
26471	 => std_logic_vector(to_unsigned(8,8) ,
26472	 => std_logic_vector(to_unsigned(16,8) ,
26473	 => std_logic_vector(to_unsigned(20,8) ,
26474	 => std_logic_vector(to_unsigned(49,8) ,
26475	 => std_logic_vector(to_unsigned(159,8) ,
26476	 => std_logic_vector(to_unsigned(142,8) ,
26477	 => std_logic_vector(to_unsigned(31,8) ,
26478	 => std_logic_vector(to_unsigned(30,8) ,
26479	 => std_logic_vector(to_unsigned(65,8) ,
26480	 => std_logic_vector(to_unsigned(78,8) ,
26481	 => std_logic_vector(to_unsigned(125,8) ,
26482	 => std_logic_vector(to_unsigned(84,8) ,
26483	 => std_logic_vector(to_unsigned(10,8) ,
26484	 => std_logic_vector(to_unsigned(4,8) ,
26485	 => std_logic_vector(to_unsigned(3,8) ,
26486	 => std_logic_vector(to_unsigned(3,8) ,
26487	 => std_logic_vector(to_unsigned(4,8) ,
26488	 => std_logic_vector(to_unsigned(5,8) ,
26489	 => std_logic_vector(to_unsigned(7,8) ,
26490	 => std_logic_vector(to_unsigned(9,8) ,
26491	 => std_logic_vector(to_unsigned(6,8) ,
26492	 => std_logic_vector(to_unsigned(6,8) ,
26493	 => std_logic_vector(to_unsigned(9,8) ,
26494	 => std_logic_vector(to_unsigned(10,8) ,
26495	 => std_logic_vector(to_unsigned(18,8) ,
26496	 => std_logic_vector(to_unsigned(24,8) ,
26497	 => std_logic_vector(to_unsigned(9,8) ,
26498	 => std_logic_vector(to_unsigned(6,8) ,
26499	 => std_logic_vector(to_unsigned(23,8) ,
26500	 => std_logic_vector(to_unsigned(19,8) ,
26501	 => std_logic_vector(to_unsigned(7,8) ,
26502	 => std_logic_vector(to_unsigned(12,8) ,
26503	 => std_logic_vector(to_unsigned(68,8) ,
26504	 => std_logic_vector(to_unsigned(104,8) ,
26505	 => std_logic_vector(to_unsigned(91,8) ,
26506	 => std_logic_vector(to_unsigned(127,8) ,
26507	 => std_logic_vector(to_unsigned(159,8) ,
26508	 => std_logic_vector(to_unsigned(179,8) ,
26509	 => std_logic_vector(to_unsigned(125,8) ,
26510	 => std_logic_vector(to_unsigned(60,8) ,
26511	 => std_logic_vector(to_unsigned(80,8) ,
26512	 => std_logic_vector(to_unsigned(49,8) ,
26513	 => std_logic_vector(to_unsigned(36,8) ,
26514	 => std_logic_vector(to_unsigned(17,8) ,
26515	 => std_logic_vector(to_unsigned(1,8) ,
26516	 => std_logic_vector(to_unsigned(1,8) ,
26517	 => std_logic_vector(to_unsigned(17,8) ,
26518	 => std_logic_vector(to_unsigned(29,8) ,
26519	 => std_logic_vector(to_unsigned(19,8) ,
26520	 => std_logic_vector(to_unsigned(9,8) ,
26521	 => std_logic_vector(to_unsigned(7,8) ,
26522	 => std_logic_vector(to_unsigned(3,8) ,
26523	 => std_logic_vector(to_unsigned(12,8) ,
26524	 => std_logic_vector(to_unsigned(104,8) ,
26525	 => std_logic_vector(to_unsigned(35,8) ,
26526	 => std_logic_vector(to_unsigned(0,8) ,
26527	 => std_logic_vector(to_unsigned(45,8) ,
26528	 => std_logic_vector(to_unsigned(164,8) ,
26529	 => std_logic_vector(to_unsigned(46,8) ,
26530	 => std_logic_vector(to_unsigned(6,8) ,
26531	 => std_logic_vector(to_unsigned(44,8) ,
26532	 => std_logic_vector(to_unsigned(59,8) ,
26533	 => std_logic_vector(to_unsigned(70,8) ,
26534	 => std_logic_vector(to_unsigned(118,8) ,
26535	 => std_logic_vector(to_unsigned(142,8) ,
26536	 => std_logic_vector(to_unsigned(119,8) ,
26537	 => std_logic_vector(to_unsigned(72,8) ,
26538	 => std_logic_vector(to_unsigned(71,8) ,
26539	 => std_logic_vector(to_unsigned(99,8) ,
26540	 => std_logic_vector(to_unsigned(109,8) ,
26541	 => std_logic_vector(to_unsigned(109,8) ,
26542	 => std_logic_vector(to_unsigned(122,8) ,
26543	 => std_logic_vector(to_unsigned(109,8) ,
26544	 => std_logic_vector(to_unsigned(107,8) ,
26545	 => std_logic_vector(to_unsigned(107,8) ,
26546	 => std_logic_vector(to_unsigned(127,8) ,
26547	 => std_logic_vector(to_unsigned(138,8) ,
26548	 => std_logic_vector(to_unsigned(127,8) ,
26549	 => std_logic_vector(to_unsigned(118,8) ,
26550	 => std_logic_vector(to_unsigned(131,8) ,
26551	 => std_logic_vector(to_unsigned(138,8) ,
26552	 => std_logic_vector(to_unsigned(139,8) ,
26553	 => std_logic_vector(to_unsigned(136,8) ,
26554	 => std_logic_vector(to_unsigned(131,8) ,
26555	 => std_logic_vector(to_unsigned(144,8) ,
26556	 => std_logic_vector(to_unsigned(163,8) ,
26557	 => std_logic_vector(to_unsigned(166,8) ,
26558	 => std_logic_vector(to_unsigned(161,8) ,
26559	 => std_logic_vector(to_unsigned(134,8) ,
26560	 => std_logic_vector(to_unsigned(121,8) ,
26561	 => std_logic_vector(to_unsigned(166,8) ,
26562	 => std_logic_vector(to_unsigned(163,8) ,
26563	 => std_logic_vector(to_unsigned(161,8) ,
26564	 => std_logic_vector(to_unsigned(164,8) ,
26565	 => std_logic_vector(to_unsigned(164,8) ,
26566	 => std_logic_vector(to_unsigned(159,8) ,
26567	 => std_logic_vector(to_unsigned(65,8) ,
26568	 => std_logic_vector(to_unsigned(32,8) ,
26569	 => std_logic_vector(to_unsigned(28,8) ,
26570	 => std_logic_vector(to_unsigned(40,8) ,
26571	 => std_logic_vector(to_unsigned(44,8) ,
26572	 => std_logic_vector(to_unsigned(35,8) ,
26573	 => std_logic_vector(to_unsigned(12,8) ,
26574	 => std_logic_vector(to_unsigned(2,8) ,
26575	 => std_logic_vector(to_unsigned(6,8) ,
26576	 => std_logic_vector(to_unsigned(14,8) ,
26577	 => std_logic_vector(to_unsigned(5,8) ,
26578	 => std_logic_vector(to_unsigned(2,8) ,
26579	 => std_logic_vector(to_unsigned(1,8) ,
26580	 => std_logic_vector(to_unsigned(2,8) ,
26581	 => std_logic_vector(to_unsigned(4,8) ,
26582	 => std_logic_vector(to_unsigned(3,8) ,
26583	 => std_logic_vector(to_unsigned(2,8) ,
26584	 => std_logic_vector(to_unsigned(2,8) ,
26585	 => std_logic_vector(to_unsigned(1,8) ,
26586	 => std_logic_vector(to_unsigned(1,8) ,
26587	 => std_logic_vector(to_unsigned(1,8) ,
26588	 => std_logic_vector(to_unsigned(0,8) ,
26589	 => std_logic_vector(to_unsigned(1,8) ,
26590	 => std_logic_vector(to_unsigned(14,8) ,
26591	 => std_logic_vector(to_unsigned(72,8) ,
26592	 => std_logic_vector(to_unsigned(133,8) ,
26593	 => std_logic_vector(to_unsigned(146,8) ,
26594	 => std_logic_vector(to_unsigned(146,8) ,
26595	 => std_logic_vector(to_unsigned(152,8) ,
26596	 => std_logic_vector(to_unsigned(149,8) ,
26597	 => std_logic_vector(to_unsigned(121,8) ,
26598	 => std_logic_vector(to_unsigned(87,8) ,
26599	 => std_logic_vector(to_unsigned(47,8) ,
26600	 => std_logic_vector(to_unsigned(84,8) ,
26601	 => std_logic_vector(to_unsigned(122,8) ,
26602	 => std_logic_vector(to_unsigned(104,8) ,
26603	 => std_logic_vector(to_unsigned(69,8) ,
26604	 => std_logic_vector(to_unsigned(15,8) ,
26605	 => std_logic_vector(to_unsigned(2,8) ,
26606	 => std_logic_vector(to_unsigned(1,8) ,
26607	 => std_logic_vector(to_unsigned(1,8) ,
26608	 => std_logic_vector(to_unsigned(0,8) ,
26609	 => std_logic_vector(to_unsigned(8,8) ,
26610	 => std_logic_vector(to_unsigned(34,8) ,
26611	 => std_logic_vector(to_unsigned(32,8) ,
26612	 => std_logic_vector(to_unsigned(65,8) ,
26613	 => std_logic_vector(to_unsigned(125,8) ,
26614	 => std_logic_vector(to_unsigned(142,8) ,
26615	 => std_logic_vector(to_unsigned(146,8) ,
26616	 => std_logic_vector(to_unsigned(168,8) ,
26617	 => std_logic_vector(to_unsigned(59,8) ,
26618	 => std_logic_vector(to_unsigned(4,8) ,
26619	 => std_logic_vector(to_unsigned(16,8) ,
26620	 => std_logic_vector(to_unsigned(20,8) ,
26621	 => std_logic_vector(to_unsigned(14,8) ,
26622	 => std_logic_vector(to_unsigned(10,8) ,
26623	 => std_logic_vector(to_unsigned(5,8) ,
26624	 => std_logic_vector(to_unsigned(5,8) ,
26625	 => std_logic_vector(to_unsigned(8,8) ,
26626	 => std_logic_vector(to_unsigned(8,8) ,
26627	 => std_logic_vector(to_unsigned(5,8) ,
26628	 => std_logic_vector(to_unsigned(4,8) ,
26629	 => std_logic_vector(to_unsigned(5,8) ,
26630	 => std_logic_vector(to_unsigned(4,8) ,
26631	 => std_logic_vector(to_unsigned(5,8) ,
26632	 => std_logic_vector(to_unsigned(7,8) ,
26633	 => std_logic_vector(to_unsigned(4,8) ,
26634	 => std_logic_vector(to_unsigned(3,8) ,
26635	 => std_logic_vector(to_unsigned(4,8) ,
26636	 => std_logic_vector(to_unsigned(2,8) ,
26637	 => std_logic_vector(to_unsigned(2,8) ,
26638	 => std_logic_vector(to_unsigned(7,8) ,
26639	 => std_logic_vector(to_unsigned(96,8) ,
26640	 => std_logic_vector(to_unsigned(144,8) ,
26641	 => std_logic_vector(to_unsigned(111,8) ,
26642	 => std_logic_vector(to_unsigned(115,8) ,
26643	 => std_logic_vector(to_unsigned(104,8) ,
26644	 => std_logic_vector(to_unsigned(100,8) ,
26645	 => std_logic_vector(to_unsigned(71,8) ,
26646	 => std_logic_vector(to_unsigned(36,8) ,
26647	 => std_logic_vector(to_unsigned(82,8) ,
26648	 => std_logic_vector(to_unsigned(170,8) ,
26649	 => std_logic_vector(to_unsigned(122,8) ,
26650	 => std_logic_vector(to_unsigned(84,8) ,
26651	 => std_logic_vector(to_unsigned(108,8) ,
26652	 => std_logic_vector(to_unsigned(138,8) ,
26653	 => std_logic_vector(to_unsigned(154,8) ,
26654	 => std_logic_vector(to_unsigned(142,8) ,
26655	 => std_logic_vector(to_unsigned(136,8) ,
26656	 => std_logic_vector(to_unsigned(147,8) ,
26657	 => std_logic_vector(to_unsigned(127,8) ,
26658	 => std_logic_vector(to_unsigned(127,8) ,
26659	 => std_logic_vector(to_unsigned(133,8) ,
26660	 => std_logic_vector(to_unsigned(159,8) ,
26661	 => std_logic_vector(to_unsigned(67,8) ,
26662	 => std_logic_vector(to_unsigned(35,8) ,
26663	 => std_logic_vector(to_unsigned(130,8) ,
26664	 => std_logic_vector(to_unsigned(108,8) ,
26665	 => std_logic_vector(to_unsigned(88,8) ,
26666	 => std_logic_vector(to_unsigned(41,8) ,
26667	 => std_logic_vector(to_unsigned(16,8) ,
26668	 => std_logic_vector(to_unsigned(118,8) ,
26669	 => std_logic_vector(to_unsigned(62,8) ,
26670	 => std_logic_vector(to_unsigned(9,8) ,
26671	 => std_logic_vector(to_unsigned(18,8) ,
26672	 => std_logic_vector(to_unsigned(57,8) ,
26673	 => std_logic_vector(to_unsigned(32,8) ,
26674	 => std_logic_vector(to_unsigned(2,8) ,
26675	 => std_logic_vector(to_unsigned(1,8) ,
26676	 => std_logic_vector(to_unsigned(1,8) ,
26677	 => std_logic_vector(to_unsigned(1,8) ,
26678	 => std_logic_vector(to_unsigned(0,8) ,
26679	 => std_logic_vector(to_unsigned(5,8) ,
26680	 => std_logic_vector(to_unsigned(16,8) ,
26681	 => std_logic_vector(to_unsigned(1,8) ,
26682	 => std_logic_vector(to_unsigned(1,8) ,
26683	 => std_logic_vector(to_unsigned(2,8) ,
26684	 => std_logic_vector(to_unsigned(8,8) ,
26685	 => std_logic_vector(to_unsigned(5,8) ,
26686	 => std_logic_vector(to_unsigned(3,8) ,
26687	 => std_logic_vector(to_unsigned(2,8) ,
26688	 => std_logic_vector(to_unsigned(10,8) ,
26689	 => std_logic_vector(to_unsigned(59,8) ,
26690	 => std_logic_vector(to_unsigned(73,8) ,
26691	 => std_logic_vector(to_unsigned(104,8) ,
26692	 => std_logic_vector(to_unsigned(103,8) ,
26693	 => std_logic_vector(to_unsigned(95,8) ,
26694	 => std_logic_vector(to_unsigned(63,8) ,
26695	 => std_logic_vector(to_unsigned(45,8) ,
26696	 => std_logic_vector(to_unsigned(119,8) ,
26697	 => std_logic_vector(to_unsigned(121,8) ,
26698	 => std_logic_vector(to_unsigned(45,8) ,
26699	 => std_logic_vector(to_unsigned(16,8) ,
26700	 => std_logic_vector(to_unsigned(12,8) ,
26701	 => std_logic_vector(to_unsigned(10,8) ,
26702	 => std_logic_vector(to_unsigned(13,8) ,
26703	 => std_logic_vector(to_unsigned(18,8) ,
26704	 => std_logic_vector(to_unsigned(32,8) ,
26705	 => std_logic_vector(to_unsigned(29,8) ,
26706	 => std_logic_vector(to_unsigned(31,8) ,
26707	 => std_logic_vector(to_unsigned(46,8) ,
26708	 => std_logic_vector(to_unsigned(25,8) ,
26709	 => std_logic_vector(to_unsigned(8,8) ,
26710	 => std_logic_vector(to_unsigned(6,8) ,
26711	 => std_logic_vector(to_unsigned(14,8) ,
26712	 => std_logic_vector(to_unsigned(14,8) ,
26713	 => std_logic_vector(to_unsigned(17,8) ,
26714	 => std_logic_vector(to_unsigned(21,8) ,
26715	 => std_logic_vector(to_unsigned(17,8) ,
26716	 => std_logic_vector(to_unsigned(15,8) ,
26717	 => std_logic_vector(to_unsigned(18,8) ,
26718	 => std_logic_vector(to_unsigned(17,8) ,
26719	 => std_logic_vector(to_unsigned(34,8) ,
26720	 => std_logic_vector(to_unsigned(37,8) ,
26721	 => std_logic_vector(to_unsigned(44,8) ,
26722	 => std_logic_vector(to_unsigned(27,8) ,
26723	 => std_logic_vector(to_unsigned(27,8) ,
26724	 => std_logic_vector(to_unsigned(18,8) ,
26725	 => std_logic_vector(to_unsigned(49,8) ,
26726	 => std_logic_vector(to_unsigned(54,8) ,
26727	 => std_logic_vector(to_unsigned(14,8) ,
26728	 => std_logic_vector(to_unsigned(4,8) ,
26729	 => std_logic_vector(to_unsigned(21,8) ,
26730	 => std_logic_vector(to_unsigned(22,8) ,
26731	 => std_logic_vector(to_unsigned(24,8) ,
26732	 => std_logic_vector(to_unsigned(25,8) ,
26733	 => std_logic_vector(to_unsigned(17,8) ,
26734	 => std_logic_vector(to_unsigned(7,8) ,
26735	 => std_logic_vector(to_unsigned(10,8) ,
26736	 => std_logic_vector(to_unsigned(29,8) ,
26737	 => std_logic_vector(to_unsigned(39,8) ,
26738	 => std_logic_vector(to_unsigned(29,8) ,
26739	 => std_logic_vector(to_unsigned(26,8) ,
26740	 => std_logic_vector(to_unsigned(20,8) ,
26741	 => std_logic_vector(to_unsigned(14,8) ,
26742	 => std_logic_vector(to_unsigned(5,8) ,
26743	 => std_logic_vector(to_unsigned(1,8) ,
26744	 => std_logic_vector(to_unsigned(12,8) ,
26745	 => std_logic_vector(to_unsigned(17,8) ,
26746	 => std_logic_vector(to_unsigned(9,8) ,
26747	 => std_logic_vector(to_unsigned(56,8) ,
26748	 => std_logic_vector(to_unsigned(92,8) ,
26749	 => std_logic_vector(to_unsigned(48,8) ,
26750	 => std_logic_vector(to_unsigned(74,8) ,
26751	 => std_logic_vector(to_unsigned(100,8) ,
26752	 => std_logic_vector(to_unsigned(131,8) ,
26753	 => std_logic_vector(to_unsigned(134,8) ,
26754	 => std_logic_vector(to_unsigned(108,8) ,
26755	 => std_logic_vector(to_unsigned(112,8) ,
26756	 => std_logic_vector(to_unsigned(146,8) ,
26757	 => std_logic_vector(to_unsigned(41,8) ,
26758	 => std_logic_vector(to_unsigned(3,8) ,
26759	 => std_logic_vector(to_unsigned(5,8) ,
26760	 => std_logic_vector(to_unsigned(2,8) ,
26761	 => std_logic_vector(to_unsigned(4,8) ,
26762	 => std_logic_vector(to_unsigned(15,8) ,
26763	 => std_logic_vector(to_unsigned(30,8) ,
26764	 => std_logic_vector(to_unsigned(63,8) ,
26765	 => std_logic_vector(to_unsigned(146,8) ,
26766	 => std_logic_vector(to_unsigned(141,8) ,
26767	 => std_logic_vector(to_unsigned(163,8) ,
26768	 => std_logic_vector(to_unsigned(37,8) ,
26769	 => std_logic_vector(to_unsigned(24,8) ,
26770	 => std_logic_vector(to_unsigned(146,8) ,
26771	 => std_logic_vector(to_unsigned(146,8) ,
26772	 => std_logic_vector(to_unsigned(157,8) ,
26773	 => std_logic_vector(to_unsigned(154,8) ,
26774	 => std_logic_vector(to_unsigned(142,8) ,
26775	 => std_logic_vector(to_unsigned(136,8) ,
26776	 => std_logic_vector(to_unsigned(139,8) ,
26777	 => std_logic_vector(to_unsigned(141,8) ,
26778	 => std_logic_vector(to_unsigned(151,8) ,
26779	 => std_logic_vector(to_unsigned(56,8) ,
26780	 => std_logic_vector(to_unsigned(6,8) ,
26781	 => std_logic_vector(to_unsigned(12,8) ,
26782	 => std_logic_vector(to_unsigned(11,8) ,
26783	 => std_logic_vector(to_unsigned(9,8) ,
26784	 => std_logic_vector(to_unsigned(73,8) ,
26785	 => std_logic_vector(to_unsigned(138,8) ,
26786	 => std_logic_vector(to_unsigned(16,8) ,
26787	 => std_logic_vector(to_unsigned(7,8) ,
26788	 => std_logic_vector(to_unsigned(10,8) ,
26789	 => std_logic_vector(to_unsigned(8,8) ,
26790	 => std_logic_vector(to_unsigned(12,8) ,
26791	 => std_logic_vector(to_unsigned(13,8) ,
26792	 => std_logic_vector(to_unsigned(24,8) ,
26793	 => std_logic_vector(to_unsigned(40,8) ,
26794	 => std_logic_vector(to_unsigned(108,8) ,
26795	 => std_logic_vector(to_unsigned(179,8) ,
26796	 => std_logic_vector(to_unsigned(85,8) ,
26797	 => std_logic_vector(to_unsigned(29,8) ,
26798	 => std_logic_vector(to_unsigned(41,8) ,
26799	 => std_logic_vector(to_unsigned(40,8) ,
26800	 => std_logic_vector(to_unsigned(61,8) ,
26801	 => std_logic_vector(to_unsigned(61,8) ,
26802	 => std_logic_vector(to_unsigned(11,8) ,
26803	 => std_logic_vector(to_unsigned(3,8) ,
26804	 => std_logic_vector(to_unsigned(7,8) ,
26805	 => std_logic_vector(to_unsigned(5,8) ,
26806	 => std_logic_vector(to_unsigned(2,8) ,
26807	 => std_logic_vector(to_unsigned(4,8) ,
26808	 => std_logic_vector(to_unsigned(9,8) ,
26809	 => std_logic_vector(to_unsigned(7,8) ,
26810	 => std_logic_vector(to_unsigned(3,8) ,
26811	 => std_logic_vector(to_unsigned(3,8) ,
26812	 => std_logic_vector(to_unsigned(7,8) ,
26813	 => std_logic_vector(to_unsigned(12,8) ,
26814	 => std_logic_vector(to_unsigned(19,8) ,
26815	 => std_logic_vector(to_unsigned(27,8) ,
26816	 => std_logic_vector(to_unsigned(15,8) ,
26817	 => std_logic_vector(to_unsigned(8,8) ,
26818	 => std_logic_vector(to_unsigned(7,8) ,
26819	 => std_logic_vector(to_unsigned(21,8) ,
26820	 => std_logic_vector(to_unsigned(22,8) ,
26821	 => std_logic_vector(to_unsigned(5,8) ,
26822	 => std_logic_vector(to_unsigned(11,8) ,
26823	 => std_logic_vector(to_unsigned(51,8) ,
26824	 => std_logic_vector(to_unsigned(79,8) ,
26825	 => std_logic_vector(to_unsigned(82,8) ,
26826	 => std_logic_vector(to_unsigned(95,8) ,
26827	 => std_logic_vector(to_unsigned(107,8) ,
26828	 => std_logic_vector(to_unsigned(141,8) ,
26829	 => std_logic_vector(to_unsigned(104,8) ,
26830	 => std_logic_vector(to_unsigned(55,8) ,
26831	 => std_logic_vector(to_unsigned(87,8) ,
26832	 => std_logic_vector(to_unsigned(48,8) ,
26833	 => std_logic_vector(to_unsigned(81,8) ,
26834	 => std_logic_vector(to_unsigned(71,8) ,
26835	 => std_logic_vector(to_unsigned(14,8) ,
26836	 => std_logic_vector(to_unsigned(36,8) ,
26837	 => std_logic_vector(to_unsigned(84,8) ,
26838	 => std_logic_vector(to_unsigned(107,8) ,
26839	 => std_logic_vector(to_unsigned(78,8) ,
26840	 => std_logic_vector(to_unsigned(35,8) ,
26841	 => std_logic_vector(to_unsigned(21,8) ,
26842	 => std_logic_vector(to_unsigned(10,8) ,
26843	 => std_logic_vector(to_unsigned(6,8) ,
26844	 => std_logic_vector(to_unsigned(65,8) ,
26845	 => std_logic_vector(to_unsigned(69,8) ,
26846	 => std_logic_vector(to_unsigned(18,8) ,
26847	 => std_logic_vector(to_unsigned(16,8) ,
26848	 => std_logic_vector(to_unsigned(49,8) ,
26849	 => std_logic_vector(to_unsigned(54,8) ,
26850	 => std_logic_vector(to_unsigned(10,8) ,
26851	 => std_logic_vector(to_unsigned(40,8) ,
26852	 => std_logic_vector(to_unsigned(59,8) ,
26853	 => std_logic_vector(to_unsigned(82,8) ,
26854	 => std_logic_vector(to_unsigned(100,8) ,
26855	 => std_logic_vector(to_unsigned(78,8) ,
26856	 => std_logic_vector(to_unsigned(105,8) ,
26857	 => std_logic_vector(to_unsigned(104,8) ,
26858	 => std_logic_vector(to_unsigned(62,8) ,
26859	 => std_logic_vector(to_unsigned(66,8) ,
26860	 => std_logic_vector(to_unsigned(124,8) ,
26861	 => std_logic_vector(to_unsigned(142,8) ,
26862	 => std_logic_vector(to_unsigned(133,8) ,
26863	 => std_logic_vector(to_unsigned(116,8) ,
26864	 => std_logic_vector(to_unsigned(115,8) ,
26865	 => std_logic_vector(to_unsigned(121,8) ,
26866	 => std_logic_vector(to_unsigned(131,8) ,
26867	 => std_logic_vector(to_unsigned(139,8) ,
26868	 => std_logic_vector(to_unsigned(136,8) ,
26869	 => std_logic_vector(to_unsigned(141,8) ,
26870	 => std_logic_vector(to_unsigned(136,8) ,
26871	 => std_logic_vector(to_unsigned(142,8) ,
26872	 => std_logic_vector(to_unsigned(151,8) ,
26873	 => std_logic_vector(to_unsigned(152,8) ,
26874	 => std_logic_vector(to_unsigned(138,8) ,
26875	 => std_logic_vector(to_unsigned(134,8) ,
26876	 => std_logic_vector(to_unsigned(156,8) ,
26877	 => std_logic_vector(to_unsigned(168,8) ,
26878	 => std_logic_vector(to_unsigned(166,8) ,
26879	 => std_logic_vector(to_unsigned(151,8) ,
26880	 => std_logic_vector(to_unsigned(139,8) ,
26881	 => std_logic_vector(to_unsigned(163,8) ,
26882	 => std_logic_vector(to_unsigned(164,8) ,
26883	 => std_logic_vector(to_unsigned(159,8) ,
26884	 => std_logic_vector(to_unsigned(159,8) ,
26885	 => std_logic_vector(to_unsigned(159,8) ,
26886	 => std_logic_vector(to_unsigned(170,8) ,
26887	 => std_logic_vector(to_unsigned(111,8) ,
26888	 => std_logic_vector(to_unsigned(22,8) ,
26889	 => std_logic_vector(to_unsigned(5,8) ,
26890	 => std_logic_vector(to_unsigned(22,8) ,
26891	 => std_logic_vector(to_unsigned(10,8) ,
26892	 => std_logic_vector(to_unsigned(0,8) ,
26893	 => std_logic_vector(to_unsigned(0,8) ,
26894	 => std_logic_vector(to_unsigned(2,8) ,
26895	 => std_logic_vector(to_unsigned(4,8) ,
26896	 => std_logic_vector(to_unsigned(4,8) ,
26897	 => std_logic_vector(to_unsigned(2,8) ,
26898	 => std_logic_vector(to_unsigned(1,8) ,
26899	 => std_logic_vector(to_unsigned(1,8) ,
26900	 => std_logic_vector(to_unsigned(2,8) ,
26901	 => std_logic_vector(to_unsigned(2,8) ,
26902	 => std_logic_vector(to_unsigned(1,8) ,
26903	 => std_logic_vector(to_unsigned(1,8) ,
26904	 => std_logic_vector(to_unsigned(1,8) ,
26905	 => std_logic_vector(to_unsigned(0,8) ,
26906	 => std_logic_vector(to_unsigned(0,8) ,
26907	 => std_logic_vector(to_unsigned(0,8) ,
26908	 => std_logic_vector(to_unsigned(0,8) ,
26909	 => std_logic_vector(to_unsigned(0,8) ,
26910	 => std_logic_vector(to_unsigned(0,8) ,
26911	 => std_logic_vector(to_unsigned(7,8) ,
26912	 => std_logic_vector(to_unsigned(57,8) ,
26913	 => std_logic_vector(to_unsigned(116,8) ,
26914	 => std_logic_vector(to_unsigned(134,8) ,
26915	 => std_logic_vector(to_unsigned(138,8) ,
26916	 => std_logic_vector(to_unsigned(142,8) ,
26917	 => std_logic_vector(to_unsigned(151,8) ,
26918	 => std_logic_vector(to_unsigned(161,8) ,
26919	 => std_logic_vector(to_unsigned(149,8) ,
26920	 => std_logic_vector(to_unsigned(124,8) ,
26921	 => std_logic_vector(to_unsigned(108,8) ,
26922	 => std_logic_vector(to_unsigned(91,8) ,
26923	 => std_logic_vector(to_unsigned(46,8) ,
26924	 => std_logic_vector(to_unsigned(9,8) ,
26925	 => std_logic_vector(to_unsigned(1,8) ,
26926	 => std_logic_vector(to_unsigned(1,8) ,
26927	 => std_logic_vector(to_unsigned(1,8) ,
26928	 => std_logic_vector(to_unsigned(0,8) ,
26929	 => std_logic_vector(to_unsigned(1,8) ,
26930	 => std_logic_vector(to_unsigned(0,8) ,
26931	 => std_logic_vector(to_unsigned(1,8) ,
26932	 => std_logic_vector(to_unsigned(27,8) ,
26933	 => std_logic_vector(to_unsigned(93,8) ,
26934	 => std_logic_vector(to_unsigned(104,8) ,
26935	 => std_logic_vector(to_unsigned(93,8) ,
26936	 => std_logic_vector(to_unsigned(108,8) ,
26937	 => std_logic_vector(to_unsigned(42,8) ,
26938	 => std_logic_vector(to_unsigned(6,8) ,
26939	 => std_logic_vector(to_unsigned(12,8) ,
26940	 => std_logic_vector(to_unsigned(21,8) ,
26941	 => std_logic_vector(to_unsigned(15,8) ,
26942	 => std_logic_vector(to_unsigned(13,8) ,
26943	 => std_logic_vector(to_unsigned(8,8) ,
26944	 => std_logic_vector(to_unsigned(5,8) ,
26945	 => std_logic_vector(to_unsigned(6,8) ,
26946	 => std_logic_vector(to_unsigned(8,8) ,
26947	 => std_logic_vector(to_unsigned(5,8) ,
26948	 => std_logic_vector(to_unsigned(6,8) ,
26949	 => std_logic_vector(to_unsigned(9,8) ,
26950	 => std_logic_vector(to_unsigned(8,8) ,
26951	 => std_logic_vector(to_unsigned(8,8) ,
26952	 => std_logic_vector(to_unsigned(6,8) ,
26953	 => std_logic_vector(to_unsigned(3,8) ,
26954	 => std_logic_vector(to_unsigned(6,8) ,
26955	 => std_logic_vector(to_unsigned(6,8) ,
26956	 => std_logic_vector(to_unsigned(3,8) ,
26957	 => std_logic_vector(to_unsigned(4,8) ,
26958	 => std_logic_vector(to_unsigned(2,8) ,
26959	 => std_logic_vector(to_unsigned(10,8) ,
26960	 => std_logic_vector(to_unsigned(82,8) ,
26961	 => std_logic_vector(to_unsigned(112,8) ,
26962	 => std_logic_vector(to_unsigned(84,8) ,
26963	 => std_logic_vector(to_unsigned(72,8) ,
26964	 => std_logic_vector(to_unsigned(73,8) ,
26965	 => std_logic_vector(to_unsigned(38,8) ,
26966	 => std_logic_vector(to_unsigned(18,8) ,
26967	 => std_logic_vector(to_unsigned(8,8) ,
26968	 => std_logic_vector(to_unsigned(60,8) ,
26969	 => std_logic_vector(to_unsigned(92,8) ,
26970	 => std_logic_vector(to_unsigned(39,8) ,
26971	 => std_logic_vector(to_unsigned(72,8) ,
26972	 => std_logic_vector(to_unsigned(127,8) ,
26973	 => std_logic_vector(to_unsigned(141,8) ,
26974	 => std_logic_vector(to_unsigned(152,8) ,
26975	 => std_logic_vector(to_unsigned(144,8) ,
26976	 => std_logic_vector(to_unsigned(156,8) ,
26977	 => std_logic_vector(to_unsigned(147,8) ,
26978	 => std_logic_vector(to_unsigned(149,8) ,
26979	 => std_logic_vector(to_unsigned(152,8) ,
26980	 => std_logic_vector(to_unsigned(144,8) ,
26981	 => std_logic_vector(to_unsigned(16,8) ,
26982	 => std_logic_vector(to_unsigned(17,8) ,
26983	 => std_logic_vector(to_unsigned(124,8) ,
26984	 => std_logic_vector(to_unsigned(90,8) ,
26985	 => std_logic_vector(to_unsigned(79,8) ,
26986	 => std_logic_vector(to_unsigned(47,8) ,
26987	 => std_logic_vector(to_unsigned(25,8) ,
26988	 => std_logic_vector(to_unsigned(95,8) ,
26989	 => std_logic_vector(to_unsigned(115,8) ,
26990	 => std_logic_vector(to_unsigned(37,8) ,
26991	 => std_logic_vector(to_unsigned(10,8) ,
26992	 => std_logic_vector(to_unsigned(20,8) ,
26993	 => std_logic_vector(to_unsigned(18,8) ,
26994	 => std_logic_vector(to_unsigned(2,8) ,
26995	 => std_logic_vector(to_unsigned(1,8) ,
26996	 => std_logic_vector(to_unsigned(1,8) ,
26997	 => std_logic_vector(to_unsigned(1,8) ,
26998	 => std_logic_vector(to_unsigned(1,8) ,
26999	 => std_logic_vector(to_unsigned(2,8) ,
27000	 => std_logic_vector(to_unsigned(5,8) ,
27001	 => std_logic_vector(to_unsigned(1,8) ,
27002	 => std_logic_vector(to_unsigned(0,8) ,
27003	 => std_logic_vector(to_unsigned(2,8) ,
27004	 => std_logic_vector(to_unsigned(3,8) ,
27005	 => std_logic_vector(to_unsigned(2,8) ,
27006	 => std_logic_vector(to_unsigned(2,8) ,
27007	 => std_logic_vector(to_unsigned(2,8) ,
27008	 => std_logic_vector(to_unsigned(12,8) ,
27009	 => std_logic_vector(to_unsigned(78,8) ,
27010	 => std_logic_vector(to_unsigned(93,8) ,
27011	 => std_logic_vector(to_unsigned(78,8) ,
27012	 => std_logic_vector(to_unsigned(85,8) ,
27013	 => std_logic_vector(to_unsigned(93,8) ,
27014	 => std_logic_vector(to_unsigned(63,8) ,
27015	 => std_logic_vector(to_unsigned(45,8) ,
27016	 => std_logic_vector(to_unsigned(103,8) ,
27017	 => std_logic_vector(to_unsigned(108,8) ,
27018	 => std_logic_vector(to_unsigned(48,8) ,
27019	 => std_logic_vector(to_unsigned(18,8) ,
27020	 => std_logic_vector(to_unsigned(10,8) ,
27021	 => std_logic_vector(to_unsigned(6,8) ,
27022	 => std_logic_vector(to_unsigned(6,8) ,
27023	 => std_logic_vector(to_unsigned(15,8) ,
27024	 => std_logic_vector(to_unsigned(24,8) ,
27025	 => std_logic_vector(to_unsigned(27,8) ,
27026	 => std_logic_vector(to_unsigned(32,8) ,
27027	 => std_logic_vector(to_unsigned(27,8) ,
27028	 => std_logic_vector(to_unsigned(11,8) ,
27029	 => std_logic_vector(to_unsigned(15,8) ,
27030	 => std_logic_vector(to_unsigned(20,8) ,
27031	 => std_logic_vector(to_unsigned(13,8) ,
27032	 => std_logic_vector(to_unsigned(9,8) ,
27033	 => std_logic_vector(to_unsigned(12,8) ,
27034	 => std_logic_vector(to_unsigned(21,8) ,
27035	 => std_logic_vector(to_unsigned(12,8) ,
27036	 => std_logic_vector(to_unsigned(10,8) ,
27037	 => std_logic_vector(to_unsigned(9,8) ,
27038	 => std_logic_vector(to_unsigned(16,8) ,
27039	 => std_logic_vector(to_unsigned(29,8) ,
27040	 => std_logic_vector(to_unsigned(36,8) ,
27041	 => std_logic_vector(to_unsigned(37,8) ,
27042	 => std_logic_vector(to_unsigned(25,8) ,
27043	 => std_logic_vector(to_unsigned(35,8) ,
27044	 => std_logic_vector(to_unsigned(15,8) ,
27045	 => std_logic_vector(to_unsigned(45,8) ,
27046	 => std_logic_vector(to_unsigned(67,8) ,
27047	 => std_logic_vector(to_unsigned(35,8) ,
27048	 => std_logic_vector(to_unsigned(4,8) ,
27049	 => std_logic_vector(to_unsigned(10,8) ,
27050	 => std_logic_vector(to_unsigned(23,8) ,
27051	 => std_logic_vector(to_unsigned(25,8) ,
27052	 => std_logic_vector(to_unsigned(24,8) ,
27053	 => std_logic_vector(to_unsigned(17,8) ,
27054	 => std_logic_vector(to_unsigned(10,8) ,
27055	 => std_logic_vector(to_unsigned(9,8) ,
27056	 => std_logic_vector(to_unsigned(17,8) ,
27057	 => std_logic_vector(to_unsigned(29,8) ,
27058	 => std_logic_vector(to_unsigned(27,8) ,
27059	 => std_logic_vector(to_unsigned(24,8) ,
27060	 => std_logic_vector(to_unsigned(17,8) ,
27061	 => std_logic_vector(to_unsigned(10,8) ,
27062	 => std_logic_vector(to_unsigned(4,8) ,
27063	 => std_logic_vector(to_unsigned(1,8) ,
27064	 => std_logic_vector(to_unsigned(6,8) ,
27065	 => std_logic_vector(to_unsigned(13,8) ,
27066	 => std_logic_vector(to_unsigned(9,8) ,
27067	 => std_logic_vector(to_unsigned(64,8) ,
27068	 => std_logic_vector(to_unsigned(128,8) ,
27069	 => std_logic_vector(to_unsigned(84,8) ,
27070	 => std_logic_vector(to_unsigned(87,8) ,
27071	 => std_logic_vector(to_unsigned(99,8) ,
27072	 => std_logic_vector(to_unsigned(131,8) ,
27073	 => std_logic_vector(to_unsigned(131,8) ,
27074	 => std_logic_vector(to_unsigned(86,8) ,
27075	 => std_logic_vector(to_unsigned(85,8) ,
27076	 => std_logic_vector(to_unsigned(154,8) ,
27077	 => std_logic_vector(to_unsigned(124,8) ,
27078	 => std_logic_vector(to_unsigned(8,8) ,
27079	 => std_logic_vector(to_unsigned(2,8) ,
27080	 => std_logic_vector(to_unsigned(3,8) ,
27081	 => std_logic_vector(to_unsigned(3,8) ,
27082	 => std_logic_vector(to_unsigned(30,8) ,
27083	 => std_logic_vector(to_unsigned(97,8) ,
27084	 => std_logic_vector(to_unsigned(134,8) ,
27085	 => std_logic_vector(to_unsigned(147,8) ,
27086	 => std_logic_vector(to_unsigned(141,8) ,
27087	 => std_logic_vector(to_unsigned(88,8) ,
27088	 => std_logic_vector(to_unsigned(42,8) ,
27089	 => std_logic_vector(to_unsigned(92,8) ,
27090	 => std_logic_vector(to_unsigned(134,8) ,
27091	 => std_logic_vector(to_unsigned(142,8) ,
27092	 => std_logic_vector(to_unsigned(157,8) ,
27093	 => std_logic_vector(to_unsigned(149,8) ,
27094	 => std_logic_vector(to_unsigned(141,8) ,
27095	 => std_logic_vector(to_unsigned(134,8) ,
27096	 => std_logic_vector(to_unsigned(133,8) ,
27097	 => std_logic_vector(to_unsigned(136,8) ,
27098	 => std_logic_vector(to_unsigned(149,8) ,
27099	 => std_logic_vector(to_unsigned(45,8) ,
27100	 => std_logic_vector(to_unsigned(4,8) ,
27101	 => std_logic_vector(to_unsigned(8,8) ,
27102	 => std_logic_vector(to_unsigned(7,8) ,
27103	 => std_logic_vector(to_unsigned(12,8) ,
27104	 => std_logic_vector(to_unsigned(100,8) ,
27105	 => std_logic_vector(to_unsigned(146,8) ,
27106	 => std_logic_vector(to_unsigned(22,8) ,
27107	 => std_logic_vector(to_unsigned(8,8) ,
27108	 => std_logic_vector(to_unsigned(14,8) ,
27109	 => std_logic_vector(to_unsigned(13,8) ,
27110	 => std_logic_vector(to_unsigned(19,8) ,
27111	 => std_logic_vector(to_unsigned(30,8) ,
27112	 => std_logic_vector(to_unsigned(20,8) ,
27113	 => std_logic_vector(to_unsigned(50,8) ,
27114	 => std_logic_vector(to_unsigned(170,8) ,
27115	 => std_logic_vector(to_unsigned(151,8) ,
27116	 => std_logic_vector(to_unsigned(47,8) ,
27117	 => std_logic_vector(to_unsigned(34,8) ,
27118	 => std_logic_vector(to_unsigned(46,8) ,
27119	 => std_logic_vector(to_unsigned(38,8) ,
27120	 => std_logic_vector(to_unsigned(20,8) ,
27121	 => std_logic_vector(to_unsigned(11,8) ,
27122	 => std_logic_vector(to_unsigned(6,8) ,
27123	 => std_logic_vector(to_unsigned(7,8) ,
27124	 => std_logic_vector(to_unsigned(7,8) ,
27125	 => std_logic_vector(to_unsigned(5,8) ,
27126	 => std_logic_vector(to_unsigned(3,8) ,
27127	 => std_logic_vector(to_unsigned(4,8) ,
27128	 => std_logic_vector(to_unsigned(3,8) ,
27129	 => std_logic_vector(to_unsigned(1,8) ,
27130	 => std_logic_vector(to_unsigned(1,8) ,
27131	 => std_logic_vector(to_unsigned(1,8) ,
27132	 => std_logic_vector(to_unsigned(4,8) ,
27133	 => std_logic_vector(to_unsigned(6,8) ,
27134	 => std_logic_vector(to_unsigned(14,8) ,
27135	 => std_logic_vector(to_unsigned(20,8) ,
27136	 => std_logic_vector(to_unsigned(12,8) ,
27137	 => std_logic_vector(to_unsigned(6,8) ,
27138	 => std_logic_vector(to_unsigned(9,8) ,
27139	 => std_logic_vector(to_unsigned(18,8) ,
27140	 => std_logic_vector(to_unsigned(44,8) ,
27141	 => std_logic_vector(to_unsigned(11,8) ,
27142	 => std_logic_vector(to_unsigned(16,8) ,
27143	 => std_logic_vector(to_unsigned(54,8) ,
27144	 => std_logic_vector(to_unsigned(52,8) ,
27145	 => std_logic_vector(to_unsigned(58,8) ,
27146	 => std_logic_vector(to_unsigned(84,8) ,
27147	 => std_logic_vector(to_unsigned(80,8) ,
27148	 => std_logic_vector(to_unsigned(82,8) ,
27149	 => std_logic_vector(to_unsigned(53,8) ,
27150	 => std_logic_vector(to_unsigned(43,8) ,
27151	 => std_logic_vector(to_unsigned(91,8) ,
27152	 => std_logic_vector(to_unsigned(125,8) ,
27153	 => std_logic_vector(to_unsigned(130,8) ,
27154	 => std_logic_vector(to_unsigned(103,8) ,
27155	 => std_logic_vector(to_unsigned(47,8) ,
27156	 => std_logic_vector(to_unsigned(48,8) ,
27157	 => std_logic_vector(to_unsigned(99,8) ,
27158	 => std_logic_vector(to_unsigned(128,8) ,
27159	 => std_logic_vector(to_unsigned(151,8) ,
27160	 => std_logic_vector(to_unsigned(108,8) ,
27161	 => std_logic_vector(to_unsigned(19,8) ,
27162	 => std_logic_vector(to_unsigned(4,8) ,
27163	 => std_logic_vector(to_unsigned(25,8) ,
27164	 => std_logic_vector(to_unsigned(72,8) ,
27165	 => std_logic_vector(to_unsigned(66,8) ,
27166	 => std_logic_vector(to_unsigned(18,8) ,
27167	 => std_logic_vector(to_unsigned(13,8) ,
27168	 => std_logic_vector(to_unsigned(14,8) ,
27169	 => std_logic_vector(to_unsigned(14,8) ,
27170	 => std_logic_vector(to_unsigned(24,8) ,
27171	 => std_logic_vector(to_unsigned(32,8) ,
27172	 => std_logic_vector(to_unsigned(45,8) ,
27173	 => std_logic_vector(to_unsigned(116,8) ,
27174	 => std_logic_vector(to_unsigned(92,8) ,
27175	 => std_logic_vector(to_unsigned(26,8) ,
27176	 => std_logic_vector(to_unsigned(73,8) ,
27177	 => std_logic_vector(to_unsigned(138,8) ,
27178	 => std_logic_vector(to_unsigned(74,8) ,
27179	 => std_logic_vector(to_unsigned(76,8) ,
27180	 => std_logic_vector(to_unsigned(146,8) ,
27181	 => std_logic_vector(to_unsigned(161,8) ,
27182	 => std_logic_vector(to_unsigned(141,8) ,
27183	 => std_logic_vector(to_unsigned(127,8) ,
27184	 => std_logic_vector(to_unsigned(131,8) ,
27185	 => std_logic_vector(to_unsigned(134,8) ,
27186	 => std_logic_vector(to_unsigned(142,8) ,
27187	 => std_logic_vector(to_unsigned(154,8) ,
27188	 => std_logic_vector(to_unsigned(152,8) ,
27189	 => std_logic_vector(to_unsigned(159,8) ,
27190	 => std_logic_vector(to_unsigned(147,8) ,
27191	 => std_logic_vector(to_unsigned(152,8) ,
27192	 => std_logic_vector(to_unsigned(156,8) ,
27193	 => std_logic_vector(to_unsigned(154,8) ,
27194	 => std_logic_vector(to_unsigned(154,8) ,
27195	 => std_logic_vector(to_unsigned(147,8) ,
27196	 => std_logic_vector(to_unsigned(146,8) ,
27197	 => std_logic_vector(to_unsigned(163,8) ,
27198	 => std_logic_vector(to_unsigned(170,8) ,
27199	 => std_logic_vector(to_unsigned(163,8) ,
27200	 => std_logic_vector(to_unsigned(156,8) ,
27201	 => std_logic_vector(to_unsigned(163,8) ,
27202	 => std_logic_vector(to_unsigned(163,8) ,
27203	 => std_logic_vector(to_unsigned(157,8) ,
27204	 => std_logic_vector(to_unsigned(161,8) ,
27205	 => std_logic_vector(to_unsigned(151,8) ,
27206	 => std_logic_vector(to_unsigned(136,8) ,
27207	 => std_logic_vector(to_unsigned(146,8) ,
27208	 => std_logic_vector(to_unsigned(71,8) ,
27209	 => std_logic_vector(to_unsigned(43,8) ,
27210	 => std_logic_vector(to_unsigned(64,8) ,
27211	 => std_logic_vector(to_unsigned(20,8) ,
27212	 => std_logic_vector(to_unsigned(8,8) ,
27213	 => std_logic_vector(to_unsigned(8,8) ,
27214	 => std_logic_vector(to_unsigned(3,8) ,
27215	 => std_logic_vector(to_unsigned(2,8) ,
27216	 => std_logic_vector(to_unsigned(1,8) ,
27217	 => std_logic_vector(to_unsigned(1,8) ,
27218	 => std_logic_vector(to_unsigned(0,8) ,
27219	 => std_logic_vector(to_unsigned(0,8) ,
27220	 => std_logic_vector(to_unsigned(1,8) ,
27221	 => std_logic_vector(to_unsigned(1,8) ,
27222	 => std_logic_vector(to_unsigned(1,8) ,
27223	 => std_logic_vector(to_unsigned(0,8) ,
27224	 => std_logic_vector(to_unsigned(0,8) ,
27225	 => std_logic_vector(to_unsigned(1,8) ,
27226	 => std_logic_vector(to_unsigned(1,8) ,
27227	 => std_logic_vector(to_unsigned(0,8) ,
27228	 => std_logic_vector(to_unsigned(0,8) ,
27229	 => std_logic_vector(to_unsigned(0,8) ,
27230	 => std_logic_vector(to_unsigned(1,8) ,
27231	 => std_logic_vector(to_unsigned(2,8) ,
27232	 => std_logic_vector(to_unsigned(11,8) ,
27233	 => std_logic_vector(to_unsigned(41,8) ,
27234	 => std_logic_vector(to_unsigned(67,8) ,
27235	 => std_logic_vector(to_unsigned(81,8) ,
27236	 => std_logic_vector(to_unsigned(80,8) ,
27237	 => std_logic_vector(to_unsigned(92,8) ,
27238	 => std_logic_vector(to_unsigned(111,8) ,
27239	 => std_logic_vector(to_unsigned(116,8) ,
27240	 => std_logic_vector(to_unsigned(112,8) ,
27241	 => std_logic_vector(to_unsigned(97,8) ,
27242	 => std_logic_vector(to_unsigned(76,8) ,
27243	 => std_logic_vector(to_unsigned(29,8) ,
27244	 => std_logic_vector(to_unsigned(3,8) ,
27245	 => std_logic_vector(to_unsigned(0,8) ,
27246	 => std_logic_vector(to_unsigned(0,8) ,
27247	 => std_logic_vector(to_unsigned(1,8) ,
27248	 => std_logic_vector(to_unsigned(1,8) ,
27249	 => std_logic_vector(to_unsigned(1,8) ,
27250	 => std_logic_vector(to_unsigned(1,8) ,
27251	 => std_logic_vector(to_unsigned(3,8) ,
27252	 => std_logic_vector(to_unsigned(53,8) ,
27253	 => std_logic_vector(to_unsigned(118,8) ,
27254	 => std_logic_vector(to_unsigned(111,8) ,
27255	 => std_logic_vector(to_unsigned(105,8) ,
27256	 => std_logic_vector(to_unsigned(86,8) ,
27257	 => std_logic_vector(to_unsigned(23,8) ,
27258	 => std_logic_vector(to_unsigned(8,8) ,
27259	 => std_logic_vector(to_unsigned(9,8) ,
27260	 => std_logic_vector(to_unsigned(18,8) ,
27261	 => std_logic_vector(to_unsigned(19,8) ,
27262	 => std_logic_vector(to_unsigned(18,8) ,
27263	 => std_logic_vector(to_unsigned(14,8) ,
27264	 => std_logic_vector(to_unsigned(9,8) ,
27265	 => std_logic_vector(to_unsigned(10,8) ,
27266	 => std_logic_vector(to_unsigned(11,8) ,
27267	 => std_logic_vector(to_unsigned(9,8) ,
27268	 => std_logic_vector(to_unsigned(10,8) ,
27269	 => std_logic_vector(to_unsigned(11,8) ,
27270	 => std_logic_vector(to_unsigned(10,8) ,
27271	 => std_logic_vector(to_unsigned(7,8) ,
27272	 => std_logic_vector(to_unsigned(3,8) ,
27273	 => std_logic_vector(to_unsigned(4,8) ,
27274	 => std_logic_vector(to_unsigned(3,8) ,
27275	 => std_logic_vector(to_unsigned(4,8) ,
27276	 => std_logic_vector(to_unsigned(5,8) ,
27277	 => std_logic_vector(to_unsigned(3,8) ,
27278	 => std_logic_vector(to_unsigned(2,8) ,
27279	 => std_logic_vector(to_unsigned(19,8) ,
27280	 => std_logic_vector(to_unsigned(124,8) ,
27281	 => std_logic_vector(to_unsigned(108,8) ,
27282	 => std_logic_vector(to_unsigned(66,8) ,
27283	 => std_logic_vector(to_unsigned(57,8) ,
27284	 => std_logic_vector(to_unsigned(49,8) ,
27285	 => std_logic_vector(to_unsigned(33,8) ,
27286	 => std_logic_vector(to_unsigned(22,8) ,
27287	 => std_logic_vector(to_unsigned(5,8) ,
27288	 => std_logic_vector(to_unsigned(32,8) ,
27289	 => std_logic_vector(to_unsigned(86,8) ,
27290	 => std_logic_vector(to_unsigned(35,8) ,
27291	 => std_logic_vector(to_unsigned(56,8) ,
27292	 => std_logic_vector(to_unsigned(78,8) ,
27293	 => std_logic_vector(to_unsigned(122,8) ,
27294	 => std_logic_vector(to_unsigned(170,8) ,
27295	 => std_logic_vector(to_unsigned(152,8) ,
27296	 => std_logic_vector(to_unsigned(118,8) ,
27297	 => std_logic_vector(to_unsigned(144,8) ,
27298	 => std_logic_vector(to_unsigned(147,8) ,
27299	 => std_logic_vector(to_unsigned(149,8) ,
27300	 => std_logic_vector(to_unsigned(149,8) ,
27301	 => std_logic_vector(to_unsigned(33,8) ,
27302	 => std_logic_vector(to_unsigned(26,8) ,
27303	 => std_logic_vector(to_unsigned(124,8) ,
27304	 => std_logic_vector(to_unsigned(78,8) ,
27305	 => std_logic_vector(to_unsigned(90,8) ,
27306	 => std_logic_vector(to_unsigned(58,8) ,
27307	 => std_logic_vector(to_unsigned(48,8) ,
27308	 => std_logic_vector(to_unsigned(86,8) ,
27309	 => std_logic_vector(to_unsigned(118,8) ,
27310	 => std_logic_vector(to_unsigned(116,8) ,
27311	 => std_logic_vector(to_unsigned(32,8) ,
27312	 => std_logic_vector(to_unsigned(7,8) ,
27313	 => std_logic_vector(to_unsigned(3,8) ,
27314	 => std_logic_vector(to_unsigned(2,8) ,
27315	 => std_logic_vector(to_unsigned(0,8) ,
27316	 => std_logic_vector(to_unsigned(0,8) ,
27317	 => std_logic_vector(to_unsigned(1,8) ,
27318	 => std_logic_vector(to_unsigned(1,8) ,
27319	 => std_logic_vector(to_unsigned(1,8) ,
27320	 => std_logic_vector(to_unsigned(1,8) ,
27321	 => std_logic_vector(to_unsigned(1,8) ,
27322	 => std_logic_vector(to_unsigned(1,8) ,
27323	 => std_logic_vector(to_unsigned(1,8) ,
27324	 => std_logic_vector(to_unsigned(2,8) ,
27325	 => std_logic_vector(to_unsigned(2,8) ,
27326	 => std_logic_vector(to_unsigned(1,8) ,
27327	 => std_logic_vector(to_unsigned(2,8) ,
27328	 => std_logic_vector(to_unsigned(9,8) ,
27329	 => std_logic_vector(to_unsigned(36,8) ,
27330	 => std_logic_vector(to_unsigned(54,8) ,
27331	 => std_logic_vector(to_unsigned(87,8) ,
27332	 => std_logic_vector(to_unsigned(103,8) ,
27333	 => std_logic_vector(to_unsigned(124,8) ,
27334	 => std_logic_vector(to_unsigned(99,8) ,
27335	 => std_logic_vector(to_unsigned(63,8) ,
27336	 => std_logic_vector(to_unsigned(87,8) ,
27337	 => std_logic_vector(to_unsigned(104,8) ,
27338	 => std_logic_vector(to_unsigned(52,8) ,
27339	 => std_logic_vector(to_unsigned(15,8) ,
27340	 => std_logic_vector(to_unsigned(11,8) ,
27341	 => std_logic_vector(to_unsigned(4,8) ,
27342	 => std_logic_vector(to_unsigned(4,8) ,
27343	 => std_logic_vector(to_unsigned(8,8) ,
27344	 => std_logic_vector(to_unsigned(14,8) ,
27345	 => std_logic_vector(to_unsigned(21,8) ,
27346	 => std_logic_vector(to_unsigned(35,8) ,
27347	 => std_logic_vector(to_unsigned(20,8) ,
27348	 => std_logic_vector(to_unsigned(15,8) ,
27349	 => std_logic_vector(to_unsigned(21,8) ,
27350	 => std_logic_vector(to_unsigned(20,8) ,
27351	 => std_logic_vector(to_unsigned(12,8) ,
27352	 => std_logic_vector(to_unsigned(9,8) ,
27353	 => std_logic_vector(to_unsigned(9,8) ,
27354	 => std_logic_vector(to_unsigned(12,8) ,
27355	 => std_logic_vector(to_unsigned(7,8) ,
27356	 => std_logic_vector(to_unsigned(3,8) ,
27357	 => std_logic_vector(to_unsigned(14,8) ,
27358	 => std_logic_vector(to_unsigned(28,8) ,
27359	 => std_logic_vector(to_unsigned(34,8) ,
27360	 => std_logic_vector(to_unsigned(47,8) ,
27361	 => std_logic_vector(to_unsigned(45,8) ,
27362	 => std_logic_vector(to_unsigned(23,8) ,
27363	 => std_logic_vector(to_unsigned(23,8) ,
27364	 => std_logic_vector(to_unsigned(15,8) ,
27365	 => std_logic_vector(to_unsigned(51,8) ,
27366	 => std_logic_vector(to_unsigned(82,8) ,
27367	 => std_logic_vector(to_unsigned(62,8) ,
27368	 => std_logic_vector(to_unsigned(9,8) ,
27369	 => std_logic_vector(to_unsigned(7,8) ,
27370	 => std_logic_vector(to_unsigned(20,8) ,
27371	 => std_logic_vector(to_unsigned(26,8) ,
27372	 => std_logic_vector(to_unsigned(27,8) ,
27373	 => std_logic_vector(to_unsigned(24,8) ,
27374	 => std_logic_vector(to_unsigned(18,8) ,
27375	 => std_logic_vector(to_unsigned(10,8) ,
27376	 => std_logic_vector(to_unsigned(12,8) ,
27377	 => std_logic_vector(to_unsigned(20,8) ,
27378	 => std_logic_vector(to_unsigned(23,8) ,
27379	 => std_logic_vector(to_unsigned(27,8) ,
27380	 => std_logic_vector(to_unsigned(17,8) ,
27381	 => std_logic_vector(to_unsigned(7,8) ,
27382	 => std_logic_vector(to_unsigned(4,8) ,
27383	 => std_logic_vector(to_unsigned(1,8) ,
27384	 => std_logic_vector(to_unsigned(4,8) ,
27385	 => std_logic_vector(to_unsigned(13,8) ,
27386	 => std_logic_vector(to_unsigned(11,8) ,
27387	 => std_logic_vector(to_unsigned(85,8) ,
27388	 => std_logic_vector(to_unsigned(142,8) ,
27389	 => std_logic_vector(to_unsigned(119,8) ,
27390	 => std_logic_vector(to_unsigned(119,8) ,
27391	 => std_logic_vector(to_unsigned(109,8) ,
27392	 => std_logic_vector(to_unsigned(142,8) ,
27393	 => std_logic_vector(to_unsigned(138,8) ,
27394	 => std_logic_vector(to_unsigned(119,8) ,
27395	 => std_logic_vector(to_unsigned(119,8) ,
27396	 => std_logic_vector(to_unsigned(122,8) ,
27397	 => std_logic_vector(to_unsigned(163,8) ,
27398	 => std_logic_vector(to_unsigned(47,8) ,
27399	 => std_logic_vector(to_unsigned(4,8) ,
27400	 => std_logic_vector(to_unsigned(6,8) ,
27401	 => std_logic_vector(to_unsigned(27,8) ,
27402	 => std_logic_vector(to_unsigned(109,8) ,
27403	 => std_logic_vector(to_unsigned(134,8) ,
27404	 => std_logic_vector(to_unsigned(146,8) ,
27405	 => std_logic_vector(to_unsigned(156,8) ,
27406	 => std_logic_vector(to_unsigned(131,8) ,
27407	 => std_logic_vector(to_unsigned(16,8) ,
27408	 => std_logic_vector(to_unsigned(19,8) ,
27409	 => std_logic_vector(to_unsigned(114,8) ,
27410	 => std_logic_vector(to_unsigned(111,8) ,
27411	 => std_logic_vector(to_unsigned(149,8) ,
27412	 => std_logic_vector(to_unsigned(156,8) ,
27413	 => std_logic_vector(to_unsigned(146,8) ,
27414	 => std_logic_vector(to_unsigned(133,8) ,
27415	 => std_logic_vector(to_unsigned(128,8) ,
27416	 => std_logic_vector(to_unsigned(133,8) ,
27417	 => std_logic_vector(to_unsigned(131,8) ,
27418	 => std_logic_vector(to_unsigned(142,8) ,
27419	 => std_logic_vector(to_unsigned(35,8) ,
27420	 => std_logic_vector(to_unsigned(5,8) ,
27421	 => std_logic_vector(to_unsigned(6,8) ,
27422	 => std_logic_vector(to_unsigned(4,8) ,
27423	 => std_logic_vector(to_unsigned(32,8) ,
27424	 => std_logic_vector(to_unsigned(144,8) ,
27425	 => std_logic_vector(to_unsigned(147,8) ,
27426	 => std_logic_vector(to_unsigned(35,8) ,
27427	 => std_logic_vector(to_unsigned(22,8) ,
27428	 => std_logic_vector(to_unsigned(27,8) ,
27429	 => std_logic_vector(to_unsigned(22,8) ,
27430	 => std_logic_vector(to_unsigned(18,8) ,
27431	 => std_logic_vector(to_unsigned(18,8) ,
27432	 => std_logic_vector(to_unsigned(20,8) ,
27433	 => std_logic_vector(to_unsigned(93,8) ,
27434	 => std_logic_vector(to_unsigned(188,8) ,
27435	 => std_logic_vector(to_unsigned(103,8) ,
27436	 => std_logic_vector(to_unsigned(27,8) ,
27437	 => std_logic_vector(to_unsigned(38,8) ,
27438	 => std_logic_vector(to_unsigned(51,8) ,
27439	 => std_logic_vector(to_unsigned(36,8) ,
27440	 => std_logic_vector(to_unsigned(12,8) ,
27441	 => std_logic_vector(to_unsigned(9,8) ,
27442	 => std_logic_vector(to_unsigned(12,8) ,
27443	 => std_logic_vector(to_unsigned(8,8) ,
27444	 => std_logic_vector(to_unsigned(7,8) ,
27445	 => std_logic_vector(to_unsigned(5,8) ,
27446	 => std_logic_vector(to_unsigned(5,8) ,
27447	 => std_logic_vector(to_unsigned(2,8) ,
27448	 => std_logic_vector(to_unsigned(8,8) ,
27449	 => std_logic_vector(to_unsigned(13,8) ,
27450	 => std_logic_vector(to_unsigned(1,8) ,
27451	 => std_logic_vector(to_unsigned(2,8) ,
27452	 => std_logic_vector(to_unsigned(6,8) ,
27453	 => std_logic_vector(to_unsigned(8,8) ,
27454	 => std_logic_vector(to_unsigned(4,8) ,
27455	 => std_logic_vector(to_unsigned(11,8) ,
27456	 => std_logic_vector(to_unsigned(14,8) ,
27457	 => std_logic_vector(to_unsigned(4,8) ,
27458	 => std_logic_vector(to_unsigned(8,8) ,
27459	 => std_logic_vector(to_unsigned(13,8) ,
27460	 => std_logic_vector(to_unsigned(22,8) ,
27461	 => std_logic_vector(to_unsigned(6,8) ,
27462	 => std_logic_vector(to_unsigned(23,8) ,
27463	 => std_logic_vector(to_unsigned(68,8) ,
27464	 => std_logic_vector(to_unsigned(53,8) ,
27465	 => std_logic_vector(to_unsigned(65,8) ,
27466	 => std_logic_vector(to_unsigned(65,8) ,
27467	 => std_logic_vector(to_unsigned(60,8) ,
27468	 => std_logic_vector(to_unsigned(64,8) ,
27469	 => std_logic_vector(to_unsigned(37,8) ,
27470	 => std_logic_vector(to_unsigned(20,8) ,
27471	 => std_logic_vector(to_unsigned(41,8) ,
27472	 => std_logic_vector(to_unsigned(111,8) ,
27473	 => std_logic_vector(to_unsigned(127,8) ,
27474	 => std_logic_vector(to_unsigned(68,8) ,
27475	 => std_logic_vector(to_unsigned(17,8) ,
27476	 => std_logic_vector(to_unsigned(3,8) ,
27477	 => std_logic_vector(to_unsigned(61,8) ,
27478	 => std_logic_vector(to_unsigned(121,8) ,
27479	 => std_logic_vector(to_unsigned(121,8) ,
27480	 => std_logic_vector(to_unsigned(80,8) ,
27481	 => std_logic_vector(to_unsigned(25,8) ,
27482	 => std_logic_vector(to_unsigned(30,8) ,
27483	 => std_logic_vector(to_unsigned(46,8) ,
27484	 => std_logic_vector(to_unsigned(27,8) ,
27485	 => std_logic_vector(to_unsigned(7,8) ,
27486	 => std_logic_vector(to_unsigned(1,8) ,
27487	 => std_logic_vector(to_unsigned(1,8) ,
27488	 => std_logic_vector(to_unsigned(26,8) ,
27489	 => std_logic_vector(to_unsigned(30,8) ,
27490	 => std_logic_vector(to_unsigned(18,8) ,
27491	 => std_logic_vector(to_unsigned(25,8) ,
27492	 => std_logic_vector(to_unsigned(62,8) ,
27493	 => std_logic_vector(to_unsigned(122,8) ,
27494	 => std_logic_vector(to_unsigned(61,8) ,
27495	 => std_logic_vector(to_unsigned(19,8) ,
27496	 => std_logic_vector(to_unsigned(82,8) ,
27497	 => std_logic_vector(to_unsigned(138,8) ,
27498	 => std_logic_vector(to_unsigned(59,8) ,
27499	 => std_logic_vector(to_unsigned(64,8) ,
27500	 => std_logic_vector(to_unsigned(164,8) ,
27501	 => std_logic_vector(to_unsigned(163,8) ,
27502	 => std_logic_vector(to_unsigned(156,8) ,
27503	 => std_logic_vector(to_unsigned(154,8) ,
27504	 => std_logic_vector(to_unsigned(144,8) ,
27505	 => std_logic_vector(to_unsigned(149,8) ,
27506	 => std_logic_vector(to_unsigned(151,8) ,
27507	 => std_logic_vector(to_unsigned(154,8) ,
27508	 => std_logic_vector(to_unsigned(151,8) ,
27509	 => std_logic_vector(to_unsigned(154,8) ,
27510	 => std_logic_vector(to_unsigned(156,8) ,
27511	 => std_logic_vector(to_unsigned(159,8) ,
27512	 => std_logic_vector(to_unsigned(159,8) ,
27513	 => std_logic_vector(to_unsigned(157,8) ,
27514	 => std_logic_vector(to_unsigned(156,8) ,
27515	 => std_logic_vector(to_unsigned(152,8) ,
27516	 => std_logic_vector(to_unsigned(152,8) ,
27517	 => std_logic_vector(to_unsigned(164,8) ,
27518	 => std_logic_vector(to_unsigned(168,8) ,
27519	 => std_logic_vector(to_unsigned(161,8) ,
27520	 => std_logic_vector(to_unsigned(163,8) ,
27521	 => std_logic_vector(to_unsigned(166,8) ,
27522	 => std_logic_vector(to_unsigned(164,8) ,
27523	 => std_logic_vector(to_unsigned(157,8) ,
27524	 => std_logic_vector(to_unsigned(141,8) ,
27525	 => std_logic_vector(to_unsigned(139,8) ,
27526	 => std_logic_vector(to_unsigned(136,8) ,
27527	 => std_logic_vector(to_unsigned(173,8) ,
27528	 => std_logic_vector(to_unsigned(198,8) ,
27529	 => std_logic_vector(to_unsigned(196,8) ,
27530	 => std_logic_vector(to_unsigned(179,8) ,
27531	 => std_logic_vector(to_unsigned(166,8) ,
27532	 => std_logic_vector(to_unsigned(152,8) ,
27533	 => std_logic_vector(to_unsigned(134,8) ,
27534	 => std_logic_vector(to_unsigned(111,8) ,
27535	 => std_logic_vector(to_unsigned(93,8) ,
27536	 => std_logic_vector(to_unsigned(79,8) ,
27537	 => std_logic_vector(to_unsigned(67,8) ,
27538	 => std_logic_vector(to_unsigned(56,8) ,
27539	 => std_logic_vector(to_unsigned(46,8) ,
27540	 => std_logic_vector(to_unsigned(36,8) ,
27541	 => std_logic_vector(to_unsigned(31,8) ,
27542	 => std_logic_vector(to_unsigned(32,8) ,
27543	 => std_logic_vector(to_unsigned(28,8) ,
27544	 => std_logic_vector(to_unsigned(15,8) ,
27545	 => std_logic_vector(to_unsigned(2,8) ,
27546	 => std_logic_vector(to_unsigned(1,8) ,
27547	 => std_logic_vector(to_unsigned(1,8) ,
27548	 => std_logic_vector(to_unsigned(0,8) ,
27549	 => std_logic_vector(to_unsigned(2,8) ,
27550	 => std_logic_vector(to_unsigned(4,8) ,
27551	 => std_logic_vector(to_unsigned(3,8) ,
27552	 => std_logic_vector(to_unsigned(8,8) ,
27553	 => std_logic_vector(to_unsigned(25,8) ,
27554	 => std_logic_vector(to_unsigned(15,8) ,
27555	 => std_logic_vector(to_unsigned(18,8) ,
27556	 => std_logic_vector(to_unsigned(26,8) ,
27557	 => std_logic_vector(to_unsigned(25,8) ,
27558	 => std_logic_vector(to_unsigned(20,8) ,
27559	 => std_logic_vector(to_unsigned(29,8) ,
27560	 => std_logic_vector(to_unsigned(42,8) ,
27561	 => std_logic_vector(to_unsigned(59,8) ,
27562	 => std_logic_vector(to_unsigned(60,8) ,
27563	 => std_logic_vector(to_unsigned(13,8) ,
27564	 => std_logic_vector(to_unsigned(1,8) ,
27565	 => std_logic_vector(to_unsigned(1,8) ,
27566	 => std_logic_vector(to_unsigned(1,8) ,
27567	 => std_logic_vector(to_unsigned(1,8) ,
27568	 => std_logic_vector(to_unsigned(2,8) ,
27569	 => std_logic_vector(to_unsigned(2,8) ,
27570	 => std_logic_vector(to_unsigned(1,8) ,
27571	 => std_logic_vector(to_unsigned(1,8) ,
27572	 => std_logic_vector(to_unsigned(37,8) ,
27573	 => std_logic_vector(to_unsigned(100,8) ,
27574	 => std_logic_vector(to_unsigned(103,8) ,
27575	 => std_logic_vector(to_unsigned(108,8) ,
27576	 => std_logic_vector(to_unsigned(80,8) ,
27577	 => std_logic_vector(to_unsigned(18,8) ,
27578	 => std_logic_vector(to_unsigned(12,8) ,
27579	 => std_logic_vector(to_unsigned(6,8) ,
27580	 => std_logic_vector(to_unsigned(18,8) ,
27581	 => std_logic_vector(to_unsigned(35,8) ,
27582	 => std_logic_vector(to_unsigned(30,8) ,
27583	 => std_logic_vector(to_unsigned(25,8) ,
27584	 => std_logic_vector(to_unsigned(19,8) ,
27585	 => std_logic_vector(to_unsigned(14,8) ,
27586	 => std_logic_vector(to_unsigned(14,8) ,
27587	 => std_logic_vector(to_unsigned(11,8) ,
27588	 => std_logic_vector(to_unsigned(10,8) ,
27589	 => std_logic_vector(to_unsigned(12,8) ,
27590	 => std_logic_vector(to_unsigned(10,8) ,
27591	 => std_logic_vector(to_unsigned(5,8) ,
27592	 => std_logic_vector(to_unsigned(5,8) ,
27593	 => std_logic_vector(to_unsigned(4,8) ,
27594	 => std_logic_vector(to_unsigned(2,8) ,
27595	 => std_logic_vector(to_unsigned(6,8) ,
27596	 => std_logic_vector(to_unsigned(9,8) ,
27597	 => std_logic_vector(to_unsigned(5,8) ,
27598	 => std_logic_vector(to_unsigned(2,8) ,
27599	 => std_logic_vector(to_unsigned(65,8) ,
27600	 => std_logic_vector(to_unsigned(164,8) ,
27601	 => std_logic_vector(to_unsigned(127,8) ,
27602	 => std_logic_vector(to_unsigned(69,8) ,
27603	 => std_logic_vector(to_unsigned(62,8) ,
27604	 => std_logic_vector(to_unsigned(49,8) ,
27605	 => std_logic_vector(to_unsigned(28,8) ,
27606	 => std_logic_vector(to_unsigned(8,8) ,
27607	 => std_logic_vector(to_unsigned(21,8) ,
27608	 => std_logic_vector(to_unsigned(93,8) ,
27609	 => std_logic_vector(to_unsigned(107,8) ,
27610	 => std_logic_vector(to_unsigned(45,8) ,
27611	 => std_logic_vector(to_unsigned(64,8) ,
27612	 => std_logic_vector(to_unsigned(125,8) ,
27613	 => std_logic_vector(to_unsigned(136,8) ,
27614	 => std_logic_vector(to_unsigned(163,8) ,
27615	 => std_logic_vector(to_unsigned(134,8) ,
27616	 => std_logic_vector(to_unsigned(71,8) ,
27617	 => std_logic_vector(to_unsigned(99,8) ,
27618	 => std_logic_vector(to_unsigned(127,8) ,
27619	 => std_logic_vector(to_unsigned(149,8) ,
27620	 => std_logic_vector(to_unsigned(144,8) ,
27621	 => std_logic_vector(to_unsigned(55,8) ,
27622	 => std_logic_vector(to_unsigned(32,8) ,
27623	 => std_logic_vector(to_unsigned(96,8) ,
27624	 => std_logic_vector(to_unsigned(91,8) ,
27625	 => std_logic_vector(to_unsigned(91,8) ,
27626	 => std_logic_vector(to_unsigned(66,8) ,
27627	 => std_logic_vector(to_unsigned(124,8) ,
27628	 => std_logic_vector(to_unsigned(82,8) ,
27629	 => std_logic_vector(to_unsigned(44,8) ,
27630	 => std_logic_vector(to_unsigned(131,8) ,
27631	 => std_logic_vector(to_unsigned(95,8) ,
27632	 => std_logic_vector(to_unsigned(32,8) ,
27633	 => std_logic_vector(to_unsigned(3,8) ,
27634	 => std_logic_vector(to_unsigned(1,8) ,
27635	 => std_logic_vector(to_unsigned(0,8) ,
27636	 => std_logic_vector(to_unsigned(0,8) ,
27637	 => std_logic_vector(to_unsigned(1,8) ,
27638	 => std_logic_vector(to_unsigned(1,8) ,
27639	 => std_logic_vector(to_unsigned(1,8) ,
27640	 => std_logic_vector(to_unsigned(1,8) ,
27641	 => std_logic_vector(to_unsigned(2,8) ,
27642	 => std_logic_vector(to_unsigned(2,8) ,
27643	 => std_logic_vector(to_unsigned(2,8) ,
27644	 => std_logic_vector(to_unsigned(2,8) ,
27645	 => std_logic_vector(to_unsigned(2,8) ,
27646	 => std_logic_vector(to_unsigned(2,8) ,
27647	 => std_logic_vector(to_unsigned(3,8) ,
27648	 => std_logic_vector(to_unsigned(9,8) ,
27649	 => std_logic_vector(to_unsigned(46,8) ,
27650	 => std_logic_vector(to_unsigned(124,8) ,
27651	 => std_logic_vector(to_unsigned(138,8) ,
27652	 => std_logic_vector(to_unsigned(107,8) ,
27653	 => std_logic_vector(to_unsigned(92,8) ,
27654	 => std_logic_vector(to_unsigned(33,8) ,
27655	 => std_logic_vector(to_unsigned(4,8) ,
27656	 => std_logic_vector(to_unsigned(38,8) ,
27657	 => std_logic_vector(to_unsigned(125,8) ,
27658	 => std_logic_vector(to_unsigned(67,8) ,
27659	 => std_logic_vector(to_unsigned(14,8) ,
27660	 => std_logic_vector(to_unsigned(15,8) ,
27661	 => std_logic_vector(to_unsigned(6,8) ,
27662	 => std_logic_vector(to_unsigned(2,8) ,
27663	 => std_logic_vector(to_unsigned(4,8) ,
27664	 => std_logic_vector(to_unsigned(9,8) ,
27665	 => std_logic_vector(to_unsigned(25,8) ,
27666	 => std_logic_vector(to_unsigned(38,8) ,
27667	 => std_logic_vector(to_unsigned(23,8) ,
27668	 => std_logic_vector(to_unsigned(20,8) ,
27669	 => std_logic_vector(to_unsigned(27,8) ,
27670	 => std_logic_vector(to_unsigned(17,8) ,
27671	 => std_logic_vector(to_unsigned(10,8) ,
27672	 => std_logic_vector(to_unsigned(11,8) ,
27673	 => std_logic_vector(to_unsigned(10,8) ,
27674	 => std_logic_vector(to_unsigned(8,8) ,
27675	 => std_logic_vector(to_unsigned(6,8) ,
27676	 => std_logic_vector(to_unsigned(5,8) ,
27677	 => std_logic_vector(to_unsigned(27,8) ,
27678	 => std_logic_vector(to_unsigned(32,8) ,
27679	 => std_logic_vector(to_unsigned(39,8) ,
27680	 => std_logic_vector(to_unsigned(47,8) ,
27681	 => std_logic_vector(to_unsigned(60,8) ,
27682	 => std_logic_vector(to_unsigned(26,8) ,
27683	 => std_logic_vector(to_unsigned(13,8) ,
27684	 => std_logic_vector(to_unsigned(17,8) ,
27685	 => std_logic_vector(to_unsigned(58,8) ,
27686	 => std_logic_vector(to_unsigned(95,8) ,
27687	 => std_logic_vector(to_unsigned(71,8) ,
27688	 => std_logic_vector(to_unsigned(33,8) ,
27689	 => std_logic_vector(to_unsigned(24,8) ,
27690	 => std_logic_vector(to_unsigned(8,8) ,
27691	 => std_logic_vector(to_unsigned(12,8) ,
27692	 => std_logic_vector(to_unsigned(20,8) ,
27693	 => std_logic_vector(to_unsigned(24,8) ,
27694	 => std_logic_vector(to_unsigned(22,8) ,
27695	 => std_logic_vector(to_unsigned(10,8) ,
27696	 => std_logic_vector(to_unsigned(6,8) ,
27697	 => std_logic_vector(to_unsigned(12,8) ,
27698	 => std_logic_vector(to_unsigned(17,8) ,
27699	 => std_logic_vector(to_unsigned(17,8) ,
27700	 => std_logic_vector(to_unsigned(8,8) ,
27701	 => std_logic_vector(to_unsigned(4,8) ,
27702	 => std_logic_vector(to_unsigned(3,8) ,
27703	 => std_logic_vector(to_unsigned(3,8) ,
27704	 => std_logic_vector(to_unsigned(3,8) ,
27705	 => std_logic_vector(to_unsigned(8,8) ,
27706	 => std_logic_vector(to_unsigned(19,8) ,
27707	 => std_logic_vector(to_unsigned(107,8) ,
27708	 => std_logic_vector(to_unsigned(142,8) ,
27709	 => std_logic_vector(to_unsigned(119,8) ,
27710	 => std_logic_vector(to_unsigned(139,8) ,
27711	 => std_logic_vector(to_unsigned(124,8) ,
27712	 => std_logic_vector(to_unsigned(141,8) ,
27713	 => std_logic_vector(to_unsigned(146,8) ,
27714	 => std_logic_vector(to_unsigned(151,8) ,
27715	 => std_logic_vector(to_unsigned(147,8) ,
27716	 => std_logic_vector(to_unsigned(115,8) ,
27717	 => std_logic_vector(to_unsigned(156,8) ,
27718	 => std_logic_vector(to_unsigned(116,8) ,
27719	 => std_logic_vector(to_unsigned(9,8) ,
27720	 => std_logic_vector(to_unsigned(9,8) ,
27721	 => std_logic_vector(to_unsigned(87,8) ,
27722	 => std_logic_vector(to_unsigned(151,8) ,
27723	 => std_logic_vector(to_unsigned(146,8) ,
27724	 => std_logic_vector(to_unsigned(152,8) ,
27725	 => std_logic_vector(to_unsigned(147,8) ,
27726	 => std_logic_vector(to_unsigned(144,8) ,
27727	 => std_logic_vector(to_unsigned(76,8) ,
27728	 => std_logic_vector(to_unsigned(55,8) ,
27729	 => std_logic_vector(to_unsigned(87,8) ,
27730	 => std_logic_vector(to_unsigned(116,8) ,
27731	 => std_logic_vector(to_unsigned(152,8) ,
27732	 => std_logic_vector(to_unsigned(151,8) ,
27733	 => std_logic_vector(to_unsigned(151,8) ,
27734	 => std_logic_vector(to_unsigned(138,8) ,
27735	 => std_logic_vector(to_unsigned(125,8) ,
27736	 => std_logic_vector(to_unsigned(128,8) ,
27737	 => std_logic_vector(to_unsigned(131,8) ,
27738	 => std_logic_vector(to_unsigned(124,8) ,
27739	 => std_logic_vector(to_unsigned(18,8) ,
27740	 => std_logic_vector(to_unsigned(7,8) ,
27741	 => std_logic_vector(to_unsigned(8,8) ,
27742	 => std_logic_vector(to_unsigned(2,8) ,
27743	 => std_logic_vector(to_unsigned(38,8) ,
27744	 => std_logic_vector(to_unsigned(163,8) ,
27745	 => std_logic_vector(to_unsigned(159,8) ,
27746	 => std_logic_vector(to_unsigned(38,8) ,
27747	 => std_logic_vector(to_unsigned(12,8) ,
27748	 => std_logic_vector(to_unsigned(29,8) ,
27749	 => std_logic_vector(to_unsigned(33,8) ,
27750	 => std_logic_vector(to_unsigned(30,8) ,
27751	 => std_logic_vector(to_unsigned(20,8) ,
27752	 => std_logic_vector(to_unsigned(66,8) ,
27753	 => std_logic_vector(to_unsigned(164,8) ,
27754	 => std_logic_vector(to_unsigned(171,8) ,
27755	 => std_logic_vector(to_unsigned(59,8) ,
27756	 => std_logic_vector(to_unsigned(14,8) ,
27757	 => std_logic_vector(to_unsigned(27,8) ,
27758	 => std_logic_vector(to_unsigned(39,8) ,
27759	 => std_logic_vector(to_unsigned(24,8) ,
27760	 => std_logic_vector(to_unsigned(13,8) ,
27761	 => std_logic_vector(to_unsigned(8,8) ,
27762	 => std_logic_vector(to_unsigned(8,8) ,
27763	 => std_logic_vector(to_unsigned(9,8) ,
27764	 => std_logic_vector(to_unsigned(5,8) ,
27765	 => std_logic_vector(to_unsigned(5,8) ,
27766	 => std_logic_vector(to_unsigned(4,8) ,
27767	 => std_logic_vector(to_unsigned(1,8) ,
27768	 => std_logic_vector(to_unsigned(3,8) ,
27769	 => std_logic_vector(to_unsigned(64,8) ,
27770	 => std_logic_vector(to_unsigned(25,8) ,
27771	 => std_logic_vector(to_unsigned(4,8) ,
27772	 => std_logic_vector(to_unsigned(9,8) ,
27773	 => std_logic_vector(to_unsigned(19,8) ,
27774	 => std_logic_vector(to_unsigned(10,8) ,
27775	 => std_logic_vector(to_unsigned(10,8) ,
27776	 => std_logic_vector(to_unsigned(12,8) ,
27777	 => std_logic_vector(to_unsigned(6,8) ,
27778	 => std_logic_vector(to_unsigned(7,8) ,
27779	 => std_logic_vector(to_unsigned(10,8) ,
27780	 => std_logic_vector(to_unsigned(17,8) ,
27781	 => std_logic_vector(to_unsigned(5,8) ,
27782	 => std_logic_vector(to_unsigned(21,8) ,
27783	 => std_logic_vector(to_unsigned(65,8) ,
27784	 => std_logic_vector(to_unsigned(51,8) ,
27785	 => std_logic_vector(to_unsigned(56,8) ,
27786	 => std_logic_vector(to_unsigned(56,8) ,
27787	 => std_logic_vector(to_unsigned(52,8) ,
27788	 => std_logic_vector(to_unsigned(58,8) ,
27789	 => std_logic_vector(to_unsigned(35,8) ,
27790	 => std_logic_vector(to_unsigned(15,8) ,
27791	 => std_logic_vector(to_unsigned(28,8) ,
27792	 => std_logic_vector(to_unsigned(25,8) ,
27793	 => std_logic_vector(to_unsigned(52,8) ,
27794	 => std_logic_vector(to_unsigned(22,8) ,
27795	 => std_logic_vector(to_unsigned(2,8) ,
27796	 => std_logic_vector(to_unsigned(2,8) ,
27797	 => std_logic_vector(to_unsigned(5,8) ,
27798	 => std_logic_vector(to_unsigned(10,8) ,
27799	 => std_logic_vector(to_unsigned(12,8) ,
27800	 => std_logic_vector(to_unsigned(6,8) ,
27801	 => std_logic_vector(to_unsigned(7,8) ,
27802	 => std_logic_vector(to_unsigned(7,8) ,
27803	 => std_logic_vector(to_unsigned(2,8) ,
27804	 => std_logic_vector(to_unsigned(1,8) ,
27805	 => std_logic_vector(to_unsigned(1,8) ,
27806	 => std_logic_vector(to_unsigned(2,8) ,
27807	 => std_logic_vector(to_unsigned(1,8) ,
27808	 => std_logic_vector(to_unsigned(20,8) ,
27809	 => std_logic_vector(to_unsigned(62,8) ,
27810	 => std_logic_vector(to_unsigned(22,8) ,
27811	 => std_logic_vector(to_unsigned(17,8) ,
27812	 => std_logic_vector(to_unsigned(54,8) ,
27813	 => std_logic_vector(to_unsigned(79,8) ,
27814	 => std_logic_vector(to_unsigned(16,8) ,
27815	 => std_logic_vector(to_unsigned(18,8) ,
27816	 => std_logic_vector(to_unsigned(108,8) ,
27817	 => std_logic_vector(to_unsigned(108,8) ,
27818	 => std_logic_vector(to_unsigned(84,8) ,
27819	 => std_logic_vector(to_unsigned(78,8) ,
27820	 => std_logic_vector(to_unsigned(149,8) ,
27821	 => std_logic_vector(to_unsigned(163,8) ,
27822	 => std_logic_vector(to_unsigned(154,8) ,
27823	 => std_logic_vector(to_unsigned(163,8) ,
27824	 => std_logic_vector(to_unsigned(164,8) ,
27825	 => std_logic_vector(to_unsigned(161,8) ,
27826	 => std_logic_vector(to_unsigned(159,8) ,
27827	 => std_logic_vector(to_unsigned(151,8) ,
27828	 => std_logic_vector(to_unsigned(149,8) ,
27829	 => std_logic_vector(to_unsigned(157,8) ,
27830	 => std_logic_vector(to_unsigned(163,8) ,
27831	 => std_logic_vector(to_unsigned(161,8) ,
27832	 => std_logic_vector(to_unsigned(163,8) ,
27833	 => std_logic_vector(to_unsigned(161,8) ,
27834	 => std_logic_vector(to_unsigned(157,8) ,
27835	 => std_logic_vector(to_unsigned(157,8) ,
27836	 => std_logic_vector(to_unsigned(157,8) ,
27837	 => std_logic_vector(to_unsigned(163,8) ,
27838	 => std_logic_vector(to_unsigned(166,8) ,
27839	 => std_logic_vector(to_unsigned(166,8) ,
27840	 => std_logic_vector(to_unsigned(163,8) ,
27841	 => std_logic_vector(to_unsigned(159,8) ,
27842	 => std_logic_vector(to_unsigned(161,8) ,
27843	 => std_logic_vector(to_unsigned(159,8) ,
27844	 => std_logic_vector(to_unsigned(134,8) ,
27845	 => std_logic_vector(to_unsigned(144,8) ,
27846	 => std_logic_vector(to_unsigned(154,8) ,
27847	 => std_logic_vector(to_unsigned(109,8) ,
27848	 => std_logic_vector(to_unsigned(107,8) ,
27849	 => std_logic_vector(to_unsigned(128,8) ,
27850	 => std_logic_vector(to_unsigned(146,8) ,
27851	 => std_logic_vector(to_unsigned(152,8) ,
27852	 => std_logic_vector(to_unsigned(164,8) ,
27853	 => std_logic_vector(to_unsigned(177,8) ,
27854	 => std_logic_vector(to_unsigned(186,8) ,
27855	 => std_logic_vector(to_unsigned(200,8) ,
27856	 => std_logic_vector(to_unsigned(202,8) ,
27857	 => std_logic_vector(to_unsigned(202,8) ,
27858	 => std_logic_vector(to_unsigned(198,8) ,
27859	 => std_logic_vector(to_unsigned(198,8) ,
27860	 => std_logic_vector(to_unsigned(175,8) ,
27861	 => std_logic_vector(to_unsigned(112,8) ,
27862	 => std_logic_vector(to_unsigned(87,8) ,
27863	 => std_logic_vector(to_unsigned(105,8) ,
27864	 => std_logic_vector(to_unsigned(72,8) ,
27865	 => std_logic_vector(to_unsigned(3,8) ,
27866	 => std_logic_vector(to_unsigned(0,8) ,
27867	 => std_logic_vector(to_unsigned(0,8) ,
27868	 => std_logic_vector(to_unsigned(1,8) ,
27869	 => std_logic_vector(to_unsigned(7,8) ,
27870	 => std_logic_vector(to_unsigned(5,8) ,
27871	 => std_logic_vector(to_unsigned(3,8) ,
27872	 => std_logic_vector(to_unsigned(8,8) ,
27873	 => std_logic_vector(to_unsigned(32,8) ,
27874	 => std_logic_vector(to_unsigned(36,8) ,
27875	 => std_logic_vector(to_unsigned(12,8) ,
27876	 => std_logic_vector(to_unsigned(5,8) ,
27877	 => std_logic_vector(to_unsigned(11,8) ,
27878	 => std_logic_vector(to_unsigned(18,8) ,
27879	 => std_logic_vector(to_unsigned(32,8) ,
27880	 => std_logic_vector(to_unsigned(64,8) ,
27881	 => std_logic_vector(to_unsigned(85,8) ,
27882	 => std_logic_vector(to_unsigned(38,8) ,
27883	 => std_logic_vector(to_unsigned(3,8) ,
27884	 => std_logic_vector(to_unsigned(1,8) ,
27885	 => std_logic_vector(to_unsigned(2,8) ,
27886	 => std_logic_vector(to_unsigned(2,8) ,
27887	 => std_logic_vector(to_unsigned(2,8) ,
27888	 => std_logic_vector(to_unsigned(2,8) ,
27889	 => std_logic_vector(to_unsigned(2,8) ,
27890	 => std_logic_vector(to_unsigned(1,8) ,
27891	 => std_logic_vector(to_unsigned(0,8) ,
27892	 => std_logic_vector(to_unsigned(23,8) ,
27893	 => std_logic_vector(to_unsigned(85,8) ,
27894	 => std_logic_vector(to_unsigned(99,8) ,
27895	 => std_logic_vector(to_unsigned(109,8) ,
27896	 => std_logic_vector(to_unsigned(57,8) ,
27897	 => std_logic_vector(to_unsigned(8,8) ,
27898	 => std_logic_vector(to_unsigned(16,8) ,
27899	 => std_logic_vector(to_unsigned(22,8) ,
27900	 => std_logic_vector(to_unsigned(13,8) ,
27901	 => std_logic_vector(to_unsigned(13,8) ,
27902	 => std_logic_vector(to_unsigned(17,8) ,
27903	 => std_logic_vector(to_unsigned(15,8) ,
27904	 => std_logic_vector(to_unsigned(15,8) ,
27905	 => std_logic_vector(to_unsigned(17,8) ,
27906	 => std_logic_vector(to_unsigned(16,8) ,
27907	 => std_logic_vector(to_unsigned(13,8) ,
27908	 => std_logic_vector(to_unsigned(9,8) ,
27909	 => std_logic_vector(to_unsigned(8,8) ,
27910	 => std_logic_vector(to_unsigned(8,8) ,
27911	 => std_logic_vector(to_unsigned(5,8) ,
27912	 => std_logic_vector(to_unsigned(6,8) ,
27913	 => std_logic_vector(to_unsigned(3,8) ,
27914	 => std_logic_vector(to_unsigned(4,8) ,
27915	 => std_logic_vector(to_unsigned(6,8) ,
27916	 => std_logic_vector(to_unsigned(4,8) ,
27917	 => std_logic_vector(to_unsigned(5,8) ,
27918	 => std_logic_vector(to_unsigned(7,8) ,
27919	 => std_logic_vector(to_unsigned(16,8) ,
27920	 => std_logic_vector(to_unsigned(59,8) ,
27921	 => std_logic_vector(to_unsigned(131,8) ,
27922	 => std_logic_vector(to_unsigned(111,8) ,
27923	 => std_logic_vector(to_unsigned(79,8) ,
27924	 => std_logic_vector(to_unsigned(45,8) ,
27925	 => std_logic_vector(to_unsigned(9,8) ,
27926	 => std_logic_vector(to_unsigned(3,8) ,
27927	 => std_logic_vector(to_unsigned(52,8) ,
27928	 => std_logic_vector(to_unsigned(114,8) ,
27929	 => std_logic_vector(to_unsigned(95,8) ,
27930	 => std_logic_vector(to_unsigned(32,8) ,
27931	 => std_logic_vector(to_unsigned(43,8) ,
27932	 => std_logic_vector(to_unsigned(144,8) ,
27933	 => std_logic_vector(to_unsigned(144,8) ,
27934	 => std_logic_vector(to_unsigned(154,8) ,
27935	 => std_logic_vector(to_unsigned(138,8) ,
27936	 => std_logic_vector(to_unsigned(108,8) ,
27937	 => std_logic_vector(to_unsigned(62,8) ,
27938	 => std_logic_vector(to_unsigned(35,8) ,
27939	 => std_logic_vector(to_unsigned(62,8) ,
27940	 => std_logic_vector(to_unsigned(115,8) ,
27941	 => std_logic_vector(to_unsigned(74,8) ,
27942	 => std_logic_vector(to_unsigned(31,8) ,
27943	 => std_logic_vector(to_unsigned(62,8) ,
27944	 => std_logic_vector(to_unsigned(125,8) ,
27945	 => std_logic_vector(to_unsigned(47,8) ,
27946	 => std_logic_vector(to_unsigned(66,8) ,
27947	 => std_logic_vector(to_unsigned(82,8) ,
27948	 => std_logic_vector(to_unsigned(19,8) ,
27949	 => std_logic_vector(to_unsigned(5,8) ,
27950	 => std_logic_vector(to_unsigned(23,8) ,
27951	 => std_logic_vector(to_unsigned(69,8) ,
27952	 => std_logic_vector(to_unsigned(71,8) ,
27953	 => std_logic_vector(to_unsigned(24,8) ,
27954	 => std_logic_vector(to_unsigned(3,8) ,
27955	 => std_logic_vector(to_unsigned(0,8) ,
27956	 => std_logic_vector(to_unsigned(1,8) ,
27957	 => std_logic_vector(to_unsigned(2,8) ,
27958	 => std_logic_vector(to_unsigned(2,8) ,
27959	 => std_logic_vector(to_unsigned(1,8) ,
27960	 => std_logic_vector(to_unsigned(1,8) ,
27961	 => std_logic_vector(to_unsigned(2,8) ,
27962	 => std_logic_vector(to_unsigned(2,8) ,
27963	 => std_logic_vector(to_unsigned(1,8) ,
27964	 => std_logic_vector(to_unsigned(1,8) ,
27965	 => std_logic_vector(to_unsigned(2,8) ,
27966	 => std_logic_vector(to_unsigned(3,8) ,
27967	 => std_logic_vector(to_unsigned(2,8) ,
27968	 => std_logic_vector(to_unsigned(27,8) ,
27969	 => std_logic_vector(to_unsigned(104,8) ,
27970	 => std_logic_vector(to_unsigned(52,8) ,
27971	 => std_logic_vector(to_unsigned(21,8) ,
27972	 => std_logic_vector(to_unsigned(9,8) ,
27973	 => std_logic_vector(to_unsigned(5,8) ,
27974	 => std_logic_vector(to_unsigned(1,8) ,
27975	 => std_logic_vector(to_unsigned(0,8) ,
27976	 => std_logic_vector(to_unsigned(41,8) ,
27977	 => std_logic_vector(to_unsigned(122,8) ,
27978	 => std_logic_vector(to_unsigned(86,8) ,
27979	 => std_logic_vector(to_unsigned(35,8) ,
27980	 => std_logic_vector(to_unsigned(13,8) ,
27981	 => std_logic_vector(to_unsigned(8,8) ,
27982	 => std_logic_vector(to_unsigned(3,8) ,
27983	 => std_logic_vector(to_unsigned(4,8) ,
27984	 => std_logic_vector(to_unsigned(7,8) ,
27985	 => std_logic_vector(to_unsigned(22,8) ,
27986	 => std_logic_vector(to_unsigned(34,8) ,
27987	 => std_logic_vector(to_unsigned(27,8) ,
27988	 => std_logic_vector(to_unsigned(30,8) ,
27989	 => std_logic_vector(to_unsigned(37,8) ,
27990	 => std_logic_vector(to_unsigned(14,8) ,
27991	 => std_logic_vector(to_unsigned(10,8) ,
27992	 => std_logic_vector(to_unsigned(10,8) ,
27993	 => std_logic_vector(to_unsigned(8,8) ,
27994	 => std_logic_vector(to_unsigned(13,8) ,
27995	 => std_logic_vector(to_unsigned(13,8) ,
27996	 => std_logic_vector(to_unsigned(12,8) ,
27997	 => std_logic_vector(to_unsigned(37,8) ,
27998	 => std_logic_vector(to_unsigned(46,8) ,
27999	 => std_logic_vector(to_unsigned(47,8) ,
28000	 => std_logic_vector(to_unsigned(61,8) ,
28001	 => std_logic_vector(to_unsigned(82,8) ,
28002	 => std_logic_vector(to_unsigned(27,8) ,
28003	 => std_logic_vector(to_unsigned(10,8) ,
28004	 => std_logic_vector(to_unsigned(27,8) ,
28005	 => std_logic_vector(to_unsigned(69,8) ,
28006	 => std_logic_vector(to_unsigned(88,8) ,
28007	 => std_logic_vector(to_unsigned(73,8) ,
28008	 => std_logic_vector(to_unsigned(41,8) ,
28009	 => std_logic_vector(to_unsigned(70,8) ,
28010	 => std_logic_vector(to_unsigned(10,8) ,
28011	 => std_logic_vector(to_unsigned(4,8) ,
28012	 => std_logic_vector(to_unsigned(17,8) ,
28013	 => std_logic_vector(to_unsigned(22,8) ,
28014	 => std_logic_vector(to_unsigned(24,8) ,
28015	 => std_logic_vector(to_unsigned(18,8) ,
28016	 => std_logic_vector(to_unsigned(7,8) ,
28017	 => std_logic_vector(to_unsigned(6,8) ,
28018	 => std_logic_vector(to_unsigned(10,8) ,
28019	 => std_logic_vector(to_unsigned(11,8) ,
28020	 => std_logic_vector(to_unsigned(5,8) ,
28021	 => std_logic_vector(to_unsigned(2,8) ,
28022	 => std_logic_vector(to_unsigned(3,8) ,
28023	 => std_logic_vector(to_unsigned(7,8) ,
28024	 => std_logic_vector(to_unsigned(3,8) ,
28025	 => std_logic_vector(to_unsigned(5,8) ,
28026	 => std_logic_vector(to_unsigned(27,8) ,
28027	 => std_logic_vector(to_unsigned(121,8) ,
28028	 => std_logic_vector(to_unsigned(144,8) ,
28029	 => std_logic_vector(to_unsigned(122,8) ,
28030	 => std_logic_vector(to_unsigned(115,8) ,
28031	 => std_logic_vector(to_unsigned(104,8) ,
28032	 => std_logic_vector(to_unsigned(128,8) ,
28033	 => std_logic_vector(to_unsigned(152,8) ,
28034	 => std_logic_vector(to_unsigned(149,8) ,
28035	 => std_logic_vector(to_unsigned(147,8) ,
28036	 => std_logic_vector(to_unsigned(133,8) ,
28037	 => std_logic_vector(to_unsigned(144,8) ,
28038	 => std_logic_vector(to_unsigned(159,8) ,
28039	 => std_logic_vector(to_unsigned(22,8) ,
28040	 => std_logic_vector(to_unsigned(25,8) ,
28041	 => std_logic_vector(to_unsigned(152,8) ,
28042	 => std_logic_vector(to_unsigned(146,8) ,
28043	 => std_logic_vector(to_unsigned(142,8) ,
28044	 => std_logic_vector(to_unsigned(154,8) ,
28045	 => std_logic_vector(to_unsigned(149,8) ,
28046	 => std_logic_vector(to_unsigned(154,8) ,
28047	 => std_logic_vector(to_unsigned(121,8) ,
28048	 => std_logic_vector(to_unsigned(66,8) ,
28049	 => std_logic_vector(to_unsigned(92,8) ,
28050	 => std_logic_vector(to_unsigned(139,8) ,
28051	 => std_logic_vector(to_unsigned(151,8) ,
28052	 => std_logic_vector(to_unsigned(151,8) ,
28053	 => std_logic_vector(to_unsigned(141,8) ,
28054	 => std_logic_vector(to_unsigned(133,8) ,
28055	 => std_logic_vector(to_unsigned(122,8) ,
28056	 => std_logic_vector(to_unsigned(122,8) ,
28057	 => std_logic_vector(to_unsigned(156,8) ,
28058	 => std_logic_vector(to_unsigned(86,8) ,
28059	 => std_logic_vector(to_unsigned(8,8) ,
28060	 => std_logic_vector(to_unsigned(8,8) ,
28061	 => std_logic_vector(to_unsigned(9,8) ,
28062	 => std_logic_vector(to_unsigned(4,8) ,
28063	 => std_logic_vector(to_unsigned(59,8) ,
28064	 => std_logic_vector(to_unsigned(163,8) ,
28065	 => std_logic_vector(to_unsigned(161,8) ,
28066	 => std_logic_vector(to_unsigned(95,8) ,
28067	 => std_logic_vector(to_unsigned(13,8) ,
28068	 => std_logic_vector(to_unsigned(6,8) ,
28069	 => std_logic_vector(to_unsigned(12,8) ,
28070	 => std_logic_vector(to_unsigned(25,8) ,
28071	 => std_logic_vector(to_unsigned(73,8) ,
28072	 => std_logic_vector(to_unsigned(156,8) ,
28073	 => std_logic_vector(to_unsigned(168,8) ,
28074	 => std_logic_vector(to_unsigned(152,8) ,
28075	 => std_logic_vector(to_unsigned(33,8) ,
28076	 => std_logic_vector(to_unsigned(13,8) ,
28077	 => std_logic_vector(to_unsigned(28,8) ,
28078	 => std_logic_vector(to_unsigned(35,8) ,
28079	 => std_logic_vector(to_unsigned(27,8) ,
28080	 => std_logic_vector(to_unsigned(10,8) ,
28081	 => std_logic_vector(to_unsigned(4,8) ,
28082	 => std_logic_vector(to_unsigned(4,8) ,
28083	 => std_logic_vector(to_unsigned(7,8) ,
28084	 => std_logic_vector(to_unsigned(9,8) ,
28085	 => std_logic_vector(to_unsigned(7,8) ,
28086	 => std_logic_vector(to_unsigned(5,8) ,
28087	 => std_logic_vector(to_unsigned(5,8) ,
28088	 => std_logic_vector(to_unsigned(0,8) ,
28089	 => std_logic_vector(to_unsigned(5,8) ,
28090	 => std_logic_vector(to_unsigned(41,8) ,
28091	 => std_logic_vector(to_unsigned(31,8) ,
28092	 => std_logic_vector(to_unsigned(23,8) ,
28093	 => std_logic_vector(to_unsigned(17,8) ,
28094	 => std_logic_vector(to_unsigned(24,8) ,
28095	 => std_logic_vector(to_unsigned(20,8) ,
28096	 => std_logic_vector(to_unsigned(10,8) ,
28097	 => std_logic_vector(to_unsigned(12,8) ,
28098	 => std_logic_vector(to_unsigned(10,8) ,
28099	 => std_logic_vector(to_unsigned(8,8) ,
28100	 => std_logic_vector(to_unsigned(20,8) ,
28101	 => std_logic_vector(to_unsigned(10,8) ,
28102	 => std_logic_vector(to_unsigned(23,8) ,
28103	 => std_logic_vector(to_unsigned(64,8) ,
28104	 => std_logic_vector(to_unsigned(43,8) ,
28105	 => std_logic_vector(to_unsigned(32,8) ,
28106	 => std_logic_vector(to_unsigned(39,8) ,
28107	 => std_logic_vector(to_unsigned(59,8) ,
28108	 => std_logic_vector(to_unsigned(60,8) ,
28109	 => std_logic_vector(to_unsigned(42,8) ,
28110	 => std_logic_vector(to_unsigned(14,8) ,
28111	 => std_logic_vector(to_unsigned(40,8) ,
28112	 => std_logic_vector(to_unsigned(47,8) ,
28113	 => std_logic_vector(to_unsigned(16,8) ,
28114	 => std_logic_vector(to_unsigned(13,8) ,
28115	 => std_logic_vector(to_unsigned(2,8) ,
28116	 => std_logic_vector(to_unsigned(5,8) ,
28117	 => std_logic_vector(to_unsigned(3,8) ,
28118	 => std_logic_vector(to_unsigned(2,8) ,
28119	 => std_logic_vector(to_unsigned(2,8) ,
28120	 => std_logic_vector(to_unsigned(2,8) ,
28121	 => std_logic_vector(to_unsigned(3,8) ,
28122	 => std_logic_vector(to_unsigned(2,8) ,
28123	 => std_logic_vector(to_unsigned(2,8) ,
28124	 => std_logic_vector(to_unsigned(2,8) ,
28125	 => std_logic_vector(to_unsigned(3,8) ,
28126	 => std_logic_vector(to_unsigned(4,8) ,
28127	 => std_logic_vector(to_unsigned(1,8) ,
28128	 => std_logic_vector(to_unsigned(19,8) ,
28129	 => std_logic_vector(to_unsigned(56,8) ,
28130	 => std_logic_vector(to_unsigned(16,8) ,
28131	 => std_logic_vector(to_unsigned(7,8) ,
28132	 => std_logic_vector(to_unsigned(14,8) ,
28133	 => std_logic_vector(to_unsigned(17,8) ,
28134	 => std_logic_vector(to_unsigned(7,8) ,
28135	 => std_logic_vector(to_unsigned(48,8) ,
28136	 => std_logic_vector(to_unsigned(107,8) ,
28137	 => std_logic_vector(to_unsigned(93,8) ,
28138	 => std_logic_vector(to_unsigned(116,8) ,
28139	 => std_logic_vector(to_unsigned(111,8) ,
28140	 => std_logic_vector(to_unsigned(144,8) ,
28141	 => std_logic_vector(to_unsigned(163,8) ,
28142	 => std_logic_vector(to_unsigned(159,8) ,
28143	 => std_logic_vector(to_unsigned(163,8) ,
28144	 => std_logic_vector(to_unsigned(163,8) ,
28145	 => std_logic_vector(to_unsigned(147,8) ,
28146	 => std_logic_vector(to_unsigned(146,8) ,
28147	 => std_logic_vector(to_unsigned(151,8) ,
28148	 => std_logic_vector(to_unsigned(149,8) ,
28149	 => std_logic_vector(to_unsigned(161,8) ,
28150	 => std_logic_vector(to_unsigned(168,8) ,
28151	 => std_logic_vector(to_unsigned(166,8) ,
28152	 => std_logic_vector(to_unsigned(166,8) ,
28153	 => std_logic_vector(to_unsigned(166,8) ,
28154	 => std_logic_vector(to_unsigned(164,8) ,
28155	 => std_logic_vector(to_unsigned(168,8) ,
28156	 => std_logic_vector(to_unsigned(166,8) ,
28157	 => std_logic_vector(to_unsigned(163,8) ,
28158	 => std_logic_vector(to_unsigned(166,8) ,
28159	 => std_logic_vector(to_unsigned(168,8) ,
28160	 => std_logic_vector(to_unsigned(163,8) ,
28161	 => std_logic_vector(to_unsigned(163,8) ,
28162	 => std_logic_vector(to_unsigned(163,8) ,
28163	 => std_logic_vector(to_unsigned(157,8) ,
28164	 => std_logic_vector(to_unsigned(159,8) ,
28165	 => std_logic_vector(to_unsigned(164,8) ,
28166	 => std_logic_vector(to_unsigned(164,8) ,
28167	 => std_logic_vector(to_unsigned(84,8) ,
28168	 => std_logic_vector(to_unsigned(20,8) ,
28169	 => std_logic_vector(to_unsigned(24,8) ,
28170	 => std_logic_vector(to_unsigned(37,8) ,
28171	 => std_logic_vector(to_unsigned(48,8) ,
28172	 => std_logic_vector(to_unsigned(61,8) ,
28173	 => std_logic_vector(to_unsigned(68,8) ,
28174	 => std_logic_vector(to_unsigned(65,8) ,
28175	 => std_logic_vector(to_unsigned(73,8) ,
28176	 => std_logic_vector(to_unsigned(88,8) ,
28177	 => std_logic_vector(to_unsigned(114,8) ,
28178	 => std_logic_vector(to_unsigned(116,8) ,
28179	 => std_logic_vector(to_unsigned(128,8) ,
28180	 => std_logic_vector(to_unsigned(141,8) ,
28181	 => std_logic_vector(to_unsigned(100,8) ,
28182	 => std_logic_vector(to_unsigned(73,8) ,
28183	 => std_logic_vector(to_unsigned(88,8) ,
28184	 => std_logic_vector(to_unsigned(91,8) ,
28185	 => std_logic_vector(to_unsigned(8,8) ,
28186	 => std_logic_vector(to_unsigned(0,8) ,
28187	 => std_logic_vector(to_unsigned(3,8) ,
28188	 => std_logic_vector(to_unsigned(17,8) ,
28189	 => std_logic_vector(to_unsigned(13,8) ,
28190	 => std_logic_vector(to_unsigned(5,8) ,
28191	 => std_logic_vector(to_unsigned(3,8) ,
28192	 => std_logic_vector(to_unsigned(7,8) ,
28193	 => std_logic_vector(to_unsigned(33,8) ,
28194	 => std_logic_vector(to_unsigned(51,8) ,
28195	 => std_logic_vector(to_unsigned(45,8) ,
28196	 => std_logic_vector(to_unsigned(23,8) ,
28197	 => std_logic_vector(to_unsigned(12,8) ,
28198	 => std_logic_vector(to_unsigned(16,8) ,
28199	 => std_logic_vector(to_unsigned(29,8) ,
28200	 => std_logic_vector(to_unsigned(47,8) ,
28201	 => std_logic_vector(to_unsigned(46,8) ,
28202	 => std_logic_vector(to_unsigned(9,8) ,
28203	 => std_logic_vector(to_unsigned(0,8) ,
28204	 => std_logic_vector(to_unsigned(0,8) ,
28205	 => std_logic_vector(to_unsigned(0,8) ,
28206	 => std_logic_vector(to_unsigned(0,8) ,
28207	 => std_logic_vector(to_unsigned(0,8) ,
28208	 => std_logic_vector(to_unsigned(0,8) ,
28209	 => std_logic_vector(to_unsigned(0,8) ,
28210	 => std_logic_vector(to_unsigned(2,8) ,
28211	 => std_logic_vector(to_unsigned(1,8) ,
28212	 => std_logic_vector(to_unsigned(17,8) ,
28213	 => std_logic_vector(to_unsigned(87,8) ,
28214	 => std_logic_vector(to_unsigned(118,8) ,
28215	 => std_logic_vector(to_unsigned(109,8) ,
28216	 => std_logic_vector(to_unsigned(51,8) ,
28217	 => std_logic_vector(to_unsigned(5,8) ,
28218	 => std_logic_vector(to_unsigned(5,8) ,
28219	 => std_logic_vector(to_unsigned(5,8) ,
28220	 => std_logic_vector(to_unsigned(1,8) ,
28221	 => std_logic_vector(to_unsigned(1,8) ,
28222	 => std_logic_vector(to_unsigned(3,8) ,
28223	 => std_logic_vector(to_unsigned(6,8) ,
28224	 => std_logic_vector(to_unsigned(10,8) ,
28225	 => std_logic_vector(to_unsigned(16,8) ,
28226	 => std_logic_vector(to_unsigned(12,8) ,
28227	 => std_logic_vector(to_unsigned(7,8) ,
28228	 => std_logic_vector(to_unsigned(3,8) ,
28229	 => std_logic_vector(to_unsigned(3,8) ,
28230	 => std_logic_vector(to_unsigned(2,8) ,
28231	 => std_logic_vector(to_unsigned(2,8) ,
28232	 => std_logic_vector(to_unsigned(2,8) ,
28233	 => std_logic_vector(to_unsigned(3,8) ,
28234	 => std_logic_vector(to_unsigned(6,8) ,
28235	 => std_logic_vector(to_unsigned(4,8) ,
28236	 => std_logic_vector(to_unsigned(3,8) ,
28237	 => std_logic_vector(to_unsigned(6,8) ,
28238	 => std_logic_vector(to_unsigned(37,8) ,
28239	 => std_logic_vector(to_unsigned(68,8) ,
28240	 => std_logic_vector(to_unsigned(35,8) ,
28241	 => std_logic_vector(to_unsigned(33,8) ,
28242	 => std_logic_vector(to_unsigned(79,8) ,
28243	 => std_logic_vector(to_unsigned(68,8) ,
28244	 => std_logic_vector(to_unsigned(15,8) ,
28245	 => std_logic_vector(to_unsigned(8,8) ,
28246	 => std_logic_vector(to_unsigned(25,8) ,
28247	 => std_logic_vector(to_unsigned(68,8) ,
28248	 => std_logic_vector(to_unsigned(69,8) ,
28249	 => std_logic_vector(to_unsigned(35,8) ,
28250	 => std_logic_vector(to_unsigned(18,8) ,
28251	 => std_logic_vector(to_unsigned(24,8) ,
28252	 => std_logic_vector(to_unsigned(103,8) ,
28253	 => std_logic_vector(to_unsigned(136,8) ,
28254	 => std_logic_vector(to_unsigned(125,8) ,
28255	 => std_logic_vector(to_unsigned(125,8) ,
28256	 => std_logic_vector(to_unsigned(130,8) ,
28257	 => std_logic_vector(to_unsigned(118,8) ,
28258	 => std_logic_vector(to_unsigned(67,8) ,
28259	 => std_logic_vector(to_unsigned(78,8) ,
28260	 => std_logic_vector(to_unsigned(99,8) ,
28261	 => std_logic_vector(to_unsigned(82,8) ,
28262	 => std_logic_vector(to_unsigned(81,8) ,
28263	 => std_logic_vector(to_unsigned(81,8) ,
28264	 => std_logic_vector(to_unsigned(82,8) ,
28265	 => std_logic_vector(to_unsigned(28,8) ,
28266	 => std_logic_vector(to_unsigned(17,8) ,
28267	 => std_logic_vector(to_unsigned(3,8) ,
28268	 => std_logic_vector(to_unsigned(6,8) ,
28269	 => std_logic_vector(to_unsigned(12,8) ,
28270	 => std_logic_vector(to_unsigned(4,8) ,
28271	 => std_logic_vector(to_unsigned(13,8) ,
28272	 => std_logic_vector(to_unsigned(39,8) ,
28273	 => std_logic_vector(to_unsigned(19,8) ,
28274	 => std_logic_vector(to_unsigned(1,8) ,
28275	 => std_logic_vector(to_unsigned(0,8) ,
28276	 => std_logic_vector(to_unsigned(1,8) ,
28277	 => std_logic_vector(to_unsigned(2,8) ,
28278	 => std_logic_vector(to_unsigned(2,8) ,
28279	 => std_logic_vector(to_unsigned(1,8) ,
28280	 => std_logic_vector(to_unsigned(1,8) ,
28281	 => std_logic_vector(to_unsigned(1,8) ,
28282	 => std_logic_vector(to_unsigned(2,8) ,
28283	 => std_logic_vector(to_unsigned(1,8) ,
28284	 => std_logic_vector(to_unsigned(1,8) ,
28285	 => std_logic_vector(to_unsigned(1,8) ,
28286	 => std_logic_vector(to_unsigned(2,8) ,
28287	 => std_logic_vector(to_unsigned(2,8) ,
28288	 => std_logic_vector(to_unsigned(16,8) ,
28289	 => std_logic_vector(to_unsigned(19,8) ,
28290	 => std_logic_vector(to_unsigned(6,8) ,
28291	 => std_logic_vector(to_unsigned(13,8) ,
28292	 => std_logic_vector(to_unsigned(11,8) ,
28293	 => std_logic_vector(to_unsigned(5,8) ,
28294	 => std_logic_vector(to_unsigned(3,8) ,
28295	 => std_logic_vector(to_unsigned(12,8) ,
28296	 => std_logic_vector(to_unsigned(92,8) ,
28297	 => std_logic_vector(to_unsigned(108,8) ,
28298	 => std_logic_vector(to_unsigned(68,8) ,
28299	 => std_logic_vector(to_unsigned(33,8) ,
28300	 => std_logic_vector(to_unsigned(12,8) ,
28301	 => std_logic_vector(to_unsigned(5,8) ,
28302	 => std_logic_vector(to_unsigned(2,8) ,
28303	 => std_logic_vector(to_unsigned(4,8) ,
28304	 => std_logic_vector(to_unsigned(8,8) ,
28305	 => std_logic_vector(to_unsigned(17,8) ,
28306	 => std_logic_vector(to_unsigned(19,8) ,
28307	 => std_logic_vector(to_unsigned(17,8) ,
28308	 => std_logic_vector(to_unsigned(24,8) ,
28309	 => std_logic_vector(to_unsigned(30,8) ,
28310	 => std_logic_vector(to_unsigned(16,8) ,
28311	 => std_logic_vector(to_unsigned(13,8) ,
28312	 => std_logic_vector(to_unsigned(13,8) ,
28313	 => std_logic_vector(to_unsigned(9,8) ,
28314	 => std_logic_vector(to_unsigned(15,8) ,
28315	 => std_logic_vector(to_unsigned(12,8) ,
28316	 => std_logic_vector(to_unsigned(9,8) ,
28317	 => std_logic_vector(to_unsigned(50,8) ,
28318	 => std_logic_vector(to_unsigned(65,8) ,
28319	 => std_logic_vector(to_unsigned(45,8) ,
28320	 => std_logic_vector(to_unsigned(76,8) ,
28321	 => std_logic_vector(to_unsigned(108,8) ,
28322	 => std_logic_vector(to_unsigned(27,8) ,
28323	 => std_logic_vector(to_unsigned(8,8) ,
28324	 => std_logic_vector(to_unsigned(33,8) ,
28325	 => std_logic_vector(to_unsigned(74,8) ,
28326	 => std_logic_vector(to_unsigned(86,8) ,
28327	 => std_logic_vector(to_unsigned(63,8) ,
28328	 => std_logic_vector(to_unsigned(35,8) ,
28329	 => std_logic_vector(to_unsigned(133,8) ,
28330	 => std_logic_vector(to_unsigned(64,8) ,
28331	 => std_logic_vector(to_unsigned(3,8) ,
28332	 => std_logic_vector(to_unsigned(12,8) ,
28333	 => std_logic_vector(to_unsigned(19,8) ,
28334	 => std_logic_vector(to_unsigned(19,8) ,
28335	 => std_logic_vector(to_unsigned(18,8) ,
28336	 => std_logic_vector(to_unsigned(9,8) ,
28337	 => std_logic_vector(to_unsigned(6,8) ,
28338	 => std_logic_vector(to_unsigned(5,8) ,
28339	 => std_logic_vector(to_unsigned(5,8) ,
28340	 => std_logic_vector(to_unsigned(2,8) ,
28341	 => std_logic_vector(to_unsigned(2,8) ,
28342	 => std_logic_vector(to_unsigned(8,8) ,
28343	 => std_logic_vector(to_unsigned(9,8) ,
28344	 => std_logic_vector(to_unsigned(3,8) ,
28345	 => std_logic_vector(to_unsigned(2,8) ,
28346	 => std_logic_vector(to_unsigned(21,8) ,
28347	 => std_logic_vector(to_unsigned(134,8) ,
28348	 => std_logic_vector(to_unsigned(149,8) ,
28349	 => std_logic_vector(to_unsigned(146,8) ,
28350	 => std_logic_vector(to_unsigned(127,8) ,
28351	 => std_logic_vector(to_unsigned(104,8) ,
28352	 => std_logic_vector(to_unsigned(116,8) ,
28353	 => std_logic_vector(to_unsigned(152,8) ,
28354	 => std_logic_vector(to_unsigned(151,8) ,
28355	 => std_logic_vector(to_unsigned(154,8) ,
28356	 => std_logic_vector(to_unsigned(146,8) ,
28357	 => std_logic_vector(to_unsigned(136,8) ,
28358	 => std_logic_vector(to_unsigned(164,8) ,
28359	 => std_logic_vector(to_unsigned(87,8) ,
28360	 => std_logic_vector(to_unsigned(88,8) ,
28361	 => std_logic_vector(to_unsigned(170,8) ,
28362	 => std_logic_vector(to_unsigned(139,8) ,
28363	 => std_logic_vector(to_unsigned(147,8) ,
28364	 => std_logic_vector(to_unsigned(154,8) ,
28365	 => std_logic_vector(to_unsigned(154,8) ,
28366	 => std_logic_vector(to_unsigned(154,8) ,
28367	 => std_logic_vector(to_unsigned(92,8) ,
28368	 => std_logic_vector(to_unsigned(62,8) ,
28369	 => std_logic_vector(to_unsigned(127,8) ,
28370	 => std_logic_vector(to_unsigned(152,8) ,
28371	 => std_logic_vector(to_unsigned(154,8) ,
28372	 => std_logic_vector(to_unsigned(157,8) ,
28373	 => std_logic_vector(to_unsigned(139,8) ,
28374	 => std_logic_vector(to_unsigned(130,8) ,
28375	 => std_logic_vector(to_unsigned(128,8) ,
28376	 => std_logic_vector(to_unsigned(133,8) ,
28377	 => std_logic_vector(to_unsigned(139,8) ,
28378	 => std_logic_vector(to_unsigned(32,8) ,
28379	 => std_logic_vector(to_unsigned(5,8) ,
28380	 => std_logic_vector(to_unsigned(8,8) ,
28381	 => std_logic_vector(to_unsigned(8,8) ,
28382	 => std_logic_vector(to_unsigned(4,8) ,
28383	 => std_logic_vector(to_unsigned(82,8) ,
28384	 => std_logic_vector(to_unsigned(166,8) ,
28385	 => std_logic_vector(to_unsigned(144,8) ,
28386	 => std_logic_vector(to_unsigned(168,8) ,
28387	 => std_logic_vector(to_unsigned(104,8) ,
28388	 => std_logic_vector(to_unsigned(35,8) ,
28389	 => std_logic_vector(to_unsigned(36,8) ,
28390	 => std_logic_vector(to_unsigned(87,8) ,
28391	 => std_logic_vector(to_unsigned(157,8) ,
28392	 => std_logic_vector(to_unsigned(157,8) ,
28393	 => std_logic_vector(to_unsigned(168,8) ,
28394	 => std_logic_vector(to_unsigned(125,8) ,
28395	 => std_logic_vector(to_unsigned(17,8) ,
28396	 => std_logic_vector(to_unsigned(16,8) ,
28397	 => std_logic_vector(to_unsigned(35,8) ,
28398	 => std_logic_vector(to_unsigned(42,8) ,
28399	 => std_logic_vector(to_unsigned(32,8) ,
28400	 => std_logic_vector(to_unsigned(8,8) ,
28401	 => std_logic_vector(to_unsigned(5,8) ,
28402	 => std_logic_vector(to_unsigned(9,8) ,
28403	 => std_logic_vector(to_unsigned(5,8) ,
28404	 => std_logic_vector(to_unsigned(10,8) ,
28405	 => std_logic_vector(to_unsigned(10,8) ,
28406	 => std_logic_vector(to_unsigned(8,8) ,
28407	 => std_logic_vector(to_unsigned(7,8) ,
28408	 => std_logic_vector(to_unsigned(3,8) ,
28409	 => std_logic_vector(to_unsigned(1,8) ,
28410	 => std_logic_vector(to_unsigned(8,8) ,
28411	 => std_logic_vector(to_unsigned(40,8) ,
28412	 => std_logic_vector(to_unsigned(24,8) ,
28413	 => std_logic_vector(to_unsigned(20,8) ,
28414	 => std_logic_vector(to_unsigned(30,8) ,
28415	 => std_logic_vector(to_unsigned(24,8) ,
28416	 => std_logic_vector(to_unsigned(13,8) ,
28417	 => std_logic_vector(to_unsigned(17,8) ,
28418	 => std_logic_vector(to_unsigned(15,8) ,
28419	 => std_logic_vector(to_unsigned(7,8) ,
28420	 => std_logic_vector(to_unsigned(13,8) ,
28421	 => std_logic_vector(to_unsigned(63,8) ,
28422	 => std_logic_vector(to_unsigned(114,8) ,
28423	 => std_logic_vector(to_unsigned(44,8) ,
28424	 => std_logic_vector(to_unsigned(27,8) ,
28425	 => std_logic_vector(to_unsigned(29,8) ,
28426	 => std_logic_vector(to_unsigned(29,8) ,
28427	 => std_logic_vector(to_unsigned(60,8) ,
28428	 => std_logic_vector(to_unsigned(59,8) ,
28429	 => std_logic_vector(to_unsigned(45,8) ,
28430	 => std_logic_vector(to_unsigned(31,8) ,
28431	 => std_logic_vector(to_unsigned(22,8) ,
28432	 => std_logic_vector(to_unsigned(93,8) ,
28433	 => std_logic_vector(to_unsigned(41,8) ,
28434	 => std_logic_vector(to_unsigned(5,8) ,
28435	 => std_logic_vector(to_unsigned(4,8) ,
28436	 => std_logic_vector(to_unsigned(5,8) ,
28437	 => std_logic_vector(to_unsigned(4,8) ,
28438	 => std_logic_vector(to_unsigned(4,8) ,
28439	 => std_logic_vector(to_unsigned(4,8) ,
28440	 => std_logic_vector(to_unsigned(4,8) ,
28441	 => std_logic_vector(to_unsigned(3,8) ,
28442	 => std_logic_vector(to_unsigned(2,8) ,
28443	 => std_logic_vector(to_unsigned(2,8) ,
28444	 => std_logic_vector(to_unsigned(2,8) ,
28445	 => std_logic_vector(to_unsigned(4,8) ,
28446	 => std_logic_vector(to_unsigned(4,8) ,
28447	 => std_logic_vector(to_unsigned(1,8) ,
28448	 => std_logic_vector(to_unsigned(13,8) ,
28449	 => std_logic_vector(to_unsigned(51,8) ,
28450	 => std_logic_vector(to_unsigned(16,8) ,
28451	 => std_logic_vector(to_unsigned(6,8) ,
28452	 => std_logic_vector(to_unsigned(6,8) ,
28453	 => std_logic_vector(to_unsigned(4,8) ,
28454	 => std_logic_vector(to_unsigned(18,8) ,
28455	 => std_logic_vector(to_unsigned(93,8) ,
28456	 => std_logic_vector(to_unsigned(100,8) ,
28457	 => std_logic_vector(to_unsigned(96,8) ,
28458	 => std_logic_vector(to_unsigned(131,8) ,
28459	 => std_logic_vector(to_unsigned(139,8) ,
28460	 => std_logic_vector(to_unsigned(151,8) ,
28461	 => std_logic_vector(to_unsigned(152,8) ,
28462	 => std_logic_vector(to_unsigned(142,8) ,
28463	 => std_logic_vector(to_unsigned(156,8) ,
28464	 => std_logic_vector(to_unsigned(163,8) ,
28465	 => std_logic_vector(to_unsigned(138,8) ,
28466	 => std_logic_vector(to_unsigned(142,8) ,
28467	 => std_logic_vector(to_unsigned(149,8) ,
28468	 => std_logic_vector(to_unsigned(154,8) ,
28469	 => std_logic_vector(to_unsigned(163,8) ,
28470	 => std_logic_vector(to_unsigned(166,8) ,
28471	 => std_logic_vector(to_unsigned(166,8) ,
28472	 => std_logic_vector(to_unsigned(168,8) ,
28473	 => std_logic_vector(to_unsigned(171,8) ,
28474	 => std_logic_vector(to_unsigned(173,8) ,
28475	 => std_logic_vector(to_unsigned(173,8) ,
28476	 => std_logic_vector(to_unsigned(175,8) ,
28477	 => std_logic_vector(to_unsigned(175,8) ,
28478	 => std_logic_vector(to_unsigned(166,8) ,
28479	 => std_logic_vector(to_unsigned(157,8) ,
28480	 => std_logic_vector(to_unsigned(156,8) ,
28481	 => std_logic_vector(to_unsigned(154,8) ,
28482	 => std_logic_vector(to_unsigned(147,8) ,
28483	 => std_logic_vector(to_unsigned(144,8) ,
28484	 => std_logic_vector(to_unsigned(151,8) ,
28485	 => std_logic_vector(to_unsigned(146,8) ,
28486	 => std_logic_vector(to_unsigned(151,8) ,
28487	 => std_logic_vector(to_unsigned(159,8) ,
28488	 => std_logic_vector(to_unsigned(70,8) ,
28489	 => std_logic_vector(to_unsigned(26,8) ,
28490	 => std_logic_vector(to_unsigned(32,8) ,
28491	 => std_logic_vector(to_unsigned(37,8) ,
28492	 => std_logic_vector(to_unsigned(43,8) ,
28493	 => std_logic_vector(to_unsigned(35,8) ,
28494	 => std_logic_vector(to_unsigned(24,8) ,
28495	 => std_logic_vector(to_unsigned(25,8) ,
28496	 => std_logic_vector(to_unsigned(29,8) ,
28497	 => std_logic_vector(to_unsigned(35,8) ,
28498	 => std_logic_vector(to_unsigned(29,8) ,
28499	 => std_logic_vector(to_unsigned(35,8) ,
28500	 => std_logic_vector(to_unsigned(36,8) ,
28501	 => std_logic_vector(to_unsigned(44,8) ,
28502	 => std_logic_vector(to_unsigned(82,8) ,
28503	 => std_logic_vector(to_unsigned(86,8) ,
28504	 => std_logic_vector(to_unsigned(78,8) ,
28505	 => std_logic_vector(to_unsigned(22,8) ,
28506	 => std_logic_vector(to_unsigned(13,8) ,
28507	 => std_logic_vector(to_unsigned(37,8) ,
28508	 => std_logic_vector(to_unsigned(18,8) ,
28509	 => std_logic_vector(to_unsigned(7,8) ,
28510	 => std_logic_vector(to_unsigned(3,8) ,
28511	 => std_logic_vector(to_unsigned(1,8) ,
28512	 => std_logic_vector(to_unsigned(2,8) ,
28513	 => std_logic_vector(to_unsigned(20,8) ,
28514	 => std_logic_vector(to_unsigned(39,8) ,
28515	 => std_logic_vector(to_unsigned(60,8) ,
28516	 => std_logic_vector(to_unsigned(70,8) ,
28517	 => std_logic_vector(to_unsigned(53,8) ,
28518	 => std_logic_vector(to_unsigned(20,8) ,
28519	 => std_logic_vector(to_unsigned(17,8) ,
28520	 => std_logic_vector(to_unsigned(6,8) ,
28521	 => std_logic_vector(to_unsigned(5,8) ,
28522	 => std_logic_vector(to_unsigned(7,8) ,
28523	 => std_logic_vector(to_unsigned(6,8) ,
28524	 => std_logic_vector(to_unsigned(5,8) ,
28525	 => std_logic_vector(to_unsigned(3,8) ,
28526	 => std_logic_vector(to_unsigned(4,8) ,
28527	 => std_logic_vector(to_unsigned(8,8) ,
28528	 => std_logic_vector(to_unsigned(10,8) ,
28529	 => std_logic_vector(to_unsigned(6,8) ,
28530	 => std_logic_vector(to_unsigned(2,8) ,
28531	 => std_logic_vector(to_unsigned(2,8) ,
28532	 => std_logic_vector(to_unsigned(15,8) ,
28533	 => std_logic_vector(to_unsigned(86,8) ,
28534	 => std_logic_vector(to_unsigned(112,8) ,
28535	 => std_logic_vector(to_unsigned(111,8) ,
28536	 => std_logic_vector(to_unsigned(73,8) ,
28537	 => std_logic_vector(to_unsigned(14,8) ,
28538	 => std_logic_vector(to_unsigned(1,8) ,
28539	 => std_logic_vector(to_unsigned(0,8) ,
28540	 => std_logic_vector(to_unsigned(0,8) ,
28541	 => std_logic_vector(to_unsigned(0,8) ,
28542	 => std_logic_vector(to_unsigned(0,8) ,
28543	 => std_logic_vector(to_unsigned(1,8) ,
28544	 => std_logic_vector(to_unsigned(4,8) ,
28545	 => std_logic_vector(to_unsigned(3,8) ,
28546	 => std_logic_vector(to_unsigned(2,8) ,
28547	 => std_logic_vector(to_unsigned(0,8) ,
28548	 => std_logic_vector(to_unsigned(0,8) ,
28549	 => std_logic_vector(to_unsigned(0,8) ,
28550	 => std_logic_vector(to_unsigned(1,8) ,
28551	 => std_logic_vector(to_unsigned(1,8) ,
28552	 => std_logic_vector(to_unsigned(1,8) ,
28553	 => std_logic_vector(to_unsigned(4,8) ,
28554	 => std_logic_vector(to_unsigned(6,8) ,
28555	 => std_logic_vector(to_unsigned(9,8) ,
28556	 => std_logic_vector(to_unsigned(7,8) ,
28557	 => std_logic_vector(to_unsigned(6,8) ,
28558	 => std_logic_vector(to_unsigned(54,8) ,
28559	 => std_logic_vector(to_unsigned(128,8) ,
28560	 => std_logic_vector(to_unsigned(104,8) ,
28561	 => std_logic_vector(to_unsigned(34,8) ,
28562	 => std_logic_vector(to_unsigned(12,8) ,
28563	 => std_logic_vector(to_unsigned(14,8) ,
28564	 => std_logic_vector(to_unsigned(8,8) ,
28565	 => std_logic_vector(to_unsigned(49,8) ,
28566	 => std_logic_vector(to_unsigned(78,8) ,
28567	 => std_logic_vector(to_unsigned(61,8) ,
28568	 => std_logic_vector(to_unsigned(30,8) ,
28569	 => std_logic_vector(to_unsigned(19,8) ,
28570	 => std_logic_vector(to_unsigned(17,8) ,
28571	 => std_logic_vector(to_unsigned(11,8) ,
28572	 => std_logic_vector(to_unsigned(51,8) ,
28573	 => std_logic_vector(to_unsigned(127,8) ,
28574	 => std_logic_vector(to_unsigned(115,8) ,
28575	 => std_logic_vector(to_unsigned(107,8) ,
28576	 => std_logic_vector(to_unsigned(107,8) ,
28577	 => std_logic_vector(to_unsigned(133,8) ,
28578	 => std_logic_vector(to_unsigned(152,8) ,
28579	 => std_logic_vector(to_unsigned(105,8) ,
28580	 => std_logic_vector(to_unsigned(56,8) ,
28581	 => std_logic_vector(to_unsigned(121,8) ,
28582	 => std_logic_vector(to_unsigned(112,8) ,
28583	 => std_logic_vector(to_unsigned(49,8) ,
28584	 => std_logic_vector(to_unsigned(35,8) ,
28585	 => std_logic_vector(to_unsigned(13,8) ,
28586	 => std_logic_vector(to_unsigned(2,8) ,
28587	 => std_logic_vector(to_unsigned(4,8) ,
28588	 => std_logic_vector(to_unsigned(14,8) ,
28589	 => std_logic_vector(to_unsigned(19,8) ,
28590	 => std_logic_vector(to_unsigned(13,8) ,
28591	 => std_logic_vector(to_unsigned(5,8) ,
28592	 => std_logic_vector(to_unsigned(3,8) ,
28593	 => std_logic_vector(to_unsigned(16,8) ,
28594	 => std_logic_vector(to_unsigned(38,8) ,
28595	 => std_logic_vector(to_unsigned(6,8) ,
28596	 => std_logic_vector(to_unsigned(1,8) ,
28597	 => std_logic_vector(to_unsigned(2,8) ,
28598	 => std_logic_vector(to_unsigned(2,8) ,
28599	 => std_logic_vector(to_unsigned(2,8) ,
28600	 => std_logic_vector(to_unsigned(1,8) ,
28601	 => std_logic_vector(to_unsigned(1,8) ,
28602	 => std_logic_vector(to_unsigned(2,8) ,
28603	 => std_logic_vector(to_unsigned(2,8) ,
28604	 => std_logic_vector(to_unsigned(2,8) ,
28605	 => std_logic_vector(to_unsigned(1,8) ,
28606	 => std_logic_vector(to_unsigned(1,8) ,
28607	 => std_logic_vector(to_unsigned(1,8) ,
28608	 => std_logic_vector(to_unsigned(2,8) ,
28609	 => std_logic_vector(to_unsigned(13,8) ,
28610	 => std_logic_vector(to_unsigned(51,8) ,
28611	 => std_logic_vector(to_unsigned(57,8) ,
28612	 => std_logic_vector(to_unsigned(38,8) ,
28613	 => std_logic_vector(to_unsigned(13,8) ,
28614	 => std_logic_vector(to_unsigned(10,8) ,
28615	 => std_logic_vector(to_unsigned(67,8) ,
28616	 => std_logic_vector(to_unsigned(105,8) ,
28617	 => std_logic_vector(to_unsigned(69,8) ,
28618	 => std_logic_vector(to_unsigned(61,8) ,
28619	 => std_logic_vector(to_unsigned(44,8) ,
28620	 => std_logic_vector(to_unsigned(15,8) ,
28621	 => std_logic_vector(to_unsigned(2,8) ,
28622	 => std_logic_vector(to_unsigned(3,8) ,
28623	 => std_logic_vector(to_unsigned(4,8) ,
28624	 => std_logic_vector(to_unsigned(7,8) ,
28625	 => std_logic_vector(to_unsigned(19,8) ,
28626	 => std_logic_vector(to_unsigned(17,8) ,
28627	 => std_logic_vector(to_unsigned(17,8) ,
28628	 => std_logic_vector(to_unsigned(33,8) ,
28629	 => std_logic_vector(to_unsigned(30,8) ,
28630	 => std_logic_vector(to_unsigned(10,8) ,
28631	 => std_logic_vector(to_unsigned(12,8) ,
28632	 => std_logic_vector(to_unsigned(17,8) ,
28633	 => std_logic_vector(to_unsigned(11,8) ,
28634	 => std_logic_vector(to_unsigned(10,8) ,
28635	 => std_logic_vector(to_unsigned(7,8) ,
28636	 => std_logic_vector(to_unsigned(15,8) ,
28637	 => std_logic_vector(to_unsigned(61,8) ,
28638	 => std_logic_vector(to_unsigned(71,8) ,
28639	 => std_logic_vector(to_unsigned(69,8) ,
28640	 => std_logic_vector(to_unsigned(93,8) ,
28641	 => std_logic_vector(to_unsigned(99,8) ,
28642	 => std_logic_vector(to_unsigned(25,8) ,
28643	 => std_logic_vector(to_unsigned(10,8) ,
28644	 => std_logic_vector(to_unsigned(35,8) ,
28645	 => std_logic_vector(to_unsigned(73,8) ,
28646	 => std_logic_vector(to_unsigned(86,8) ,
28647	 => std_logic_vector(to_unsigned(55,8) ,
28648	 => std_logic_vector(to_unsigned(38,8) ,
28649	 => std_logic_vector(to_unsigned(142,8) ,
28650	 => std_logic_vector(to_unsigned(144,8) ,
28651	 => std_logic_vector(to_unsigned(9,8) ,
28652	 => std_logic_vector(to_unsigned(2,8) ,
28653	 => std_logic_vector(to_unsigned(10,8) ,
28654	 => std_logic_vector(to_unsigned(25,8) ,
28655	 => std_logic_vector(to_unsigned(24,8) ,
28656	 => std_logic_vector(to_unsigned(13,8) ,
28657	 => std_logic_vector(to_unsigned(10,8) ,
28658	 => std_logic_vector(to_unsigned(5,8) ,
28659	 => std_logic_vector(to_unsigned(4,8) ,
28660	 => std_logic_vector(to_unsigned(4,8) ,
28661	 => std_logic_vector(to_unsigned(8,8) ,
28662	 => std_logic_vector(to_unsigned(8,8) ,
28663	 => std_logic_vector(to_unsigned(5,8) ,
28664	 => std_logic_vector(to_unsigned(4,8) ,
28665	 => std_logic_vector(to_unsigned(1,8) ,
28666	 => std_logic_vector(to_unsigned(29,8) ,
28667	 => std_logic_vector(to_unsigned(159,8) ,
28668	 => std_logic_vector(to_unsigned(142,8) ,
28669	 => std_logic_vector(to_unsigned(151,8) ,
28670	 => std_logic_vector(to_unsigned(147,8) ,
28671	 => std_logic_vector(to_unsigned(130,8) ,
28672	 => std_logic_vector(to_unsigned(96,8) ,
28673	 => std_logic_vector(to_unsigned(139,8) ,
28674	 => std_logic_vector(to_unsigned(154,8) ,
28675	 => std_logic_vector(to_unsigned(156,8) ,
28676	 => std_logic_vector(to_unsigned(152,8) ,
28677	 => std_logic_vector(to_unsigned(144,8) ,
28678	 => std_logic_vector(to_unsigned(141,8) ,
28679	 => std_logic_vector(to_unsigned(141,8) ,
28680	 => std_logic_vector(to_unsigned(152,8) ,
28681	 => std_logic_vector(to_unsigned(152,8) ,
28682	 => std_logic_vector(to_unsigned(146,8) ,
28683	 => std_logic_vector(to_unsigned(154,8) ,
28684	 => std_logic_vector(to_unsigned(151,8) ,
28685	 => std_logic_vector(to_unsigned(154,8) ,
28686	 => std_logic_vector(to_unsigned(147,8) ,
28687	 => std_logic_vector(to_unsigned(104,8) ,
28688	 => std_logic_vector(to_unsigned(87,8) ,
28689	 => std_logic_vector(to_unsigned(147,8) ,
28690	 => std_logic_vector(to_unsigned(157,8) ,
28691	 => std_logic_vector(to_unsigned(156,8) ,
28692	 => std_logic_vector(to_unsigned(138,8) ,
28693	 => std_logic_vector(to_unsigned(141,8) ,
28694	 => std_logic_vector(to_unsigned(141,8) ,
28695	 => std_logic_vector(to_unsigned(122,8) ,
28696	 => std_logic_vector(to_unsigned(130,8) ,
28697	 => std_logic_vector(to_unsigned(84,8) ,
28698	 => std_logic_vector(to_unsigned(9,8) ,
28699	 => std_logic_vector(to_unsigned(6,8) ,
28700	 => std_logic_vector(to_unsigned(10,8) ,
28701	 => std_logic_vector(to_unsigned(6,8) ,
28702	 => std_logic_vector(to_unsigned(4,8) ,
28703	 => std_logic_vector(to_unsigned(99,8) ,
28704	 => std_logic_vector(to_unsigned(163,8) ,
28705	 => std_logic_vector(to_unsigned(146,8) ,
28706	 => std_logic_vector(to_unsigned(146,8) ,
28707	 => std_logic_vector(to_unsigned(156,8) ,
28708	 => std_logic_vector(to_unsigned(157,8) ,
28709	 => std_logic_vector(to_unsigned(163,8) ,
28710	 => std_logic_vector(to_unsigned(171,8) ,
28711	 => std_logic_vector(to_unsigned(157,8) ,
28712	 => std_logic_vector(to_unsigned(151,8) ,
28713	 => std_logic_vector(to_unsigned(171,8) ,
28714	 => std_logic_vector(to_unsigned(85,8) ,
28715	 => std_logic_vector(to_unsigned(8,8) ,
28716	 => std_logic_vector(to_unsigned(15,8) ,
28717	 => std_logic_vector(to_unsigned(34,8) ,
28718	 => std_logic_vector(to_unsigned(41,8) ,
28719	 => std_logic_vector(to_unsigned(27,8) ,
28720	 => std_logic_vector(to_unsigned(6,8) ,
28721	 => std_logic_vector(to_unsigned(5,8) ,
28722	 => std_logic_vector(to_unsigned(11,8) ,
28723	 => std_logic_vector(to_unsigned(7,8) ,
28724	 => std_logic_vector(to_unsigned(5,8) ,
28725	 => std_logic_vector(to_unsigned(12,8) ,
28726	 => std_logic_vector(to_unsigned(9,8) ,
28727	 => std_logic_vector(to_unsigned(7,8) ,
28728	 => std_logic_vector(to_unsigned(9,8) ,
28729	 => std_logic_vector(to_unsigned(11,8) ,
28730	 => std_logic_vector(to_unsigned(10,8) ,
28731	 => std_logic_vector(to_unsigned(10,8) ,
28732	 => std_logic_vector(to_unsigned(12,8) ,
28733	 => std_logic_vector(to_unsigned(15,8) ,
28734	 => std_logic_vector(to_unsigned(22,8) ,
28735	 => std_logic_vector(to_unsigned(19,8) ,
28736	 => std_logic_vector(to_unsigned(22,8) ,
28737	 => std_logic_vector(to_unsigned(23,8) ,
28738	 => std_logic_vector(to_unsigned(23,8) ,
28739	 => std_logic_vector(to_unsigned(10,8) ,
28740	 => std_logic_vector(to_unsigned(7,8) ,
28741	 => std_logic_vector(to_unsigned(56,8) ,
28742	 => std_logic_vector(to_unsigned(157,8) ,
28743	 => std_logic_vector(to_unsigned(87,8) ,
28744	 => std_logic_vector(to_unsigned(73,8) ,
28745	 => std_logic_vector(to_unsigned(64,8) ,
28746	 => std_logic_vector(to_unsigned(41,8) ,
28747	 => std_logic_vector(to_unsigned(76,8) ,
28748	 => std_logic_vector(to_unsigned(79,8) ,
28749	 => std_logic_vector(to_unsigned(45,8) ,
28750	 => std_logic_vector(to_unsigned(51,8) ,
28751	 => std_logic_vector(to_unsigned(32,8) ,
28752	 => std_logic_vector(to_unsigned(46,8) ,
28753	 => std_logic_vector(to_unsigned(50,8) ,
28754	 => std_logic_vector(to_unsigned(2,8) ,
28755	 => std_logic_vector(to_unsigned(4,8) ,
28756	 => std_logic_vector(to_unsigned(5,8) ,
28757	 => std_logic_vector(to_unsigned(4,8) ,
28758	 => std_logic_vector(to_unsigned(4,8) ,
28759	 => std_logic_vector(to_unsigned(4,8) ,
28760	 => std_logic_vector(to_unsigned(4,8) ,
28761	 => std_logic_vector(to_unsigned(3,8) ,
28762	 => std_logic_vector(to_unsigned(2,8) ,
28763	 => std_logic_vector(to_unsigned(1,8) ,
28764	 => std_logic_vector(to_unsigned(2,8) ,
28765	 => std_logic_vector(to_unsigned(5,8) ,
28766	 => std_logic_vector(to_unsigned(3,8) ,
28767	 => std_logic_vector(to_unsigned(1,8) ,
28768	 => std_logic_vector(to_unsigned(10,8) ,
28769	 => std_logic_vector(to_unsigned(45,8) ,
28770	 => std_logic_vector(to_unsigned(16,8) ,
28771	 => std_logic_vector(to_unsigned(7,8) ,
28772	 => std_logic_vector(to_unsigned(5,8) ,
28773	 => std_logic_vector(to_unsigned(3,8) ,
28774	 => std_logic_vector(to_unsigned(37,8) ,
28775	 => std_logic_vector(to_unsigned(73,8) ,
28776	 => std_logic_vector(to_unsigned(74,8) ,
28777	 => std_logic_vector(to_unsigned(101,8) ,
28778	 => std_logic_vector(to_unsigned(139,8) ,
28779	 => std_logic_vector(to_unsigned(159,8) ,
28780	 => std_logic_vector(to_unsigned(157,8) ,
28781	 => std_logic_vector(to_unsigned(142,8) ,
28782	 => std_logic_vector(to_unsigned(134,8) ,
28783	 => std_logic_vector(to_unsigned(147,8) ,
28784	 => std_logic_vector(to_unsigned(163,8) ,
28785	 => std_logic_vector(to_unsigned(157,8) ,
28786	 => std_logic_vector(to_unsigned(156,8) ,
28787	 => std_logic_vector(to_unsigned(163,8) ,
28788	 => std_logic_vector(to_unsigned(163,8) ,
28789	 => std_logic_vector(to_unsigned(170,8) ,
28790	 => std_logic_vector(to_unsigned(168,8) ,
28791	 => std_logic_vector(to_unsigned(166,8) ,
28792	 => std_logic_vector(to_unsigned(164,8) ,
28793	 => std_logic_vector(to_unsigned(166,8) ,
28794	 => std_logic_vector(to_unsigned(168,8) ,
28795	 => std_logic_vector(to_unsigned(163,8) ,
28796	 => std_logic_vector(to_unsigned(166,8) ,
28797	 => std_logic_vector(to_unsigned(171,8) ,
28798	 => std_logic_vector(to_unsigned(164,8) ,
28799	 => std_logic_vector(to_unsigned(157,8) ,
28800	 => std_logic_vector(to_unsigned(157,8) ,
28801	 => std_logic_vector(to_unsigned(146,8) ,
28802	 => std_logic_vector(to_unsigned(144,8) ,
28803	 => std_logic_vector(to_unsigned(144,8) ,
28804	 => std_logic_vector(to_unsigned(134,8) ,
28805	 => std_logic_vector(to_unsigned(130,8) ,
28806	 => std_logic_vector(to_unsigned(131,8) ,
28807	 => std_logic_vector(to_unsigned(146,8) ,
28808	 => std_logic_vector(to_unsigned(115,8) ,
28809	 => std_logic_vector(to_unsigned(88,8) ,
28810	 => std_logic_vector(to_unsigned(104,8) ,
28811	 => std_logic_vector(to_unsigned(96,8) ,
28812	 => std_logic_vector(to_unsigned(87,8) ,
28813	 => std_logic_vector(to_unsigned(73,8) ,
28814	 => std_logic_vector(to_unsigned(61,8) ,
28815	 => std_logic_vector(to_unsigned(62,8) ,
28816	 => std_logic_vector(to_unsigned(59,8) ,
28817	 => std_logic_vector(to_unsigned(54,8) ,
28818	 => std_logic_vector(to_unsigned(47,8) ,
28819	 => std_logic_vector(to_unsigned(35,8) ,
28820	 => std_logic_vector(to_unsigned(17,8) ,
28821	 => std_logic_vector(to_unsigned(23,8) ,
28822	 => std_logic_vector(to_unsigned(69,8) ,
28823	 => std_logic_vector(to_unsigned(70,8) ,
28824	 => std_logic_vector(to_unsigned(65,8) ,
28825	 => std_logic_vector(to_unsigned(41,8) ,
28826	 => std_logic_vector(to_unsigned(39,8) ,
28827	 => std_logic_vector(to_unsigned(29,8) ,
28828	 => std_logic_vector(to_unsigned(6,8) ,
28829	 => std_logic_vector(to_unsigned(3,8) ,
28830	 => std_logic_vector(to_unsigned(2,8) ,
28831	 => std_logic_vector(to_unsigned(0,8) ,
28832	 => std_logic_vector(to_unsigned(1,8) ,
28833	 => std_logic_vector(to_unsigned(9,8) ,
28834	 => std_logic_vector(to_unsigned(15,8) ,
28835	 => std_logic_vector(to_unsigned(41,8) ,
28836	 => std_logic_vector(to_unsigned(70,8) ,
28837	 => std_logic_vector(to_unsigned(61,8) ,
28838	 => std_logic_vector(to_unsigned(52,8) ,
28839	 => std_logic_vector(to_unsigned(56,8) ,
28840	 => std_logic_vector(to_unsigned(41,8) ,
28841	 => std_logic_vector(to_unsigned(45,8) ,
28842	 => std_logic_vector(to_unsigned(51,8) ,
28843	 => std_logic_vector(to_unsigned(66,8) ,
28844	 => std_logic_vector(to_unsigned(91,8) ,
28845	 => std_logic_vector(to_unsigned(99,8) ,
28846	 => std_logic_vector(to_unsigned(121,8) ,
28847	 => std_logic_vector(to_unsigned(139,8) ,
28848	 => std_logic_vector(to_unsigned(147,8) ,
28849	 => std_logic_vector(to_unsigned(131,8) ,
28850	 => std_logic_vector(to_unsigned(37,8) ,
28851	 => std_logic_vector(to_unsigned(4,8) ,
28852	 => std_logic_vector(to_unsigned(7,8) ,
28853	 => std_logic_vector(to_unsigned(59,8) ,
28854	 => std_logic_vector(to_unsigned(99,8) ,
28855	 => std_logic_vector(to_unsigned(115,8) ,
28856	 => std_logic_vector(to_unsigned(107,8) ,
28857	 => std_logic_vector(to_unsigned(80,8) ,
28858	 => std_logic_vector(to_unsigned(23,8) ,
28859	 => std_logic_vector(to_unsigned(9,8) ,
28860	 => std_logic_vector(to_unsigned(36,8) ,
28861	 => std_logic_vector(to_unsigned(42,8) ,
28862	 => std_logic_vector(to_unsigned(8,8) ,
28863	 => std_logic_vector(to_unsigned(1,8) ,
28864	 => std_logic_vector(to_unsigned(0,8) ,
28865	 => std_logic_vector(to_unsigned(0,8) ,
28866	 => std_logic_vector(to_unsigned(1,8) ,
28867	 => std_logic_vector(to_unsigned(1,8) ,
28868	 => std_logic_vector(to_unsigned(1,8) ,
28869	 => std_logic_vector(to_unsigned(3,8) ,
28870	 => std_logic_vector(to_unsigned(3,8) ,
28871	 => std_logic_vector(to_unsigned(5,8) ,
28872	 => std_logic_vector(to_unsigned(2,8) ,
28873	 => std_logic_vector(to_unsigned(2,8) ,
28874	 => std_logic_vector(to_unsigned(6,8) ,
28875	 => std_logic_vector(to_unsigned(8,8) ,
28876	 => std_logic_vector(to_unsigned(6,8) ,
28877	 => std_logic_vector(to_unsigned(6,8) ,
28878	 => std_logic_vector(to_unsigned(44,8) ,
28879	 => std_logic_vector(to_unsigned(93,8) ,
28880	 => std_logic_vector(to_unsigned(82,8) ,
28881	 => std_logic_vector(to_unsigned(72,8) ,
28882	 => std_logic_vector(to_unsigned(28,8) ,
28883	 => std_logic_vector(to_unsigned(26,8) ,
28884	 => std_logic_vector(to_unsigned(91,8) ,
28885	 => std_logic_vector(to_unsigned(72,8) ,
28886	 => std_logic_vector(to_unsigned(37,8) ,
28887	 => std_logic_vector(to_unsigned(14,8) ,
28888	 => std_logic_vector(to_unsigned(13,8) ,
28889	 => std_logic_vector(to_unsigned(20,8) ,
28890	 => std_logic_vector(to_unsigned(13,8) ,
28891	 => std_logic_vector(to_unsigned(4,8) ,
28892	 => std_logic_vector(to_unsigned(20,8) ,
28893	 => std_logic_vector(to_unsigned(139,8) ,
28894	 => std_logic_vector(to_unsigned(125,8) ,
28895	 => std_logic_vector(to_unsigned(116,8) ,
28896	 => std_logic_vector(to_unsigned(124,8) ,
28897	 => std_logic_vector(to_unsigned(164,8) ,
28898	 => std_logic_vector(to_unsigned(107,8) ,
28899	 => std_logic_vector(to_unsigned(6,8) ,
28900	 => std_logic_vector(to_unsigned(12,8) ,
28901	 => std_logic_vector(to_unsigned(42,8) ,
28902	 => std_logic_vector(to_unsigned(16,8) ,
28903	 => std_logic_vector(to_unsigned(41,8) ,
28904	 => std_logic_vector(to_unsigned(76,8) ,
28905	 => std_logic_vector(to_unsigned(48,8) ,
28906	 => std_logic_vector(to_unsigned(16,8) ,
28907	 => std_logic_vector(to_unsigned(16,8) ,
28908	 => std_logic_vector(to_unsigned(14,8) ,
28909	 => std_logic_vector(to_unsigned(13,8) ,
28910	 => std_logic_vector(to_unsigned(12,8) ,
28911	 => std_logic_vector(to_unsigned(6,8) ,
28912	 => std_logic_vector(to_unsigned(2,8) ,
28913	 => std_logic_vector(to_unsigned(93,8) ,
28914	 => std_logic_vector(to_unsigned(179,8) ,
28915	 => std_logic_vector(to_unsigned(25,8) ,
28916	 => std_logic_vector(to_unsigned(1,8) ,
28917	 => std_logic_vector(to_unsigned(3,8) ,
28918	 => std_logic_vector(to_unsigned(2,8) ,
28919	 => std_logic_vector(to_unsigned(2,8) ,
28920	 => std_logic_vector(to_unsigned(1,8) ,
28921	 => std_logic_vector(to_unsigned(1,8) ,
28922	 => std_logic_vector(to_unsigned(2,8) ,
28923	 => std_logic_vector(to_unsigned(2,8) ,
28924	 => std_logic_vector(to_unsigned(2,8) ,
28925	 => std_logic_vector(to_unsigned(1,8) ,
28926	 => std_logic_vector(to_unsigned(1,8) ,
28927	 => std_logic_vector(to_unsigned(0,8) ,
28928	 => std_logic_vector(to_unsigned(2,8) ,
28929	 => std_logic_vector(to_unsigned(39,8) ,
28930	 => std_logic_vector(to_unsigned(72,8) ,
28931	 => std_logic_vector(to_unsigned(53,8) ,
28932	 => std_logic_vector(to_unsigned(37,8) ,
28933	 => std_logic_vector(to_unsigned(17,8) ,
28934	 => std_logic_vector(to_unsigned(6,8) ,
28935	 => std_logic_vector(to_unsigned(40,8) ,
28936	 => std_logic_vector(to_unsigned(77,8) ,
28937	 => std_logic_vector(to_unsigned(53,8) ,
28938	 => std_logic_vector(to_unsigned(45,8) ,
28939	 => std_logic_vector(to_unsigned(37,8) ,
28940	 => std_logic_vector(to_unsigned(13,8) ,
28941	 => std_logic_vector(to_unsigned(2,8) ,
28942	 => std_logic_vector(to_unsigned(2,8) ,
28943	 => std_logic_vector(to_unsigned(2,8) ,
28944	 => std_logic_vector(to_unsigned(7,8) ,
28945	 => std_logic_vector(to_unsigned(15,8) ,
28946	 => std_logic_vector(to_unsigned(13,8) ,
28947	 => std_logic_vector(to_unsigned(20,8) ,
28948	 => std_logic_vector(to_unsigned(37,8) ,
28949	 => std_logic_vector(to_unsigned(25,8) ,
28950	 => std_logic_vector(to_unsigned(12,8) ,
28951	 => std_logic_vector(to_unsigned(17,8) ,
28952	 => std_logic_vector(to_unsigned(17,8) ,
28953	 => std_logic_vector(to_unsigned(10,8) ,
28954	 => std_logic_vector(to_unsigned(10,8) ,
28955	 => std_logic_vector(to_unsigned(6,8) ,
28956	 => std_logic_vector(to_unsigned(26,8) ,
28957	 => std_logic_vector(to_unsigned(71,8) ,
28958	 => std_logic_vector(to_unsigned(73,8) ,
28959	 => std_logic_vector(to_unsigned(82,8) ,
28960	 => std_logic_vector(to_unsigned(93,8) ,
28961	 => std_logic_vector(to_unsigned(70,8) ,
28962	 => std_logic_vector(to_unsigned(20,8) ,
28963	 => std_logic_vector(to_unsigned(11,8) ,
28964	 => std_logic_vector(to_unsigned(43,8) ,
28965	 => std_logic_vector(to_unsigned(70,8) ,
28966	 => std_logic_vector(to_unsigned(59,8) ,
28967	 => std_logic_vector(to_unsigned(36,8) ,
28968	 => std_logic_vector(to_unsigned(50,8) ,
28969	 => std_logic_vector(to_unsigned(157,8) ,
28970	 => std_logic_vector(to_unsigned(151,8) ,
28971	 => std_logic_vector(to_unsigned(18,8) ,
28972	 => std_logic_vector(to_unsigned(2,8) ,
28973	 => std_logic_vector(to_unsigned(12,8) ,
28974	 => std_logic_vector(to_unsigned(37,8) ,
28975	 => std_logic_vector(to_unsigned(39,8) ,
28976	 => std_logic_vector(to_unsigned(20,8) ,
28977	 => std_logic_vector(to_unsigned(16,8) ,
28978	 => std_logic_vector(to_unsigned(15,8) ,
28979	 => std_logic_vector(to_unsigned(15,8) ,
28980	 => std_logic_vector(to_unsigned(14,8) ,
28981	 => std_logic_vector(to_unsigned(8,8) ,
28982	 => std_logic_vector(to_unsigned(5,8) ,
28983	 => std_logic_vector(to_unsigned(6,8) ,
28984	 => std_logic_vector(to_unsigned(4,8) ,
28985	 => std_logic_vector(to_unsigned(2,8) ,
28986	 => std_logic_vector(to_unsigned(53,8) ,
28987	 => std_logic_vector(to_unsigned(170,8) ,
28988	 => std_logic_vector(to_unsigned(142,8) ,
28989	 => std_logic_vector(to_unsigned(149,8) ,
28990	 => std_logic_vector(to_unsigned(151,8) ,
28991	 => std_logic_vector(to_unsigned(156,8) ,
28992	 => std_logic_vector(to_unsigned(87,8) ,
28993	 => std_logic_vector(to_unsigned(93,8) ,
28994	 => std_logic_vector(to_unsigned(166,8) ,
28995	 => std_logic_vector(to_unsigned(154,8) ,
28996	 => std_logic_vector(to_unsigned(154,8) ,
28997	 => std_logic_vector(to_unsigned(152,8) ,
28998	 => std_logic_vector(to_unsigned(142,8) ,
28999	 => std_logic_vector(to_unsigned(134,8) ,
29000	 => std_logic_vector(to_unsigned(151,8) ,
29001	 => std_logic_vector(to_unsigned(154,8) ,
29002	 => std_logic_vector(to_unsigned(147,8) ,
29003	 => std_logic_vector(to_unsigned(149,8) ,
29004	 => std_logic_vector(to_unsigned(152,8) ,
29005	 => std_logic_vector(to_unsigned(152,8) ,
29006	 => std_logic_vector(to_unsigned(139,8) ,
29007	 => std_logic_vector(to_unsigned(111,8) ,
29008	 => std_logic_vector(to_unsigned(114,8) ,
29009	 => std_logic_vector(to_unsigned(154,8) ,
29010	 => std_logic_vector(to_unsigned(154,8) ,
29011	 => std_logic_vector(to_unsigned(156,8) ,
29012	 => std_logic_vector(to_unsigned(101,8) ,
29013	 => std_logic_vector(to_unsigned(115,8) ,
29014	 => std_logic_vector(to_unsigned(147,8) ,
29015	 => std_logic_vector(to_unsigned(127,8) ,
29016	 => std_logic_vector(to_unsigned(133,8) ,
29017	 => std_logic_vector(to_unsigned(53,8) ,
29018	 => std_logic_vector(to_unsigned(4,8) ,
29019	 => std_logic_vector(to_unsigned(8,8) ,
29020	 => std_logic_vector(to_unsigned(9,8) ,
29021	 => std_logic_vector(to_unsigned(5,8) ,
29022	 => std_logic_vector(to_unsigned(5,8) ,
29023	 => std_logic_vector(to_unsigned(104,8) ,
29024	 => std_logic_vector(to_unsigned(151,8) ,
29025	 => std_logic_vector(to_unsigned(144,8) ,
29026	 => std_logic_vector(to_unsigned(144,8) ,
29027	 => std_logic_vector(to_unsigned(139,8) ,
29028	 => std_logic_vector(to_unsigned(146,8) ,
29029	 => std_logic_vector(to_unsigned(149,8) ,
29030	 => std_logic_vector(to_unsigned(152,8) ,
29031	 => std_logic_vector(to_unsigned(154,8) ,
29032	 => std_logic_vector(to_unsigned(154,8) ,
29033	 => std_logic_vector(to_unsigned(175,8) ,
29034	 => std_logic_vector(to_unsigned(66,8) ,
29035	 => std_logic_vector(to_unsigned(3,8) ,
29036	 => std_logic_vector(to_unsigned(11,8) ,
29037	 => std_logic_vector(to_unsigned(30,8) ,
29038	 => std_logic_vector(to_unsigned(36,8) ,
29039	 => std_logic_vector(to_unsigned(23,8) ,
29040	 => std_logic_vector(to_unsigned(6,8) ,
29041	 => std_logic_vector(to_unsigned(5,8) ,
29042	 => std_logic_vector(to_unsigned(6,8) ,
29043	 => std_logic_vector(to_unsigned(11,8) ,
29044	 => std_logic_vector(to_unsigned(7,8) ,
29045	 => std_logic_vector(to_unsigned(9,8) ,
29046	 => std_logic_vector(to_unsigned(11,8) ,
29047	 => std_logic_vector(to_unsigned(8,8) ,
29048	 => std_logic_vector(to_unsigned(10,8) ,
29049	 => std_logic_vector(to_unsigned(9,8) ,
29050	 => std_logic_vector(to_unsigned(9,8) ,
29051	 => std_logic_vector(to_unsigned(7,8) ,
29052	 => std_logic_vector(to_unsigned(4,8) ,
29053	 => std_logic_vector(to_unsigned(7,8) ,
29054	 => std_logic_vector(to_unsigned(8,8) ,
29055	 => std_logic_vector(to_unsigned(10,8) ,
29056	 => std_logic_vector(to_unsigned(14,8) ,
29057	 => std_logic_vector(to_unsigned(17,8) ,
29058	 => std_logic_vector(to_unsigned(16,8) ,
29059	 => std_logic_vector(to_unsigned(9,8) ,
29060	 => std_logic_vector(to_unsigned(9,8) ,
29061	 => std_logic_vector(to_unsigned(58,8) ,
29062	 => std_logic_vector(to_unsigned(112,8) ,
29063	 => std_logic_vector(to_unsigned(97,8) ,
29064	 => std_logic_vector(to_unsigned(136,8) ,
29065	 => std_logic_vector(to_unsigned(90,8) ,
29066	 => std_logic_vector(to_unsigned(22,8) ,
29067	 => std_logic_vector(to_unsigned(24,8) ,
29068	 => std_logic_vector(to_unsigned(58,8) ,
29069	 => std_logic_vector(to_unsigned(40,8) ,
29070	 => std_logic_vector(to_unsigned(45,8) ,
29071	 => std_logic_vector(to_unsigned(80,8) ,
29072	 => std_logic_vector(to_unsigned(45,8) ,
29073	 => std_logic_vector(to_unsigned(62,8) ,
29074	 => std_logic_vector(to_unsigned(9,8) ,
29075	 => std_logic_vector(to_unsigned(1,8) ,
29076	 => std_logic_vector(to_unsigned(4,8) ,
29077	 => std_logic_vector(to_unsigned(4,8) ,
29078	 => std_logic_vector(to_unsigned(5,8) ,
29079	 => std_logic_vector(to_unsigned(4,8) ,
29080	 => std_logic_vector(to_unsigned(3,8) ,
29081	 => std_logic_vector(to_unsigned(3,8) ,
29082	 => std_logic_vector(to_unsigned(1,8) ,
29083	 => std_logic_vector(to_unsigned(1,8) ,
29084	 => std_logic_vector(to_unsigned(3,8) ,
29085	 => std_logic_vector(to_unsigned(4,8) ,
29086	 => std_logic_vector(to_unsigned(4,8) ,
29087	 => std_logic_vector(to_unsigned(2,8) ,
29088	 => std_logic_vector(to_unsigned(12,8) ,
29089	 => std_logic_vector(to_unsigned(29,8) ,
29090	 => std_logic_vector(to_unsigned(9,8) ,
29091	 => std_logic_vector(to_unsigned(6,8) ,
29092	 => std_logic_vector(to_unsigned(4,8) ,
29093	 => std_logic_vector(to_unsigned(5,8) ,
29094	 => std_logic_vector(to_unsigned(39,8) ,
29095	 => std_logic_vector(to_unsigned(48,8) ,
29096	 => std_logic_vector(to_unsigned(87,8) ,
29097	 => std_logic_vector(to_unsigned(101,8) ,
29098	 => std_logic_vector(to_unsigned(141,8) ,
29099	 => std_logic_vector(to_unsigned(170,8) ,
29100	 => std_logic_vector(to_unsigned(161,8) ,
29101	 => std_logic_vector(to_unsigned(138,8) ,
29102	 => std_logic_vector(to_unsigned(134,8) ,
29103	 => std_logic_vector(to_unsigned(147,8) ,
29104	 => std_logic_vector(to_unsigned(151,8) ,
29105	 => std_logic_vector(to_unsigned(156,8) ,
29106	 => std_logic_vector(to_unsigned(154,8) ,
29107	 => std_logic_vector(to_unsigned(164,8) ,
29108	 => std_logic_vector(to_unsigned(166,8) ,
29109	 => std_logic_vector(to_unsigned(171,8) ,
29110	 => std_logic_vector(to_unsigned(171,8) ,
29111	 => std_logic_vector(to_unsigned(170,8) ,
29112	 => std_logic_vector(to_unsigned(170,8) ,
29113	 => std_logic_vector(to_unsigned(166,8) ,
29114	 => std_logic_vector(to_unsigned(159,8) ,
29115	 => std_logic_vector(to_unsigned(151,8) ,
29116	 => std_logic_vector(to_unsigned(161,8) ,
29117	 => std_logic_vector(to_unsigned(164,8) ,
29118	 => std_logic_vector(to_unsigned(147,8) ,
29119	 => std_logic_vector(to_unsigned(144,8) ,
29120	 => std_logic_vector(to_unsigned(147,8) ,
29121	 => std_logic_vector(to_unsigned(86,8) ,
29122	 => std_logic_vector(to_unsigned(97,8) ,
29123	 => std_logic_vector(to_unsigned(108,8) ,
29124	 => std_logic_vector(to_unsigned(115,8) ,
29125	 => std_logic_vector(to_unsigned(130,8) ,
29126	 => std_logic_vector(to_unsigned(142,8) ,
29127	 => std_logic_vector(to_unsigned(95,8) ,
29128	 => std_logic_vector(to_unsigned(25,8) ,
29129	 => std_logic_vector(to_unsigned(81,8) ,
29130	 => std_logic_vector(to_unsigned(183,8) ,
29131	 => std_logic_vector(to_unsigned(147,8) ,
29132	 => std_logic_vector(to_unsigned(146,8) ,
29133	 => std_logic_vector(to_unsigned(142,8) ,
29134	 => std_logic_vector(to_unsigned(139,8) ,
29135	 => std_logic_vector(to_unsigned(138,8) ,
29136	 => std_logic_vector(to_unsigned(128,8) ,
29137	 => std_logic_vector(to_unsigned(118,8) ,
29138	 => std_logic_vector(to_unsigned(116,8) ,
29139	 => std_logic_vector(to_unsigned(32,8) ,
29140	 => std_logic_vector(to_unsigned(9,8) ,
29141	 => std_logic_vector(to_unsigned(22,8) ,
29142	 => std_logic_vector(to_unsigned(31,8) ,
29143	 => std_logic_vector(to_unsigned(51,8) ,
29144	 => std_logic_vector(to_unsigned(60,8) ,
29145	 => std_logic_vector(to_unsigned(23,8) ,
29146	 => std_logic_vector(to_unsigned(8,8) ,
29147	 => std_logic_vector(to_unsigned(3,8) ,
29148	 => std_logic_vector(to_unsigned(3,8) ,
29149	 => std_logic_vector(to_unsigned(2,8) ,
29150	 => std_logic_vector(to_unsigned(0,8) ,
29151	 => std_logic_vector(to_unsigned(0,8) ,
29152	 => std_logic_vector(to_unsigned(0,8) ,
29153	 => std_logic_vector(to_unsigned(3,8) ,
29154	 => std_logic_vector(to_unsigned(7,8) ,
29155	 => std_logic_vector(to_unsigned(13,8) ,
29156	 => std_logic_vector(to_unsigned(33,8) ,
29157	 => std_logic_vector(to_unsigned(46,8) ,
29158	 => std_logic_vector(to_unsigned(72,8) ,
29159	 => std_logic_vector(to_unsigned(91,8) ,
29160	 => std_logic_vector(to_unsigned(105,8) ,
29161	 => std_logic_vector(to_unsigned(119,8) ,
29162	 => std_logic_vector(to_unsigned(119,8) ,
29163	 => std_logic_vector(to_unsigned(141,8) ,
29164	 => std_logic_vector(to_unsigned(147,8) ,
29165	 => std_logic_vector(to_unsigned(151,8) ,
29166	 => std_logic_vector(to_unsigned(170,8) ,
29167	 => std_logic_vector(to_unsigned(170,8) ,
29168	 => std_logic_vector(to_unsigned(147,8) ,
29169	 => std_logic_vector(to_unsigned(144,8) ,
29170	 => std_logic_vector(to_unsigned(139,8) ,
29171	 => std_logic_vector(to_unsigned(42,8) ,
29172	 => std_logic_vector(to_unsigned(5,8) ,
29173	 => std_logic_vector(to_unsigned(22,8) ,
29174	 => std_logic_vector(to_unsigned(62,8) ,
29175	 => std_logic_vector(to_unsigned(97,8) ,
29176	 => std_logic_vector(to_unsigned(115,8) ,
29177	 => std_logic_vector(to_unsigned(116,8) ,
29178	 => std_logic_vector(to_unsigned(115,8) ,
29179	 => std_logic_vector(to_unsigned(141,8) ,
29180	 => std_logic_vector(to_unsigned(163,8) ,
29181	 => std_logic_vector(to_unsigned(164,8) ,
29182	 => std_logic_vector(to_unsigned(130,8) ,
29183	 => std_logic_vector(to_unsigned(73,8) ,
29184	 => std_logic_vector(to_unsigned(17,8) ,
29185	 => std_logic_vector(to_unsigned(3,8) ,
29186	 => std_logic_vector(to_unsigned(3,8) ,
29187	 => std_logic_vector(to_unsigned(3,8) ,
29188	 => std_logic_vector(to_unsigned(7,8) ,
29189	 => std_logic_vector(to_unsigned(7,8) ,
29190	 => std_logic_vector(to_unsigned(2,8) ,
29191	 => std_logic_vector(to_unsigned(6,8) ,
29192	 => std_logic_vector(to_unsigned(13,8) ,
29193	 => std_logic_vector(to_unsigned(7,8) ,
29194	 => std_logic_vector(to_unsigned(3,8) ,
29195	 => std_logic_vector(to_unsigned(6,8) ,
29196	 => std_logic_vector(to_unsigned(4,8) ,
29197	 => std_logic_vector(to_unsigned(3,8) ,
29198	 => std_logic_vector(to_unsigned(68,8) ,
29199	 => std_logic_vector(to_unsigned(173,8) ,
29200	 => std_logic_vector(to_unsigned(100,8) ,
29201	 => std_logic_vector(to_unsigned(45,8) ,
29202	 => std_logic_vector(to_unsigned(39,8) ,
29203	 => std_logic_vector(to_unsigned(127,8) ,
29204	 => std_logic_vector(to_unsigned(97,8) ,
29205	 => std_logic_vector(to_unsigned(15,8) ,
29206	 => std_logic_vector(to_unsigned(13,8) ,
29207	 => std_logic_vector(to_unsigned(3,8) ,
29208	 => std_logic_vector(to_unsigned(10,8) ,
29209	 => std_logic_vector(to_unsigned(13,8) ,
29210	 => std_logic_vector(to_unsigned(8,8) ,
29211	 => std_logic_vector(to_unsigned(3,8) ,
29212	 => std_logic_vector(to_unsigned(30,8) ,
29213	 => std_logic_vector(to_unsigned(121,8) ,
29214	 => std_logic_vector(to_unsigned(107,8) ,
29215	 => std_logic_vector(to_unsigned(130,8) ,
29216	 => std_logic_vector(to_unsigned(138,8) ,
29217	 => std_logic_vector(to_unsigned(93,8) ,
29218	 => std_logic_vector(to_unsigned(19,8) ,
29219	 => std_logic_vector(to_unsigned(4,8) ,
29220	 => std_logic_vector(to_unsigned(9,8) ,
29221	 => std_logic_vector(to_unsigned(6,8) ,
29222	 => std_logic_vector(to_unsigned(36,8) ,
29223	 => std_logic_vector(to_unsigned(91,8) ,
29224	 => std_logic_vector(to_unsigned(77,8) ,
29225	 => std_logic_vector(to_unsigned(51,8) ,
29226	 => std_logic_vector(to_unsigned(27,8) ,
29227	 => std_logic_vector(to_unsigned(19,8) ,
29228	 => std_logic_vector(to_unsigned(16,8) ,
29229	 => std_logic_vector(to_unsigned(10,8) ,
29230	 => std_logic_vector(to_unsigned(11,8) ,
29231	 => std_logic_vector(to_unsigned(3,8) ,
29232	 => std_logic_vector(to_unsigned(13,8) ,
29233	 => std_logic_vector(to_unsigned(149,8) ,
29234	 => std_logic_vector(to_unsigned(103,8) ,
29235	 => std_logic_vector(to_unsigned(4,8) ,
29236	 => std_logic_vector(to_unsigned(1,8) ,
29237	 => std_logic_vector(to_unsigned(2,8) ,
29238	 => std_logic_vector(to_unsigned(1,8) ,
29239	 => std_logic_vector(to_unsigned(1,8) ,
29240	 => std_logic_vector(to_unsigned(1,8) ,
29241	 => std_logic_vector(to_unsigned(1,8) ,
29242	 => std_logic_vector(to_unsigned(1,8) ,
29243	 => std_logic_vector(to_unsigned(2,8) ,
29244	 => std_logic_vector(to_unsigned(1,8) ,
29245	 => std_logic_vector(to_unsigned(1,8) ,
29246	 => std_logic_vector(to_unsigned(1,8) ,
29247	 => std_logic_vector(to_unsigned(0,8) ,
29248	 => std_logic_vector(to_unsigned(1,8) ,
29249	 => std_logic_vector(to_unsigned(36,8) ,
29250	 => std_logic_vector(to_unsigned(70,8) ,
29251	 => std_logic_vector(to_unsigned(53,8) ,
29252	 => std_logic_vector(to_unsigned(30,8) ,
29253	 => std_logic_vector(to_unsigned(11,8) ,
29254	 => std_logic_vector(to_unsigned(12,8) ,
29255	 => std_logic_vector(to_unsigned(39,8) ,
29256	 => std_logic_vector(to_unsigned(37,8) ,
29257	 => std_logic_vector(to_unsigned(37,8) ,
29258	 => std_logic_vector(to_unsigned(48,8) ,
29259	 => std_logic_vector(to_unsigned(22,8) ,
29260	 => std_logic_vector(to_unsigned(8,8) ,
29261	 => std_logic_vector(to_unsigned(36,8) ,
29262	 => std_logic_vector(to_unsigned(5,8) ,
29263	 => std_logic_vector(to_unsigned(1,8) ,
29264	 => std_logic_vector(to_unsigned(7,8) ,
29265	 => std_logic_vector(to_unsigned(9,8) ,
29266	 => std_logic_vector(to_unsigned(6,8) ,
29267	 => std_logic_vector(to_unsigned(12,8) ,
29268	 => std_logic_vector(to_unsigned(24,8) ,
29269	 => std_logic_vector(to_unsigned(19,8) ,
29270	 => std_logic_vector(to_unsigned(24,8) ,
29271	 => std_logic_vector(to_unsigned(23,8) ,
29272	 => std_logic_vector(to_unsigned(16,8) ,
29273	 => std_logic_vector(to_unsigned(11,8) ,
29274	 => std_logic_vector(to_unsigned(8,8) ,
29275	 => std_logic_vector(to_unsigned(2,8) ,
29276	 => std_logic_vector(to_unsigned(19,8) ,
29277	 => std_logic_vector(to_unsigned(81,8) ,
29278	 => std_logic_vector(to_unsigned(91,8) ,
29279	 => std_logic_vector(to_unsigned(84,8) ,
29280	 => std_logic_vector(to_unsigned(69,8) ,
29281	 => std_logic_vector(to_unsigned(32,8) ,
29282	 => std_logic_vector(to_unsigned(10,8) ,
29283	 => std_logic_vector(to_unsigned(17,8) ,
29284	 => std_logic_vector(to_unsigned(59,8) ,
29285	 => std_logic_vector(to_unsigned(77,8) ,
29286	 => std_logic_vector(to_unsigned(44,8) ,
29287	 => std_logic_vector(to_unsigned(22,8) ,
29288	 => std_logic_vector(to_unsigned(71,8) ,
29289	 => std_logic_vector(to_unsigned(166,8) ,
29290	 => std_logic_vector(to_unsigned(159,8) ,
29291	 => std_logic_vector(to_unsigned(25,8) ,
29292	 => std_logic_vector(to_unsigned(1,8) ,
29293	 => std_logic_vector(to_unsigned(10,8) ,
29294	 => std_logic_vector(to_unsigned(17,8) ,
29295	 => std_logic_vector(to_unsigned(12,8) ,
29296	 => std_logic_vector(to_unsigned(6,8) ,
29297	 => std_logic_vector(to_unsigned(11,8) ,
29298	 => std_logic_vector(to_unsigned(15,8) ,
29299	 => std_logic_vector(to_unsigned(17,8) ,
29300	 => std_logic_vector(to_unsigned(13,8) ,
29301	 => std_logic_vector(to_unsigned(8,8) ,
29302	 => std_logic_vector(to_unsigned(8,8) ,
29303	 => std_logic_vector(to_unsigned(10,8) ,
29304	 => std_logic_vector(to_unsigned(3,8) ,
29305	 => std_logic_vector(to_unsigned(3,8) ,
29306	 => std_logic_vector(to_unsigned(78,8) ,
29307	 => std_logic_vector(to_unsigned(164,8) ,
29308	 => std_logic_vector(to_unsigned(151,8) ,
29309	 => std_logic_vector(to_unsigned(151,8) ,
29310	 => std_logic_vector(to_unsigned(151,8) ,
29311	 => std_logic_vector(to_unsigned(152,8) ,
29312	 => std_logic_vector(to_unsigned(92,8) ,
29313	 => std_logic_vector(to_unsigned(66,8) ,
29314	 => std_logic_vector(to_unsigned(161,8) ,
29315	 => std_logic_vector(to_unsigned(154,8) ,
29316	 => std_logic_vector(to_unsigned(156,8) ,
29317	 => std_logic_vector(to_unsigned(156,8) ,
29318	 => std_logic_vector(to_unsigned(151,8) ,
29319	 => std_logic_vector(to_unsigned(141,8) ,
29320	 => std_logic_vector(to_unsigned(146,8) ,
29321	 => std_logic_vector(to_unsigned(149,8) ,
29322	 => std_logic_vector(to_unsigned(142,8) ,
29323	 => std_logic_vector(to_unsigned(147,8) ,
29324	 => std_logic_vector(to_unsigned(151,8) ,
29325	 => std_logic_vector(to_unsigned(147,8) ,
29326	 => std_logic_vector(to_unsigned(139,8) ,
29327	 => std_logic_vector(to_unsigned(79,8) ,
29328	 => std_logic_vector(to_unsigned(99,8) ,
29329	 => std_logic_vector(to_unsigned(159,8) ,
29330	 => std_logic_vector(to_unsigned(154,8) ,
29331	 => std_logic_vector(to_unsigned(159,8) ,
29332	 => std_logic_vector(to_unsigned(149,8) ,
29333	 => std_logic_vector(to_unsigned(139,8) ,
29334	 => std_logic_vector(to_unsigned(134,8) ,
29335	 => std_logic_vector(to_unsigned(146,8) ,
29336	 => std_logic_vector(to_unsigned(152,8) ,
29337	 => std_logic_vector(to_unsigned(31,8) ,
29338	 => std_logic_vector(to_unsigned(3,8) ,
29339	 => std_logic_vector(to_unsigned(9,8) ,
29340	 => std_logic_vector(to_unsigned(12,8) ,
29341	 => std_logic_vector(to_unsigned(4,8) ,
29342	 => std_logic_vector(to_unsigned(6,8) ,
29343	 => std_logic_vector(to_unsigned(100,8) ,
29344	 => std_logic_vector(to_unsigned(142,8) ,
29345	 => std_logic_vector(to_unsigned(138,8) ,
29346	 => std_logic_vector(to_unsigned(144,8) ,
29347	 => std_logic_vector(to_unsigned(147,8) ,
29348	 => std_logic_vector(to_unsigned(147,8) ,
29349	 => std_logic_vector(to_unsigned(149,8) ,
29350	 => std_logic_vector(to_unsigned(152,8) ,
29351	 => std_logic_vector(to_unsigned(157,8) ,
29352	 => std_logic_vector(to_unsigned(152,8) ,
29353	 => std_logic_vector(to_unsigned(171,8) ,
29354	 => std_logic_vector(to_unsigned(60,8) ,
29355	 => std_logic_vector(to_unsigned(1,8) ,
29356	 => std_logic_vector(to_unsigned(4,8) ,
29357	 => std_logic_vector(to_unsigned(19,8) ,
29358	 => std_logic_vector(to_unsigned(24,8) ,
29359	 => std_logic_vector(to_unsigned(16,8) ,
29360	 => std_logic_vector(to_unsigned(4,8) ,
29361	 => std_logic_vector(to_unsigned(6,8) ,
29362	 => std_logic_vector(to_unsigned(11,8) ,
29363	 => std_logic_vector(to_unsigned(11,8) ,
29364	 => std_logic_vector(to_unsigned(15,8) ,
29365	 => std_logic_vector(to_unsigned(7,8) ,
29366	 => std_logic_vector(to_unsigned(10,8) ,
29367	 => std_logic_vector(to_unsigned(9,8) ,
29368	 => std_logic_vector(to_unsigned(8,8) ,
29369	 => std_logic_vector(to_unsigned(5,8) ,
29370	 => std_logic_vector(to_unsigned(2,8) ,
29371	 => std_logic_vector(to_unsigned(9,8) ,
29372	 => std_logic_vector(to_unsigned(11,8) ,
29373	 => std_logic_vector(to_unsigned(13,8) ,
29374	 => std_logic_vector(to_unsigned(17,8) ,
29375	 => std_logic_vector(to_unsigned(9,8) ,
29376	 => std_logic_vector(to_unsigned(8,8) ,
29377	 => std_logic_vector(to_unsigned(8,8) ,
29378	 => std_logic_vector(to_unsigned(13,8) ,
29379	 => std_logic_vector(to_unsigned(28,8) ,
29380	 => std_logic_vector(to_unsigned(30,8) ,
29381	 => std_logic_vector(to_unsigned(54,8) ,
29382	 => std_logic_vector(to_unsigned(77,8) ,
29383	 => std_logic_vector(to_unsigned(70,8) ,
29384	 => std_logic_vector(to_unsigned(87,8) ,
29385	 => std_logic_vector(to_unsigned(37,8) ,
29386	 => std_logic_vector(to_unsigned(10,8) ,
29387	 => std_logic_vector(to_unsigned(16,8) ,
29388	 => std_logic_vector(to_unsigned(29,8) ,
29389	 => std_logic_vector(to_unsigned(42,8) ,
29390	 => std_logic_vector(to_unsigned(22,8) ,
29391	 => std_logic_vector(to_unsigned(61,8) ,
29392	 => std_logic_vector(to_unsigned(69,8) ,
29393	 => std_logic_vector(to_unsigned(37,8) ,
29394	 => std_logic_vector(to_unsigned(14,8) ,
29395	 => std_logic_vector(to_unsigned(1,8) ,
29396	 => std_logic_vector(to_unsigned(5,8) ,
29397	 => std_logic_vector(to_unsigned(4,8) ,
29398	 => std_logic_vector(to_unsigned(4,8) ,
29399	 => std_logic_vector(to_unsigned(4,8) ,
29400	 => std_logic_vector(to_unsigned(3,8) ,
29401	 => std_logic_vector(to_unsigned(2,8) ,
29402	 => std_logic_vector(to_unsigned(2,8) ,
29403	 => std_logic_vector(to_unsigned(2,8) ,
29404	 => std_logic_vector(to_unsigned(4,8) ,
29405	 => std_logic_vector(to_unsigned(3,8) ,
29406	 => std_logic_vector(to_unsigned(3,8) ,
29407	 => std_logic_vector(to_unsigned(2,8) ,
29408	 => std_logic_vector(to_unsigned(10,8) ,
29409	 => std_logic_vector(to_unsigned(18,8) ,
29410	 => std_logic_vector(to_unsigned(5,8) ,
29411	 => std_logic_vector(to_unsigned(5,8) ,
29412	 => std_logic_vector(to_unsigned(2,8) ,
29413	 => std_logic_vector(to_unsigned(13,8) ,
29414	 => std_logic_vector(to_unsigned(72,8) ,
29415	 => std_logic_vector(to_unsigned(96,8) ,
29416	 => std_logic_vector(to_unsigned(111,8) ,
29417	 => std_logic_vector(to_unsigned(90,8) ,
29418	 => std_logic_vector(to_unsigned(128,8) ,
29419	 => std_logic_vector(to_unsigned(170,8) ,
29420	 => std_logic_vector(to_unsigned(161,8) ,
29421	 => std_logic_vector(to_unsigned(139,8) ,
29422	 => std_logic_vector(to_unsigned(136,8) ,
29423	 => std_logic_vector(to_unsigned(147,8) ,
29424	 => std_logic_vector(to_unsigned(147,8) ,
29425	 => std_logic_vector(to_unsigned(147,8) ,
29426	 => std_logic_vector(to_unsigned(156,8) ,
29427	 => std_logic_vector(to_unsigned(164,8) ,
29428	 => std_logic_vector(to_unsigned(168,8) ,
29429	 => std_logic_vector(to_unsigned(168,8) ,
29430	 => std_logic_vector(to_unsigned(168,8) ,
29431	 => std_logic_vector(to_unsigned(166,8) ,
29432	 => std_logic_vector(to_unsigned(173,8) ,
29433	 => std_logic_vector(to_unsigned(171,8) ,
29434	 => std_logic_vector(to_unsigned(159,8) ,
29435	 => std_logic_vector(to_unsigned(154,8) ,
29436	 => std_logic_vector(to_unsigned(166,8) ,
29437	 => std_logic_vector(to_unsigned(166,8) ,
29438	 => std_logic_vector(to_unsigned(146,8) ,
29439	 => std_logic_vector(to_unsigned(138,8) ,
29440	 => std_logic_vector(to_unsigned(139,8) ,
29441	 => std_logic_vector(to_unsigned(4,8) ,
29442	 => std_logic_vector(to_unsigned(4,8) ,
29443	 => std_logic_vector(to_unsigned(6,8) ,
29444	 => std_logic_vector(to_unsigned(8,8) ,
29445	 => std_logic_vector(to_unsigned(9,8) ,
29446	 => std_logic_vector(to_unsigned(17,8) ,
29447	 => std_logic_vector(to_unsigned(14,8) ,
29448	 => std_logic_vector(to_unsigned(3,8) ,
29449	 => std_logic_vector(to_unsigned(55,8) ,
29450	 => std_logic_vector(to_unsigned(192,8) ,
29451	 => std_logic_vector(to_unsigned(166,8) ,
29452	 => std_logic_vector(to_unsigned(171,8) ,
29453	 => std_logic_vector(to_unsigned(173,8) ,
29454	 => std_logic_vector(to_unsigned(173,8) ,
29455	 => std_logic_vector(to_unsigned(177,8) ,
29456	 => std_logic_vector(to_unsigned(171,8) ,
29457	 => std_logic_vector(to_unsigned(168,8) ,
29458	 => std_logic_vector(to_unsigned(184,8) ,
29459	 => std_logic_vector(to_unsigned(64,8) ,
29460	 => std_logic_vector(to_unsigned(12,8) ,
29461	 => std_logic_vector(to_unsigned(21,8) ,
29462	 => std_logic_vector(to_unsigned(17,8) ,
29463	 => std_logic_vector(to_unsigned(37,8) ,
29464	 => std_logic_vector(to_unsigned(70,8) ,
29465	 => std_logic_vector(to_unsigned(17,8) ,
29466	 => std_logic_vector(to_unsigned(1,8) ,
29467	 => std_logic_vector(to_unsigned(1,8) ,
29468	 => std_logic_vector(to_unsigned(2,8) ,
29469	 => std_logic_vector(to_unsigned(1,8) ,
29470	 => std_logic_vector(to_unsigned(0,8) ,
29471	 => std_logic_vector(to_unsigned(0,8) ,
29472	 => std_logic_vector(to_unsigned(2,8) ,
29473	 => std_logic_vector(to_unsigned(3,8) ,
29474	 => std_logic_vector(to_unsigned(4,8) ,
29475	 => std_logic_vector(to_unsigned(3,8) ,
29476	 => std_logic_vector(to_unsigned(7,8) ,
29477	 => std_logic_vector(to_unsigned(11,8) ,
29478	 => std_logic_vector(to_unsigned(24,8) ,
29479	 => std_logic_vector(to_unsigned(32,8) ,
29480	 => std_logic_vector(to_unsigned(35,8) ,
29481	 => std_logic_vector(to_unsigned(55,8) ,
29482	 => std_logic_vector(to_unsigned(79,8) ,
29483	 => std_logic_vector(to_unsigned(118,8) ,
29484	 => std_logic_vector(to_unsigned(149,8) ,
29485	 => std_logic_vector(to_unsigned(164,8) ,
29486	 => std_logic_vector(to_unsigned(156,8) ,
29487	 => std_logic_vector(to_unsigned(147,8) ,
29488	 => std_logic_vector(to_unsigned(142,8) ,
29489	 => std_logic_vector(to_unsigned(141,8) ,
29490	 => std_logic_vector(to_unsigned(82,8) ,
29491	 => std_logic_vector(to_unsigned(11,8) ,
29492	 => std_logic_vector(to_unsigned(1,8) ,
29493	 => std_logic_vector(to_unsigned(6,8) ,
29494	 => std_logic_vector(to_unsigned(28,8) ,
29495	 => std_logic_vector(to_unsigned(59,8) ,
29496	 => std_logic_vector(to_unsigned(93,8) ,
29497	 => std_logic_vector(to_unsigned(97,8) ,
29498	 => std_logic_vector(to_unsigned(128,8) ,
29499	 => std_logic_vector(to_unsigned(177,8) ,
29500	 => std_logic_vector(to_unsigned(141,8) ,
29501	 => std_logic_vector(to_unsigned(124,8) ,
29502	 => std_logic_vector(to_unsigned(134,8) ,
29503	 => std_logic_vector(to_unsigned(168,8) ,
29504	 => std_logic_vector(to_unsigned(147,8) ,
29505	 => std_logic_vector(to_unsigned(91,8) ,
29506	 => std_logic_vector(to_unsigned(25,8) ,
29507	 => std_logic_vector(to_unsigned(21,8) ,
29508	 => std_logic_vector(to_unsigned(17,8) ,
29509	 => std_logic_vector(to_unsigned(1,8) ,
29510	 => std_logic_vector(to_unsigned(0,8) ,
29511	 => std_logic_vector(to_unsigned(5,8) ,
29512	 => std_logic_vector(to_unsigned(14,8) ,
29513	 => std_logic_vector(to_unsigned(7,8) ,
29514	 => std_logic_vector(to_unsigned(4,8) ,
29515	 => std_logic_vector(to_unsigned(8,8) ,
29516	 => std_logic_vector(to_unsigned(8,8) ,
29517	 => std_logic_vector(to_unsigned(3,8) ,
29518	 => std_logic_vector(to_unsigned(73,8) ,
29519	 => std_logic_vector(to_unsigned(183,8) ,
29520	 => std_logic_vector(to_unsigned(152,8) ,
29521	 => std_logic_vector(to_unsigned(122,8) ,
29522	 => std_logic_vector(to_unsigned(114,8) ,
29523	 => std_logic_vector(to_unsigned(108,8) ,
29524	 => std_logic_vector(to_unsigned(32,8) ,
29525	 => std_logic_vector(to_unsigned(6,8) ,
29526	 => std_logic_vector(to_unsigned(5,8) ,
29527	 => std_logic_vector(to_unsigned(2,8) ,
29528	 => std_logic_vector(to_unsigned(2,8) ,
29529	 => std_logic_vector(to_unsigned(6,8) ,
29530	 => std_logic_vector(to_unsigned(4,8) ,
29531	 => std_logic_vector(to_unsigned(1,8) ,
29532	 => std_logic_vector(to_unsigned(8,8) ,
29533	 => std_logic_vector(to_unsigned(15,8) ,
29534	 => std_logic_vector(to_unsigned(31,8) ,
29535	 => std_logic_vector(to_unsigned(53,8) ,
29536	 => std_logic_vector(to_unsigned(53,8) ,
29537	 => std_logic_vector(to_unsigned(28,8) ,
29538	 => std_logic_vector(to_unsigned(21,8) ,
29539	 => std_logic_vector(to_unsigned(32,8) ,
29540	 => std_logic_vector(to_unsigned(29,8) ,
29541	 => std_logic_vector(to_unsigned(57,8) ,
29542	 => std_logic_vector(to_unsigned(81,8) ,
29543	 => std_logic_vector(to_unsigned(77,8) ,
29544	 => std_logic_vector(to_unsigned(57,8) ,
29545	 => std_logic_vector(to_unsigned(25,8) ,
29546	 => std_logic_vector(to_unsigned(12,8) ,
29547	 => std_logic_vector(to_unsigned(21,8) ,
29548	 => std_logic_vector(to_unsigned(23,8) ,
29549	 => std_logic_vector(to_unsigned(15,8) ,
29550	 => std_logic_vector(to_unsigned(7,8) ,
29551	 => std_logic_vector(to_unsigned(3,8) ,
29552	 => std_logic_vector(to_unsigned(64,8) ,
29553	 => std_logic_vector(to_unsigned(170,8) ,
29554	 => std_logic_vector(to_unsigned(81,8) ,
29555	 => std_logic_vector(to_unsigned(2,8) ,
29556	 => std_logic_vector(to_unsigned(0,8) ,
29557	 => std_logic_vector(to_unsigned(1,8) ,
29558	 => std_logic_vector(to_unsigned(2,8) ,
29559	 => std_logic_vector(to_unsigned(1,8) ,
29560	 => std_logic_vector(to_unsigned(1,8) ,
29561	 => std_logic_vector(to_unsigned(1,8) ,
29562	 => std_logic_vector(to_unsigned(1,8) ,
29563	 => std_logic_vector(to_unsigned(1,8) ,
29564	 => std_logic_vector(to_unsigned(1,8) ,
29565	 => std_logic_vector(to_unsigned(1,8) ,
29566	 => std_logic_vector(to_unsigned(0,8) ,
29567	 => std_logic_vector(to_unsigned(0,8) ,
29568	 => std_logic_vector(to_unsigned(1,8) ,
29569	 => std_logic_vector(to_unsigned(30,8) ,
29570	 => std_logic_vector(to_unsigned(63,8) ,
29571	 => std_logic_vector(to_unsigned(47,8) ,
29572	 => std_logic_vector(to_unsigned(17,8) ,
29573	 => std_logic_vector(to_unsigned(7,8) ,
29574	 => std_logic_vector(to_unsigned(50,8) ,
29575	 => std_logic_vector(to_unsigned(93,8) ,
29576	 => std_logic_vector(to_unsigned(51,8) ,
29577	 => std_logic_vector(to_unsigned(33,8) ,
29578	 => std_logic_vector(to_unsigned(32,8) ,
29579	 => std_logic_vector(to_unsigned(18,8) ,
29580	 => std_logic_vector(to_unsigned(6,8) ,
29581	 => std_logic_vector(to_unsigned(74,8) ,
29582	 => std_logic_vector(to_unsigned(29,8) ,
29583	 => std_logic_vector(to_unsigned(2,8) ,
29584	 => std_logic_vector(to_unsigned(11,8) ,
29585	 => std_logic_vector(to_unsigned(8,8) ,
29586	 => std_logic_vector(to_unsigned(6,8) ,
29587	 => std_logic_vector(to_unsigned(12,8) ,
29588	 => std_logic_vector(to_unsigned(16,8) ,
29589	 => std_logic_vector(to_unsigned(25,8) ,
29590	 => std_logic_vector(to_unsigned(35,8) ,
29591	 => std_logic_vector(to_unsigned(27,8) ,
29592	 => std_logic_vector(to_unsigned(19,8) ,
29593	 => std_logic_vector(to_unsigned(11,8) ,
29594	 => std_logic_vector(to_unsigned(7,8) ,
29595	 => std_logic_vector(to_unsigned(4,8) ,
29596	 => std_logic_vector(to_unsigned(34,8) ,
29597	 => std_logic_vector(to_unsigned(67,8) ,
29598	 => std_logic_vector(to_unsigned(86,8) ,
29599	 => std_logic_vector(to_unsigned(115,8) ,
29600	 => std_logic_vector(to_unsigned(100,8) ,
29601	 => std_logic_vector(to_unsigned(46,8) ,
29602	 => std_logic_vector(to_unsigned(6,8) ,
29603	 => std_logic_vector(to_unsigned(23,8) ,
29604	 => std_logic_vector(to_unsigned(66,8) ,
29605	 => std_logic_vector(to_unsigned(79,8) ,
29606	 => std_logic_vector(to_unsigned(49,8) ,
29607	 => std_logic_vector(to_unsigned(27,8) ,
29608	 => std_logic_vector(to_unsigned(103,8) ,
29609	 => std_logic_vector(to_unsigned(164,8) ,
29610	 => std_logic_vector(to_unsigned(164,8) ,
29611	 => std_logic_vector(to_unsigned(34,8) ,
29612	 => std_logic_vector(to_unsigned(1,8) ,
29613	 => std_logic_vector(to_unsigned(4,8) ,
29614	 => std_logic_vector(to_unsigned(11,8) ,
29615	 => std_logic_vector(to_unsigned(13,8) ,
29616	 => std_logic_vector(to_unsigned(9,8) ,
29617	 => std_logic_vector(to_unsigned(8,8) ,
29618	 => std_logic_vector(to_unsigned(10,8) ,
29619	 => std_logic_vector(to_unsigned(12,8) ,
29620	 => std_logic_vector(to_unsigned(13,8) ,
29621	 => std_logic_vector(to_unsigned(9,8) ,
29622	 => std_logic_vector(to_unsigned(10,8) ,
29623	 => std_logic_vector(to_unsigned(12,8) ,
29624	 => std_logic_vector(to_unsigned(3,8) ,
29625	 => std_logic_vector(to_unsigned(4,8) ,
29626	 => std_logic_vector(to_unsigned(90,8) ,
29627	 => std_logic_vector(to_unsigned(164,8) ,
29628	 => std_logic_vector(to_unsigned(147,8) ,
29629	 => std_logic_vector(to_unsigned(149,8) ,
29630	 => std_logic_vector(to_unsigned(146,8) ,
29631	 => std_logic_vector(to_unsigned(136,8) ,
29632	 => std_logic_vector(to_unsigned(51,8) ,
29633	 => std_logic_vector(to_unsigned(52,8) ,
29634	 => std_logic_vector(to_unsigned(142,8) ,
29635	 => std_logic_vector(to_unsigned(144,8) ,
29636	 => std_logic_vector(to_unsigned(147,8) ,
29637	 => std_logic_vector(to_unsigned(147,8) ,
29638	 => std_logic_vector(to_unsigned(146,8) ,
29639	 => std_logic_vector(to_unsigned(147,8) ,
29640	 => std_logic_vector(to_unsigned(142,8) ,
29641	 => std_logic_vector(to_unsigned(142,8) ,
29642	 => std_logic_vector(to_unsigned(141,8) ,
29643	 => std_logic_vector(to_unsigned(139,8) ,
29644	 => std_logic_vector(to_unsigned(134,8) ,
29645	 => std_logic_vector(to_unsigned(141,8) ,
29646	 => std_logic_vector(to_unsigned(112,8) ,
29647	 => std_logic_vector(to_unsigned(58,8) ,
29648	 => std_logic_vector(to_unsigned(91,8) ,
29649	 => std_logic_vector(to_unsigned(152,8) ,
29650	 => std_logic_vector(to_unsigned(152,8) ,
29651	 => std_logic_vector(to_unsigned(151,8) ,
29652	 => std_logic_vector(to_unsigned(159,8) ,
29653	 => std_logic_vector(to_unsigned(149,8) ,
29654	 => std_logic_vector(to_unsigned(134,8) ,
29655	 => std_logic_vector(to_unsigned(154,8) ,
29656	 => std_logic_vector(to_unsigned(170,8) ,
29657	 => std_logic_vector(to_unsigned(35,8) ,
29658	 => std_logic_vector(to_unsigned(2,8) ,
29659	 => std_logic_vector(to_unsigned(6,8) ,
29660	 => std_logic_vector(to_unsigned(9,8) ,
29661	 => std_logic_vector(to_unsigned(3,8) ,
29662	 => std_logic_vector(to_unsigned(38,8) ,
29663	 => std_logic_vector(to_unsigned(107,8) ,
29664	 => std_logic_vector(to_unsigned(111,8) ,
29665	 => std_logic_vector(to_unsigned(141,8) ,
29666	 => std_logic_vector(to_unsigned(134,8) ,
29667	 => std_logic_vector(to_unsigned(134,8) ,
29668	 => std_logic_vector(to_unsigned(147,8) ,
29669	 => std_logic_vector(to_unsigned(152,8) ,
29670	 => std_logic_vector(to_unsigned(156,8) ,
29671	 => std_logic_vector(to_unsigned(161,8) ,
29672	 => std_logic_vector(to_unsigned(146,8) ,
29673	 => std_logic_vector(to_unsigned(170,8) ,
29674	 => std_logic_vector(to_unsigned(77,8) ,
29675	 => std_logic_vector(to_unsigned(1,8) ,
29676	 => std_logic_vector(to_unsigned(8,8) ,
29677	 => std_logic_vector(to_unsigned(25,8) ,
29678	 => std_logic_vector(to_unsigned(20,8) ,
29679	 => std_logic_vector(to_unsigned(12,8) ,
29680	 => std_logic_vector(to_unsigned(2,8) ,
29681	 => std_logic_vector(to_unsigned(4,8) ,
29682	 => std_logic_vector(to_unsigned(17,8) ,
29683	 => std_logic_vector(to_unsigned(10,8) ,
29684	 => std_logic_vector(to_unsigned(11,8) ,
29685	 => std_logic_vector(to_unsigned(11,8) ,
29686	 => std_logic_vector(to_unsigned(11,8) ,
29687	 => std_logic_vector(to_unsigned(9,8) ,
29688	 => std_logic_vector(to_unsigned(7,8) ,
29689	 => std_logic_vector(to_unsigned(3,8) ,
29690	 => std_logic_vector(to_unsigned(1,8) ,
29691	 => std_logic_vector(to_unsigned(4,8) ,
29692	 => std_logic_vector(to_unsigned(18,8) ,
29693	 => std_logic_vector(to_unsigned(32,8) ,
29694	 => std_logic_vector(to_unsigned(14,8) ,
29695	 => std_logic_vector(to_unsigned(6,8) ,
29696	 => std_logic_vector(to_unsigned(4,8) ,
29697	 => std_logic_vector(to_unsigned(9,8) ,
29698	 => std_logic_vector(to_unsigned(18,8) ,
29699	 => std_logic_vector(to_unsigned(18,8) ,
29700	 => std_logic_vector(to_unsigned(5,8) ,
29701	 => std_logic_vector(to_unsigned(10,8) ,
29702	 => std_logic_vector(to_unsigned(81,8) ,
29703	 => std_logic_vector(to_unsigned(97,8) ,
29704	 => std_logic_vector(to_unsigned(67,8) ,
29705	 => std_logic_vector(to_unsigned(35,8) ,
29706	 => std_logic_vector(to_unsigned(60,8) ,
29707	 => std_logic_vector(to_unsigned(82,8) ,
29708	 => std_logic_vector(to_unsigned(33,8) ,
29709	 => std_logic_vector(to_unsigned(53,8) ,
29710	 => std_logic_vector(to_unsigned(27,8) ,
29711	 => std_logic_vector(to_unsigned(55,8) ,
29712	 => std_logic_vector(to_unsigned(115,8) ,
29713	 => std_logic_vector(to_unsigned(51,8) ,
29714	 => std_logic_vector(to_unsigned(22,8) ,
29715	 => std_logic_vector(to_unsigned(3,8) ,
29716	 => std_logic_vector(to_unsigned(4,8) ,
29717	 => std_logic_vector(to_unsigned(4,8) ,
29718	 => std_logic_vector(to_unsigned(5,8) ,
29719	 => std_logic_vector(to_unsigned(3,8) ,
29720	 => std_logic_vector(to_unsigned(2,8) ,
29721	 => std_logic_vector(to_unsigned(5,8) ,
29722	 => std_logic_vector(to_unsigned(3,8) ,
29723	 => std_logic_vector(to_unsigned(3,8) ,
29724	 => std_logic_vector(to_unsigned(3,8) ,
29725	 => std_logic_vector(to_unsigned(3,8) ,
29726	 => std_logic_vector(to_unsigned(4,8) ,
29727	 => std_logic_vector(to_unsigned(3,8) ,
29728	 => std_logic_vector(to_unsigned(6,8) ,
29729	 => std_logic_vector(to_unsigned(10,8) ,
29730	 => std_logic_vector(to_unsigned(4,8) ,
29731	 => std_logic_vector(to_unsigned(2,8) ,
29732	 => std_logic_vector(to_unsigned(3,8) ,
29733	 => std_logic_vector(to_unsigned(41,8) ,
29734	 => std_logic_vector(to_unsigned(95,8) ,
29735	 => std_logic_vector(to_unsigned(99,8) ,
29736	 => std_logic_vector(to_unsigned(116,8) ,
29737	 => std_logic_vector(to_unsigned(105,8) ,
29738	 => std_logic_vector(to_unsigned(124,8) ,
29739	 => std_logic_vector(to_unsigned(149,8) ,
29740	 => std_logic_vector(to_unsigned(121,8) ,
29741	 => std_logic_vector(to_unsigned(146,8) ,
29742	 => std_logic_vector(to_unsigned(154,8) ,
29743	 => std_logic_vector(to_unsigned(147,8) ,
29744	 => std_logic_vector(to_unsigned(152,8) ,
29745	 => std_logic_vector(to_unsigned(151,8) ,
29746	 => std_logic_vector(to_unsigned(154,8) ,
29747	 => std_logic_vector(to_unsigned(161,8) ,
29748	 => std_logic_vector(to_unsigned(164,8) ,
29749	 => std_logic_vector(to_unsigned(161,8) ,
29750	 => std_logic_vector(to_unsigned(159,8) ,
29751	 => std_logic_vector(to_unsigned(159,8) ,
29752	 => std_logic_vector(to_unsigned(164,8) ,
29753	 => std_logic_vector(to_unsigned(164,8) ,
29754	 => std_logic_vector(to_unsigned(157,8) ,
29755	 => std_logic_vector(to_unsigned(156,8) ,
29756	 => std_logic_vector(to_unsigned(164,8) ,
29757	 => std_logic_vector(to_unsigned(164,8) ,
29758	 => std_logic_vector(to_unsigned(157,8) ,
29759	 => std_logic_vector(to_unsigned(157,8) ,
29760	 => std_logic_vector(to_unsigned(159,8) ,
29761	 => std_logic_vector(to_unsigned(57,8) ,
29762	 => std_logic_vector(to_unsigned(45,8) ,
29763	 => std_logic_vector(to_unsigned(37,8) ,
29764	 => std_logic_vector(to_unsigned(26,8) ,
29765	 => std_logic_vector(to_unsigned(23,8) ,
29766	 => std_logic_vector(to_unsigned(15,8) ,
29767	 => std_logic_vector(to_unsigned(8,8) ,
29768	 => std_logic_vector(to_unsigned(8,8) ,
29769	 => std_logic_vector(to_unsigned(12,8) ,
29770	 => std_logic_vector(to_unsigned(26,8) ,
29771	 => std_logic_vector(to_unsigned(30,8) ,
29772	 => std_logic_vector(to_unsigned(38,8) ,
29773	 => std_logic_vector(to_unsigned(45,8) ,
29774	 => std_logic_vector(to_unsigned(51,8) ,
29775	 => std_logic_vector(to_unsigned(64,8) ,
29776	 => std_logic_vector(to_unsigned(82,8) ,
29777	 => std_logic_vector(to_unsigned(95,8) ,
29778	 => std_logic_vector(to_unsigned(112,8) ,
29779	 => std_logic_vector(to_unsigned(96,8) ,
29780	 => std_logic_vector(to_unsigned(40,8) ,
29781	 => std_logic_vector(to_unsigned(36,8) ,
29782	 => std_logic_vector(to_unsigned(39,8) ,
29783	 => std_logic_vector(to_unsigned(41,8) ,
29784	 => std_logic_vector(to_unsigned(36,8) ,
29785	 => std_logic_vector(to_unsigned(4,8) ,
29786	 => std_logic_vector(to_unsigned(0,8) ,
29787	 => std_logic_vector(to_unsigned(1,8) ,
29788	 => std_logic_vector(to_unsigned(2,8) ,
29789	 => std_logic_vector(to_unsigned(2,8) ,
29790	 => std_logic_vector(to_unsigned(2,8) ,
29791	 => std_logic_vector(to_unsigned(3,8) ,
29792	 => std_logic_vector(to_unsigned(7,8) ,
29793	 => std_logic_vector(to_unsigned(6,8) ,
29794	 => std_logic_vector(to_unsigned(5,8) ,
29795	 => std_logic_vector(to_unsigned(4,8) ,
29796	 => std_logic_vector(to_unsigned(3,8) ,
29797	 => std_logic_vector(to_unsigned(2,8) ,
29798	 => std_logic_vector(to_unsigned(1,8) ,
29799	 => std_logic_vector(to_unsigned(1,8) ,
29800	 => std_logic_vector(to_unsigned(1,8) ,
29801	 => std_logic_vector(to_unsigned(1,8) ,
29802	 => std_logic_vector(to_unsigned(2,8) ,
29803	 => std_logic_vector(to_unsigned(4,8) ,
29804	 => std_logic_vector(to_unsigned(29,8) ,
29805	 => std_logic_vector(to_unsigned(114,8) ,
29806	 => std_logic_vector(to_unsigned(177,8) ,
29807	 => std_logic_vector(to_unsigned(159,8) ,
29808	 => std_logic_vector(to_unsigned(151,8) ,
29809	 => std_logic_vector(to_unsigned(151,8) ,
29810	 => std_logic_vector(to_unsigned(35,8) ,
29811	 => std_logic_vector(to_unsigned(3,8) ,
29812	 => std_logic_vector(to_unsigned(1,8) ,
29813	 => std_logic_vector(to_unsigned(1,8) ,
29814	 => std_logic_vector(to_unsigned(12,8) ,
29815	 => std_logic_vector(to_unsigned(41,8) ,
29816	 => std_logic_vector(to_unsigned(72,8) ,
29817	 => std_logic_vector(to_unsigned(54,8) ,
29818	 => std_logic_vector(to_unsigned(95,8) ,
29819	 => std_logic_vector(to_unsigned(147,8) ,
29820	 => std_logic_vector(to_unsigned(119,8) ,
29821	 => std_logic_vector(to_unsigned(108,8) ,
29822	 => std_logic_vector(to_unsigned(116,8) ,
29823	 => std_logic_vector(to_unsigned(133,8) ,
29824	 => std_logic_vector(to_unsigned(161,8) ,
29825	 => std_logic_vector(to_unsigned(118,8) ,
29826	 => std_logic_vector(to_unsigned(53,8) ,
29827	 => std_logic_vector(to_unsigned(32,8) ,
29828	 => std_logic_vector(to_unsigned(18,8) ,
29829	 => std_logic_vector(to_unsigned(4,8) ,
29830	 => std_logic_vector(to_unsigned(4,8) ,
29831	 => std_logic_vector(to_unsigned(3,8) ,
29832	 => std_logic_vector(to_unsigned(5,8) ,
29833	 => std_logic_vector(to_unsigned(4,8) ,
29834	 => std_logic_vector(to_unsigned(9,8) ,
29835	 => std_logic_vector(to_unsigned(12,8) ,
29836	 => std_logic_vector(to_unsigned(11,8) ,
29837	 => std_logic_vector(to_unsigned(11,8) ,
29838	 => std_logic_vector(to_unsigned(79,8) ,
29839	 => std_logic_vector(to_unsigned(179,8) ,
29840	 => std_logic_vector(to_unsigned(159,8) ,
29841	 => std_logic_vector(to_unsigned(161,8) ,
29842	 => std_logic_vector(to_unsigned(163,8) ,
29843	 => std_logic_vector(to_unsigned(173,8) ,
29844	 => std_logic_vector(to_unsigned(166,8) ,
29845	 => std_logic_vector(to_unsigned(131,8) ,
29846	 => std_logic_vector(to_unsigned(81,8) ,
29847	 => std_logic_vector(to_unsigned(37,8) ,
29848	 => std_logic_vector(to_unsigned(16,8) ,
29849	 => std_logic_vector(to_unsigned(3,8) ,
29850	 => std_logic_vector(to_unsigned(0,8) ,
29851	 => std_logic_vector(to_unsigned(0,8) ,
29852	 => std_logic_vector(to_unsigned(0,8) ,
29853	 => std_logic_vector(to_unsigned(0,8) ,
29854	 => std_logic_vector(to_unsigned(2,8) ,
29855	 => std_logic_vector(to_unsigned(3,8) ,
29856	 => std_logic_vector(to_unsigned(3,8) ,
29857	 => std_logic_vector(to_unsigned(17,8) ,
29858	 => std_logic_vector(to_unsigned(37,8) ,
29859	 => std_logic_vector(to_unsigned(37,8) ,
29860	 => std_logic_vector(to_unsigned(51,8) ,
29861	 => std_logic_vector(to_unsigned(82,8) ,
29862	 => std_logic_vector(to_unsigned(95,8) ,
29863	 => std_logic_vector(to_unsigned(72,8) ,
29864	 => std_logic_vector(to_unsigned(47,8) ,
29865	 => std_logic_vector(to_unsigned(19,8) ,
29866	 => std_logic_vector(to_unsigned(4,8) ,
29867	 => std_logic_vector(to_unsigned(30,8) ,
29868	 => std_logic_vector(to_unsigned(39,8) ,
29869	 => std_logic_vector(to_unsigned(14,8) ,
29870	 => std_logic_vector(to_unsigned(2,8) ,
29871	 => std_logic_vector(to_unsigned(7,8) ,
29872	 => std_logic_vector(to_unsigned(136,8) ,
29873	 => std_logic_vector(to_unsigned(175,8) ,
29874	 => std_logic_vector(to_unsigned(41,8) ,
29875	 => std_logic_vector(to_unsigned(1,8) ,
29876	 => std_logic_vector(to_unsigned(1,8) ,
29877	 => std_logic_vector(to_unsigned(1,8) ,
29878	 => std_logic_vector(to_unsigned(1,8) ,
29879	 => std_logic_vector(to_unsigned(0,8) ,
29880	 => std_logic_vector(to_unsigned(1,8) ,
29881	 => std_logic_vector(to_unsigned(1,8) ,
29882	 => std_logic_vector(to_unsigned(0,8) ,
29883	 => std_logic_vector(to_unsigned(0,8) ,
29884	 => std_logic_vector(to_unsigned(0,8) ,
29885	 => std_logic_vector(to_unsigned(1,8) ,
29886	 => std_logic_vector(to_unsigned(0,8) ,
29887	 => std_logic_vector(to_unsigned(0,8) ,
29888	 => std_logic_vector(to_unsigned(1,8) ,
29889	 => std_logic_vector(to_unsigned(27,8) ,
29890	 => std_logic_vector(to_unsigned(62,8) ,
29891	 => std_logic_vector(to_unsigned(34,8) ,
29892	 => std_logic_vector(to_unsigned(10,8) ,
29893	 => std_logic_vector(to_unsigned(9,8) ,
29894	 => std_logic_vector(to_unsigned(33,8) ,
29895	 => std_logic_vector(to_unsigned(43,8) ,
29896	 => std_logic_vector(to_unsigned(36,8) ,
29897	 => std_logic_vector(to_unsigned(41,8) ,
29898	 => std_logic_vector(to_unsigned(27,8) ,
29899	 => std_logic_vector(to_unsigned(8,8) ,
29900	 => std_logic_vector(to_unsigned(4,8) ,
29901	 => std_logic_vector(to_unsigned(105,8) ,
29902	 => std_logic_vector(to_unsigned(77,8) ,
29903	 => std_logic_vector(to_unsigned(2,8) ,
29904	 => std_logic_vector(to_unsigned(8,8) ,
29905	 => std_logic_vector(to_unsigned(6,8) ,
29906	 => std_logic_vector(to_unsigned(9,8) ,
29907	 => std_logic_vector(to_unsigned(17,8) ,
29908	 => std_logic_vector(to_unsigned(8,8) ,
29909	 => std_logic_vector(to_unsigned(20,8) ,
29910	 => std_logic_vector(to_unsigned(30,8) ,
29911	 => std_logic_vector(to_unsigned(18,8) ,
29912	 => std_logic_vector(to_unsigned(20,8) ,
29913	 => std_logic_vector(to_unsigned(11,8) ,
29914	 => std_logic_vector(to_unsigned(4,8) ,
29915	 => std_logic_vector(to_unsigned(12,8) ,
29916	 => std_logic_vector(to_unsigned(49,8) ,
29917	 => std_logic_vector(to_unsigned(56,8) ,
29918	 => std_logic_vector(to_unsigned(48,8) ,
29919	 => std_logic_vector(to_unsigned(57,8) ,
29920	 => std_logic_vector(to_unsigned(64,8) ,
29921	 => std_logic_vector(to_unsigned(67,8) ,
29922	 => std_logic_vector(to_unsigned(29,8) ,
29923	 => std_logic_vector(to_unsigned(24,8) ,
29924	 => std_logic_vector(to_unsigned(69,8) ,
29925	 => std_logic_vector(to_unsigned(81,8) ,
29926	 => std_logic_vector(to_unsigned(51,8) ,
29927	 => std_logic_vector(to_unsigned(42,8) ,
29928	 => std_logic_vector(to_unsigned(127,8) ,
29929	 => std_logic_vector(to_unsigned(151,8) ,
29930	 => std_logic_vector(to_unsigned(147,8) ,
29931	 => std_logic_vector(to_unsigned(28,8) ,
29932	 => std_logic_vector(to_unsigned(2,8) ,
29933	 => std_logic_vector(to_unsigned(3,8) ,
29934	 => std_logic_vector(to_unsigned(5,8) ,
29935	 => std_logic_vector(to_unsigned(11,8) ,
29936	 => std_logic_vector(to_unsigned(10,8) ,
29937	 => std_logic_vector(to_unsigned(7,8) ,
29938	 => std_logic_vector(to_unsigned(10,8) ,
29939	 => std_logic_vector(to_unsigned(11,8) ,
29940	 => std_logic_vector(to_unsigned(12,8) ,
29941	 => std_logic_vector(to_unsigned(12,8) ,
29942	 => std_logic_vector(to_unsigned(12,8) ,
29943	 => std_logic_vector(to_unsigned(9,8) ,
29944	 => std_logic_vector(to_unsigned(2,8) ,
29945	 => std_logic_vector(to_unsigned(10,8) ,
29946	 => std_logic_vector(to_unsigned(111,8) ,
29947	 => std_logic_vector(to_unsigned(157,8) ,
29948	 => std_logic_vector(to_unsigned(142,8) ,
29949	 => std_logic_vector(to_unsigned(152,8) ,
29950	 => std_logic_vector(to_unsigned(141,8) ,
29951	 => std_logic_vector(to_unsigned(134,8) ,
29952	 => std_logic_vector(to_unsigned(48,8) ,
29953	 => std_logic_vector(to_unsigned(19,8) ,
29954	 => std_logic_vector(to_unsigned(78,8) ,
29955	 => std_logic_vector(to_unsigned(142,8) ,
29956	 => std_logic_vector(to_unsigned(147,8) ,
29957	 => std_logic_vector(to_unsigned(146,8) ,
29958	 => std_logic_vector(to_unsigned(147,8) ,
29959	 => std_logic_vector(to_unsigned(142,8) ,
29960	 => std_logic_vector(to_unsigned(151,8) ,
29961	 => std_logic_vector(to_unsigned(146,8) ,
29962	 => std_logic_vector(to_unsigned(131,8) ,
29963	 => std_logic_vector(to_unsigned(149,8) ,
29964	 => std_logic_vector(to_unsigned(115,8) ,
29965	 => std_logic_vector(to_unsigned(103,8) ,
29966	 => std_logic_vector(to_unsigned(100,8) ,
29967	 => std_logic_vector(to_unsigned(56,8) ,
29968	 => std_logic_vector(to_unsigned(45,8) ,
29969	 => std_logic_vector(to_unsigned(127,8) ,
29970	 => std_logic_vector(to_unsigned(157,8) ,
29971	 => std_logic_vector(to_unsigned(151,8) ,
29972	 => std_logic_vector(to_unsigned(154,8) ,
29973	 => std_logic_vector(to_unsigned(149,8) ,
29974	 => std_logic_vector(to_unsigned(151,8) ,
29975	 => std_logic_vector(to_unsigned(157,8) ,
29976	 => std_logic_vector(to_unsigned(164,8) ,
29977	 => std_logic_vector(to_unsigned(149,8) ,
29978	 => std_logic_vector(to_unsigned(73,8) ,
29979	 => std_logic_vector(to_unsigned(26,8) ,
29980	 => std_logic_vector(to_unsigned(3,8) ,
29981	 => std_logic_vector(to_unsigned(10,8) ,
29982	 => std_logic_vector(to_unsigned(115,8) ,
29983	 => std_logic_vector(to_unsigned(99,8) ,
29984	 => std_logic_vector(to_unsigned(65,8) ,
29985	 => std_logic_vector(to_unsigned(109,8) ,
29986	 => std_logic_vector(to_unsigned(128,8) ,
29987	 => std_logic_vector(to_unsigned(133,8) ,
29988	 => std_logic_vector(to_unsigned(146,8) ,
29989	 => std_logic_vector(to_unsigned(141,8) ,
29990	 => std_logic_vector(to_unsigned(146,8) ,
29991	 => std_logic_vector(to_unsigned(156,8) ,
29992	 => std_logic_vector(to_unsigned(144,8) ,
29993	 => std_logic_vector(to_unsigned(146,8) ,
29994	 => std_logic_vector(to_unsigned(87,8) ,
29995	 => std_logic_vector(to_unsigned(6,8) ,
29996	 => std_logic_vector(to_unsigned(28,8) ,
29997	 => std_logic_vector(to_unsigned(47,8) ,
29998	 => std_logic_vector(to_unsigned(29,8) ,
29999	 => std_logic_vector(to_unsigned(9,8) ,
30000	 => std_logic_vector(to_unsigned(1,8) ,
30001	 => std_logic_vector(to_unsigned(4,8) ,
30002	 => std_logic_vector(to_unsigned(15,8) ,
30003	 => std_logic_vector(to_unsigned(17,8) ,
30004	 => std_logic_vector(to_unsigned(11,8) ,
30005	 => std_logic_vector(to_unsigned(12,8) ,
30006	 => std_logic_vector(to_unsigned(10,8) ,
30007	 => std_logic_vector(to_unsigned(8,8) ,
30008	 => std_logic_vector(to_unsigned(3,8) ,
30009	 => std_logic_vector(to_unsigned(2,8) ,
30010	 => std_logic_vector(to_unsigned(2,8) ,
30011	 => std_logic_vector(to_unsigned(1,8) ,
30012	 => std_logic_vector(to_unsigned(1,8) ,
30013	 => std_logic_vector(to_unsigned(3,8) ,
30014	 => std_logic_vector(to_unsigned(2,8) ,
30015	 => std_logic_vector(to_unsigned(0,8) ,
30016	 => std_logic_vector(to_unsigned(17,8) ,
30017	 => std_logic_vector(to_unsigned(52,8) ,
30018	 => std_logic_vector(to_unsigned(13,8) ,
30019	 => std_logic_vector(to_unsigned(18,8) ,
30020	 => std_logic_vector(to_unsigned(23,8) ,
30021	 => std_logic_vector(to_unsigned(24,8) ,
30022	 => std_logic_vector(to_unsigned(105,8) ,
30023	 => std_logic_vector(to_unsigned(58,8) ,
30024	 => std_logic_vector(to_unsigned(28,8) ,
30025	 => std_logic_vector(to_unsigned(13,8) ,
30026	 => std_logic_vector(to_unsigned(24,8) ,
30027	 => std_logic_vector(to_unsigned(35,8) ,
30028	 => std_logic_vector(to_unsigned(30,8) ,
30029	 => std_logic_vector(to_unsigned(55,8) ,
30030	 => std_logic_vector(to_unsigned(38,8) ,
30031	 => std_logic_vector(to_unsigned(82,8) ,
30032	 => std_logic_vector(to_unsigned(142,8) ,
30033	 => std_logic_vector(to_unsigned(111,8) ,
30034	 => std_logic_vector(to_unsigned(39,8) ,
30035	 => std_logic_vector(to_unsigned(2,8) ,
30036	 => std_logic_vector(to_unsigned(2,8) ,
30037	 => std_logic_vector(to_unsigned(3,8) ,
30038	 => std_logic_vector(to_unsigned(4,8) ,
30039	 => std_logic_vector(to_unsigned(3,8) ,
30040	 => std_logic_vector(to_unsigned(4,8) ,
30041	 => std_logic_vector(to_unsigned(8,8) ,
30042	 => std_logic_vector(to_unsigned(7,8) ,
30043	 => std_logic_vector(to_unsigned(4,8) ,
30044	 => std_logic_vector(to_unsigned(3,8) ,
30045	 => std_logic_vector(to_unsigned(3,8) ,
30046	 => std_logic_vector(to_unsigned(2,8) ,
30047	 => std_logic_vector(to_unsigned(1,8) ,
30048	 => std_logic_vector(to_unsigned(1,8) ,
30049	 => std_logic_vector(to_unsigned(5,8) ,
30050	 => std_logic_vector(to_unsigned(2,8) ,
30051	 => std_logic_vector(to_unsigned(0,8) ,
30052	 => std_logic_vector(to_unsigned(6,8) ,
30053	 => std_logic_vector(to_unsigned(73,8) ,
30054	 => std_logic_vector(to_unsigned(96,8) ,
30055	 => std_logic_vector(to_unsigned(91,8) ,
30056	 => std_logic_vector(to_unsigned(130,8) ,
30057	 => std_logic_vector(to_unsigned(138,8) ,
30058	 => std_logic_vector(to_unsigned(146,8) ,
30059	 => std_logic_vector(to_unsigned(144,8) ,
30060	 => std_logic_vector(to_unsigned(134,8) ,
30061	 => std_logic_vector(to_unsigned(166,8) ,
30062	 => std_logic_vector(to_unsigned(166,8) ,
30063	 => std_logic_vector(to_unsigned(161,8) ,
30064	 => std_logic_vector(to_unsigned(156,8) ,
30065	 => std_logic_vector(to_unsigned(154,8) ,
30066	 => std_logic_vector(to_unsigned(157,8) ,
30067	 => std_logic_vector(to_unsigned(159,8) ,
30068	 => std_logic_vector(to_unsigned(163,8) ,
30069	 => std_logic_vector(to_unsigned(159,8) ,
30070	 => std_logic_vector(to_unsigned(157,8) ,
30071	 => std_logic_vector(to_unsigned(156,8) ,
30072	 => std_logic_vector(to_unsigned(156,8) ,
30073	 => std_logic_vector(to_unsigned(157,8) ,
30074	 => std_logic_vector(to_unsigned(156,8) ,
30075	 => std_logic_vector(to_unsigned(156,8) ,
30076	 => std_logic_vector(to_unsigned(156,8) ,
30077	 => std_logic_vector(to_unsigned(154,8) ,
30078	 => std_logic_vector(to_unsigned(156,8) ,
30079	 => std_logic_vector(to_unsigned(154,8) ,
30080	 => std_logic_vector(to_unsigned(151,8) ,
30081	 => std_logic_vector(to_unsigned(206,8) ,
30082	 => std_logic_vector(to_unsigned(208,8) ,
30083	 => std_logic_vector(to_unsigned(206,8) ,
30084	 => std_logic_vector(to_unsigned(210,8) ,
30085	 => std_logic_vector(to_unsigned(210,8) ,
30086	 => std_logic_vector(to_unsigned(69,8) ,
30087	 => std_logic_vector(to_unsigned(7,8) ,
30088	 => std_logic_vector(to_unsigned(8,8) ,
30089	 => std_logic_vector(to_unsigned(4,8) ,
30090	 => std_logic_vector(to_unsigned(1,8) ,
30091	 => std_logic_vector(to_unsigned(1,8) ,
30092	 => std_logic_vector(to_unsigned(0,8) ,
30093	 => std_logic_vector(to_unsigned(0,8) ,
30094	 => std_logic_vector(to_unsigned(0,8) ,
30095	 => std_logic_vector(to_unsigned(0,8) ,
30096	 => std_logic_vector(to_unsigned(1,8) ,
30097	 => std_logic_vector(to_unsigned(2,8) ,
30098	 => std_logic_vector(to_unsigned(3,8) ,
30099	 => std_logic_vector(to_unsigned(8,8) ,
30100	 => std_logic_vector(to_unsigned(8,8) ,
30101	 => std_logic_vector(to_unsigned(11,8) ,
30102	 => std_logic_vector(to_unsigned(15,8) ,
30103	 => std_logic_vector(to_unsigned(14,8) ,
30104	 => std_logic_vector(to_unsigned(8,8) ,
30105	 => std_logic_vector(to_unsigned(1,8) ,
30106	 => std_logic_vector(to_unsigned(2,8) ,
30107	 => std_logic_vector(to_unsigned(1,8) ,
30108	 => std_logic_vector(to_unsigned(2,8) ,
30109	 => std_logic_vector(to_unsigned(7,8) ,
30110	 => std_logic_vector(to_unsigned(13,8) ,
30111	 => std_logic_vector(to_unsigned(10,8) ,
30112	 => std_logic_vector(to_unsigned(8,8) ,
30113	 => std_logic_vector(to_unsigned(7,8) ,
30114	 => std_logic_vector(to_unsigned(7,8) ,
30115	 => std_logic_vector(to_unsigned(7,8) ,
30116	 => std_logic_vector(to_unsigned(5,8) ,
30117	 => std_logic_vector(to_unsigned(5,8) ,
30118	 => std_logic_vector(to_unsigned(3,8) ,
30119	 => std_logic_vector(to_unsigned(2,8) ,
30120	 => std_logic_vector(to_unsigned(1,8) ,
30121	 => std_logic_vector(to_unsigned(1,8) ,
30122	 => std_logic_vector(to_unsigned(2,8) ,
30123	 => std_logic_vector(to_unsigned(7,8) ,
30124	 => std_logic_vector(to_unsigned(11,8) ,
30125	 => std_logic_vector(to_unsigned(11,8) ,
30126	 => std_logic_vector(to_unsigned(61,8) ,
30127	 => std_logic_vector(to_unsigned(139,8) ,
30128	 => std_logic_vector(to_unsigned(128,8) ,
30129	 => std_logic_vector(to_unsigned(62,8) ,
30130	 => std_logic_vector(to_unsigned(10,8) ,
30131	 => std_logic_vector(to_unsigned(4,8) ,
30132	 => std_logic_vector(to_unsigned(1,8) ,
30133	 => std_logic_vector(to_unsigned(1,8) ,
30134	 => std_logic_vector(to_unsigned(3,8) ,
30135	 => std_logic_vector(to_unsigned(10,8) ,
30136	 => std_logic_vector(to_unsigned(31,8) ,
30137	 => std_logic_vector(to_unsigned(16,8) ,
30138	 => std_logic_vector(to_unsigned(30,8) ,
30139	 => std_logic_vector(to_unsigned(74,8) ,
30140	 => std_logic_vector(to_unsigned(69,8) ,
30141	 => std_logic_vector(to_unsigned(96,8) ,
30142	 => std_logic_vector(to_unsigned(131,8) ,
30143	 => std_logic_vector(to_unsigned(144,8) ,
30144	 => std_logic_vector(to_unsigned(112,8) ,
30145	 => std_logic_vector(to_unsigned(43,8) ,
30146	 => std_logic_vector(to_unsigned(81,8) ,
30147	 => std_logic_vector(to_unsigned(45,8) ,
30148	 => std_logic_vector(to_unsigned(6,8) ,
30149	 => std_logic_vector(to_unsigned(6,8) ,
30150	 => std_logic_vector(to_unsigned(12,8) ,
30151	 => std_logic_vector(to_unsigned(6,8) ,
30152	 => std_logic_vector(to_unsigned(4,8) ,
30153	 => std_logic_vector(to_unsigned(10,8) ,
30154	 => std_logic_vector(to_unsigned(19,8) ,
30155	 => std_logic_vector(to_unsigned(13,8) ,
30156	 => std_logic_vector(to_unsigned(16,8) ,
30157	 => std_logic_vector(to_unsigned(13,8) ,
30158	 => std_logic_vector(to_unsigned(24,8) ,
30159	 => std_logic_vector(to_unsigned(121,8) ,
30160	 => std_logic_vector(to_unsigned(170,8) ,
30161	 => std_logic_vector(to_unsigned(82,8) ,
30162	 => std_logic_vector(to_unsigned(68,8) ,
30163	 => std_logic_vector(to_unsigned(107,8) ,
30164	 => std_logic_vector(to_unsigned(136,8) ,
30165	 => std_logic_vector(to_unsigned(168,8) ,
30166	 => std_logic_vector(to_unsigned(192,8) ,
30167	 => std_logic_vector(to_unsigned(202,8) ,
30168	 => std_logic_vector(to_unsigned(171,8) ,
30169	 => std_logic_vector(to_unsigned(107,8) ,
30170	 => std_logic_vector(to_unsigned(51,8) ,
30171	 => std_logic_vector(to_unsigned(30,8) ,
30172	 => std_logic_vector(to_unsigned(9,8) ,
30173	 => std_logic_vector(to_unsigned(1,8) ,
30174	 => std_logic_vector(to_unsigned(1,8) ,
30175	 => std_logic_vector(to_unsigned(12,8) ,
30176	 => std_logic_vector(to_unsigned(19,8) ,
30177	 => std_logic_vector(to_unsigned(25,8) ,
30178	 => std_logic_vector(to_unsigned(31,8) ,
30179	 => std_logic_vector(to_unsigned(32,8) ,
30180	 => std_logic_vector(to_unsigned(43,8) ,
30181	 => std_logic_vector(to_unsigned(43,8) ,
30182	 => std_logic_vector(to_unsigned(68,8) ,
30183	 => std_logic_vector(to_unsigned(64,8) ,
30184	 => std_logic_vector(to_unsigned(19,8) ,
30185	 => std_logic_vector(to_unsigned(2,8) ,
30186	 => std_logic_vector(to_unsigned(3,8) ,
30187	 => std_logic_vector(to_unsigned(41,8) ,
30188	 => std_logic_vector(to_unsigned(60,8) ,
30189	 => std_logic_vector(to_unsigned(24,8) ,
30190	 => std_logic_vector(to_unsigned(5,8) ,
30191	 => std_logic_vector(to_unsigned(6,8) ,
30192	 => std_logic_vector(to_unsigned(66,8) ,
30193	 => std_logic_vector(to_unsigned(55,8) ,
30194	 => std_logic_vector(to_unsigned(2,8) ,
30195	 => std_logic_vector(to_unsigned(1,8) ,
30196	 => std_logic_vector(to_unsigned(1,8) ,
30197	 => std_logic_vector(to_unsigned(0,8) ,
30198	 => std_logic_vector(to_unsigned(0,8) ,
30199	 => std_logic_vector(to_unsigned(0,8) ,
30200	 => std_logic_vector(to_unsigned(0,8) ,
30201	 => std_logic_vector(to_unsigned(0,8) ,
30202	 => std_logic_vector(to_unsigned(0,8) ,
30203	 => std_logic_vector(to_unsigned(0,8) ,
30204	 => std_logic_vector(to_unsigned(0,8) ,
30205	 => std_logic_vector(to_unsigned(0,8) ,
30206	 => std_logic_vector(to_unsigned(0,8) ,
30207	 => std_logic_vector(to_unsigned(0,8) ,
30208	 => std_logic_vector(to_unsigned(0,8) ,
30209	 => std_logic_vector(to_unsigned(14,8) ,
30210	 => std_logic_vector(to_unsigned(70,8) ,
30211	 => std_logic_vector(to_unsigned(34,8) ,
30212	 => std_logic_vector(to_unsigned(13,8) ,
30213	 => std_logic_vector(to_unsigned(29,8) ,
30214	 => std_logic_vector(to_unsigned(32,8) ,
30215	 => std_logic_vector(to_unsigned(23,8) ,
30216	 => std_logic_vector(to_unsigned(16,8) ,
30217	 => std_logic_vector(to_unsigned(12,8) ,
30218	 => std_logic_vector(to_unsigned(24,8) ,
30219	 => std_logic_vector(to_unsigned(5,8) ,
30220	 => std_logic_vector(to_unsigned(14,8) ,
30221	 => std_logic_vector(to_unsigned(159,8) ,
30222	 => std_logic_vector(to_unsigned(125,8) ,
30223	 => std_logic_vector(to_unsigned(5,8) ,
30224	 => std_logic_vector(to_unsigned(4,8) ,
30225	 => std_logic_vector(to_unsigned(7,8) ,
30226	 => std_logic_vector(to_unsigned(6,8) ,
30227	 => std_logic_vector(to_unsigned(12,8) ,
30228	 => std_logic_vector(to_unsigned(12,8) ,
30229	 => std_logic_vector(to_unsigned(16,8) ,
30230	 => std_logic_vector(to_unsigned(11,8) ,
30231	 => std_logic_vector(to_unsigned(7,8) ,
30232	 => std_logic_vector(to_unsigned(13,8) ,
30233	 => std_logic_vector(to_unsigned(22,8) ,
30234	 => std_logic_vector(to_unsigned(27,8) ,
30235	 => std_logic_vector(to_unsigned(38,8) ,
30236	 => std_logic_vector(to_unsigned(28,8) ,
30237	 => std_logic_vector(to_unsigned(20,8) ,
30238	 => std_logic_vector(to_unsigned(22,8) ,
30239	 => std_logic_vector(to_unsigned(13,8) ,
30240	 => std_logic_vector(to_unsigned(5,8) ,
30241	 => std_logic_vector(to_unsigned(5,8) ,
30242	 => std_logic_vector(to_unsigned(23,8) ,
30243	 => std_logic_vector(to_unsigned(37,8) ,
30244	 => std_logic_vector(to_unsigned(71,8) ,
30245	 => std_logic_vector(to_unsigned(80,8) ,
30246	 => std_logic_vector(to_unsigned(53,8) ,
30247	 => std_logic_vector(to_unsigned(63,8) ,
30248	 => std_logic_vector(to_unsigned(149,8) ,
30249	 => std_logic_vector(to_unsigned(175,8) ,
30250	 => std_logic_vector(to_unsigned(130,8) ,
30251	 => std_logic_vector(to_unsigned(8,8) ,
30252	 => std_logic_vector(to_unsigned(1,8) ,
30253	 => std_logic_vector(to_unsigned(7,8) ,
30254	 => std_logic_vector(to_unsigned(8,8) ,
30255	 => std_logic_vector(to_unsigned(8,8) ,
30256	 => std_logic_vector(to_unsigned(8,8) ,
30257	 => std_logic_vector(to_unsigned(6,8) ,
30258	 => std_logic_vector(to_unsigned(7,8) ,
30259	 => std_logic_vector(to_unsigned(12,8) ,
30260	 => std_logic_vector(to_unsigned(15,8) ,
30261	 => std_logic_vector(to_unsigned(17,8) ,
30262	 => std_logic_vector(to_unsigned(8,8) ,
30263	 => std_logic_vector(to_unsigned(2,8) ,
30264	 => std_logic_vector(to_unsigned(5,8) ,
30265	 => std_logic_vector(to_unsigned(42,8) ,
30266	 => std_logic_vector(to_unsigned(134,8) ,
30267	 => std_logic_vector(to_unsigned(156,8) ,
30268	 => std_logic_vector(to_unsigned(151,8) ,
30269	 => std_logic_vector(to_unsigned(149,8) ,
30270	 => std_logic_vector(to_unsigned(139,8) ,
30271	 => std_logic_vector(to_unsigned(93,8) ,
30272	 => std_logic_vector(to_unsigned(61,8) ,
30273	 => std_logic_vector(to_unsigned(8,8) ,
30274	 => std_logic_vector(to_unsigned(23,8) ,
30275	 => std_logic_vector(to_unsigned(105,8) ,
30276	 => std_logic_vector(to_unsigned(133,8) ,
30277	 => std_logic_vector(to_unsigned(144,8) ,
30278	 => std_logic_vector(to_unsigned(151,8) ,
30279	 => std_logic_vector(to_unsigned(141,8) ,
30280	 => std_logic_vector(to_unsigned(156,8) ,
30281	 => std_logic_vector(to_unsigned(151,8) ,
30282	 => std_logic_vector(to_unsigned(78,8) ,
30283	 => std_logic_vector(to_unsigned(90,8) ,
30284	 => std_logic_vector(to_unsigned(93,8) ,
30285	 => std_logic_vector(to_unsigned(72,8) ,
30286	 => std_logic_vector(to_unsigned(33,8) ,
30287	 => std_logic_vector(to_unsigned(3,8) ,
30288	 => std_logic_vector(to_unsigned(11,8) ,
30289	 => std_logic_vector(to_unsigned(101,8) ,
30290	 => std_logic_vector(to_unsigned(151,8) ,
30291	 => std_logic_vector(to_unsigned(154,8) ,
30292	 => std_logic_vector(to_unsigned(151,8) ,
30293	 => std_logic_vector(to_unsigned(152,8) ,
30294	 => std_logic_vector(to_unsigned(159,8) ,
30295	 => std_logic_vector(to_unsigned(157,8) ,
30296	 => std_logic_vector(to_unsigned(161,8) ,
30297	 => std_logic_vector(to_unsigned(166,8) ,
30298	 => std_logic_vector(to_unsigned(183,8) ,
30299	 => std_logic_vector(to_unsigned(163,8) ,
30300	 => std_logic_vector(to_unsigned(73,8) ,
30301	 => std_logic_vector(to_unsigned(90,8) ,
30302	 => std_logic_vector(to_unsigned(138,8) ,
30303	 => std_logic_vector(to_unsigned(111,8) ,
30304	 => std_logic_vector(to_unsigned(76,8) ,
30305	 => std_logic_vector(to_unsigned(77,8) ,
30306	 => std_logic_vector(to_unsigned(121,8) ,
30307	 => std_logic_vector(to_unsigned(133,8) ,
30308	 => std_logic_vector(to_unsigned(139,8) ,
30309	 => std_logic_vector(to_unsigned(131,8) ,
30310	 => std_logic_vector(to_unsigned(128,8) ,
30311	 => std_logic_vector(to_unsigned(133,8) ,
30312	 => std_logic_vector(to_unsigned(122,8) ,
30313	 => std_logic_vector(to_unsigned(88,8) ,
30314	 => std_logic_vector(to_unsigned(31,8) ,
30315	 => std_logic_vector(to_unsigned(18,8) ,
30316	 => std_logic_vector(to_unsigned(50,8) ,
30317	 => std_logic_vector(to_unsigned(65,8) ,
30318	 => std_logic_vector(to_unsigned(43,8) ,
30319	 => std_logic_vector(to_unsigned(6,8) ,
30320	 => std_logic_vector(to_unsigned(1,8) ,
30321	 => std_logic_vector(to_unsigned(8,8) ,
30322	 => std_logic_vector(to_unsigned(16,8) ,
30323	 => std_logic_vector(to_unsigned(20,8) ,
30324	 => std_logic_vector(to_unsigned(15,8) ,
30325	 => std_logic_vector(to_unsigned(12,8) ,
30326	 => std_logic_vector(to_unsigned(9,8) ,
30327	 => std_logic_vector(to_unsigned(5,8) ,
30328	 => std_logic_vector(to_unsigned(2,8) ,
30329	 => std_logic_vector(to_unsigned(3,8) ,
30330	 => std_logic_vector(to_unsigned(2,8) ,
30331	 => std_logic_vector(to_unsigned(2,8) ,
30332	 => std_logic_vector(to_unsigned(1,8) ,
30333	 => std_logic_vector(to_unsigned(1,8) ,
30334	 => std_logic_vector(to_unsigned(3,8) ,
30335	 => std_logic_vector(to_unsigned(3,8) ,
30336	 => std_logic_vector(to_unsigned(14,8) ,
30337	 => std_logic_vector(to_unsigned(66,8) ,
30338	 => std_logic_vector(to_unsigned(77,8) ,
30339	 => std_logic_vector(to_unsigned(68,8) ,
30340	 => std_logic_vector(to_unsigned(29,8) ,
30341	 => std_logic_vector(to_unsigned(10,8) ,
30342	 => std_logic_vector(to_unsigned(41,8) ,
30343	 => std_logic_vector(to_unsigned(23,8) ,
30344	 => std_logic_vector(to_unsigned(12,8) ,
30345	 => std_logic_vector(to_unsigned(24,8) ,
30346	 => std_logic_vector(to_unsigned(32,8) ,
30347	 => std_logic_vector(to_unsigned(30,8) ,
30348	 => std_logic_vector(to_unsigned(51,8) ,
30349	 => std_logic_vector(to_unsigned(33,8) ,
30350	 => std_logic_vector(to_unsigned(41,8) ,
30351	 => std_logic_vector(to_unsigned(96,8) ,
30352	 => std_logic_vector(to_unsigned(138,8) ,
30353	 => std_logic_vector(to_unsigned(136,8) ,
30354	 => std_logic_vector(to_unsigned(73,8) ,
30355	 => std_logic_vector(to_unsigned(4,8) ,
30356	 => std_logic_vector(to_unsigned(1,8) ,
30357	 => std_logic_vector(to_unsigned(1,8) ,
30358	 => std_logic_vector(to_unsigned(6,8) ,
30359	 => std_logic_vector(to_unsigned(8,8) ,
30360	 => std_logic_vector(to_unsigned(5,8) ,
30361	 => std_logic_vector(to_unsigned(5,8) ,
30362	 => std_logic_vector(to_unsigned(5,8) ,
30363	 => std_logic_vector(to_unsigned(4,8) ,
30364	 => std_logic_vector(to_unsigned(4,8) ,
30365	 => std_logic_vector(to_unsigned(3,8) ,
30366	 => std_logic_vector(to_unsigned(2,8) ,
30367	 => std_logic_vector(to_unsigned(1,8) ,
30368	 => std_logic_vector(to_unsigned(1,8) ,
30369	 => std_logic_vector(to_unsigned(2,8) ,
30370	 => std_logic_vector(to_unsigned(6,8) ,
30371	 => std_logic_vector(to_unsigned(7,8) ,
30372	 => std_logic_vector(to_unsigned(3,8) ,
30373	 => std_logic_vector(to_unsigned(74,8) ,
30374	 => std_logic_vector(to_unsigned(127,8) ,
30375	 => std_logic_vector(to_unsigned(91,8) ,
30376	 => std_logic_vector(to_unsigned(142,8) ,
30377	 => std_logic_vector(to_unsigned(136,8) ,
30378	 => std_logic_vector(to_unsigned(118,8) ,
30379	 => std_logic_vector(to_unsigned(151,8) ,
30380	 => std_logic_vector(to_unsigned(171,8) ,
30381	 => std_logic_vector(to_unsigned(173,8) ,
30382	 => std_logic_vector(to_unsigned(171,8) ,
30383	 => std_logic_vector(to_unsigned(168,8) ,
30384	 => std_logic_vector(to_unsigned(161,8) ,
30385	 => std_logic_vector(to_unsigned(161,8) ,
30386	 => std_logic_vector(to_unsigned(157,8) ,
30387	 => std_logic_vector(to_unsigned(156,8) ,
30388	 => std_logic_vector(to_unsigned(159,8) ,
30389	 => std_logic_vector(to_unsigned(161,8) ,
30390	 => std_logic_vector(to_unsigned(157,8) ,
30391	 => std_logic_vector(to_unsigned(156,8) ,
30392	 => std_logic_vector(to_unsigned(157,8) ,
30393	 => std_logic_vector(to_unsigned(159,8) ,
30394	 => std_logic_vector(to_unsigned(157,8) ,
30395	 => std_logic_vector(to_unsigned(157,8) ,
30396	 => std_logic_vector(to_unsigned(154,8) ,
30397	 => std_logic_vector(to_unsigned(149,8) ,
30398	 => std_logic_vector(to_unsigned(149,8) ,
30399	 => std_logic_vector(to_unsigned(152,8) ,
30400	 => std_logic_vector(to_unsigned(156,8) ,
30401	 => std_logic_vector(to_unsigned(69,8) ,
30402	 => std_logic_vector(to_unsigned(82,8) ,
30403	 => std_logic_vector(to_unsigned(88,8) ,
30404	 => std_logic_vector(to_unsigned(118,8) ,
30405	 => std_logic_vector(to_unsigned(81,8) ,
30406	 => std_logic_vector(to_unsigned(11,8) ,
30407	 => std_logic_vector(to_unsigned(7,8) ,
30408	 => std_logic_vector(to_unsigned(7,8) ,
30409	 => std_logic_vector(to_unsigned(6,8) ,
30410	 => std_logic_vector(to_unsigned(4,8) ,
30411	 => std_logic_vector(to_unsigned(2,8) ,
30412	 => std_logic_vector(to_unsigned(2,8) ,
30413	 => std_logic_vector(to_unsigned(1,8) ,
30414	 => std_logic_vector(to_unsigned(0,8) ,
30415	 => std_logic_vector(to_unsigned(0,8) ,
30416	 => std_logic_vector(to_unsigned(0,8) ,
30417	 => std_logic_vector(to_unsigned(0,8) ,
30418	 => std_logic_vector(to_unsigned(0,8) ,
30419	 => std_logic_vector(to_unsigned(0,8) ,
30420	 => std_logic_vector(to_unsigned(0,8) ,
30421	 => std_logic_vector(to_unsigned(1,8) ,
30422	 => std_logic_vector(to_unsigned(3,8) ,
30423	 => std_logic_vector(to_unsigned(3,8) ,
30424	 => std_logic_vector(to_unsigned(3,8) ,
30425	 => std_logic_vector(to_unsigned(3,8) ,
30426	 => std_logic_vector(to_unsigned(4,8) ,
30427	 => std_logic_vector(to_unsigned(13,8) ,
30428	 => std_logic_vector(to_unsigned(21,8) ,
30429	 => std_logic_vector(to_unsigned(15,8) ,
30430	 => std_logic_vector(to_unsigned(12,8) ,
30431	 => std_logic_vector(to_unsigned(11,8) ,
30432	 => std_logic_vector(to_unsigned(9,8) ,
30433	 => std_logic_vector(to_unsigned(8,8) ,
30434	 => std_logic_vector(to_unsigned(5,8) ,
30435	 => std_logic_vector(to_unsigned(3,8) ,
30436	 => std_logic_vector(to_unsigned(3,8) ,
30437	 => std_logic_vector(to_unsigned(5,8) ,
30438	 => std_logic_vector(to_unsigned(4,8) ,
30439	 => std_logic_vector(to_unsigned(3,8) ,
30440	 => std_logic_vector(to_unsigned(10,8) ,
30441	 => std_logic_vector(to_unsigned(27,8) ,
30442	 => std_logic_vector(to_unsigned(29,8) ,
30443	 => std_logic_vector(to_unsigned(27,8) ,
30444	 => std_logic_vector(to_unsigned(27,8) ,
30445	 => std_logic_vector(to_unsigned(11,8) ,
30446	 => std_logic_vector(to_unsigned(6,8) ,
30447	 => std_logic_vector(to_unsigned(17,8) ,
30448	 => std_logic_vector(to_unsigned(51,8) ,
30449	 => std_logic_vector(to_unsigned(19,8) ,
30450	 => std_logic_vector(to_unsigned(6,8) ,
30451	 => std_logic_vector(to_unsigned(6,8) ,
30452	 => std_logic_vector(to_unsigned(2,8) ,
30453	 => std_logic_vector(to_unsigned(3,8) ,
30454	 => std_logic_vector(to_unsigned(2,8) ,
30455	 => std_logic_vector(to_unsigned(5,8) ,
30456	 => std_logic_vector(to_unsigned(18,8) ,
30457	 => std_logic_vector(to_unsigned(6,8) ,
30458	 => std_logic_vector(to_unsigned(9,8) ,
30459	 => std_logic_vector(to_unsigned(24,8) ,
30460	 => std_logic_vector(to_unsigned(31,8) ,
30461	 => std_logic_vector(to_unsigned(58,8) ,
30462	 => std_logic_vector(to_unsigned(88,8) ,
30463	 => std_logic_vector(to_unsigned(149,8) ,
30464	 => std_logic_vector(to_unsigned(86,8) ,
30465	 => std_logic_vector(to_unsigned(70,8) ,
30466	 => std_logic_vector(to_unsigned(157,8) ,
30467	 => std_logic_vector(to_unsigned(54,8) ,
30468	 => std_logic_vector(to_unsigned(15,8) ,
30469	 => std_logic_vector(to_unsigned(3,8) ,
30470	 => std_logic_vector(to_unsigned(1,8) ,
30471	 => std_logic_vector(to_unsigned(3,8) ,
30472	 => std_logic_vector(to_unsigned(8,8) ,
30473	 => std_logic_vector(to_unsigned(9,8) ,
30474	 => std_logic_vector(to_unsigned(15,8) ,
30475	 => std_logic_vector(to_unsigned(18,8) ,
30476	 => std_logic_vector(to_unsigned(20,8) ,
30477	 => std_logic_vector(to_unsigned(14,8) ,
30478	 => std_logic_vector(to_unsigned(7,8) ,
30479	 => std_logic_vector(to_unsigned(25,8) ,
30480	 => std_logic_vector(to_unsigned(131,8) ,
30481	 => std_logic_vector(to_unsigned(100,8) ,
30482	 => std_logic_vector(to_unsigned(74,8) ,
30483	 => std_logic_vector(to_unsigned(36,8) ,
30484	 => std_logic_vector(to_unsigned(24,8) ,
30485	 => std_logic_vector(to_unsigned(51,8) ,
30486	 => std_logic_vector(to_unsigned(67,8) ,
30487	 => std_logic_vector(to_unsigned(99,8) ,
30488	 => std_logic_vector(to_unsigned(141,8) ,
30489	 => std_logic_vector(to_unsigned(166,8) ,
30490	 => std_logic_vector(to_unsigned(175,8) ,
30491	 => std_logic_vector(to_unsigned(206,8) ,
30492	 => std_logic_vector(to_unsigned(64,8) ,
30493	 => std_logic_vector(to_unsigned(2,8) ,
30494	 => std_logic_vector(to_unsigned(18,8) ,
30495	 => std_logic_vector(to_unsigned(58,8) ,
30496	 => std_logic_vector(to_unsigned(47,8) ,
30497	 => std_logic_vector(to_unsigned(45,8) ,
30498	 => std_logic_vector(to_unsigned(59,8) ,
30499	 => std_logic_vector(to_unsigned(56,8) ,
30500	 => std_logic_vector(to_unsigned(41,8) ,
30501	 => std_logic_vector(to_unsigned(32,8) ,
30502	 => std_logic_vector(to_unsigned(25,8) ,
30503	 => std_logic_vector(to_unsigned(12,8) ,
30504	 => std_logic_vector(to_unsigned(2,8) ,
30505	 => std_logic_vector(to_unsigned(0,8) ,
30506	 => std_logic_vector(to_unsigned(5,8) ,
30507	 => std_logic_vector(to_unsigned(47,8) ,
30508	 => std_logic_vector(to_unsigned(65,8) ,
30509	 => std_logic_vector(to_unsigned(39,8) ,
30510	 => std_logic_vector(to_unsigned(18,8) ,
30511	 => std_logic_vector(to_unsigned(8,8) ,
30512	 => std_logic_vector(to_unsigned(2,8) ,
30513	 => std_logic_vector(to_unsigned(1,8) ,
30514	 => std_logic_vector(to_unsigned(1,8) ,
30515	 => std_logic_vector(to_unsigned(2,8) ,
30516	 => std_logic_vector(to_unsigned(1,8) ,
30517	 => std_logic_vector(to_unsigned(1,8) ,
30518	 => std_logic_vector(to_unsigned(1,8) ,
30519	 => std_logic_vector(to_unsigned(1,8) ,
30520	 => std_logic_vector(to_unsigned(1,8) ,
30521	 => std_logic_vector(to_unsigned(1,8) ,
30522	 => std_logic_vector(to_unsigned(1,8) ,
30523	 => std_logic_vector(to_unsigned(1,8) ,
30524	 => std_logic_vector(to_unsigned(1,8) ,
30525	 => std_logic_vector(to_unsigned(1,8) ,
30526	 => std_logic_vector(to_unsigned(1,8) ,
30527	 => std_logic_vector(to_unsigned(0,8) ,
30528	 => std_logic_vector(to_unsigned(2,8) ,
30529	 => std_logic_vector(to_unsigned(30,8) ,
30530	 => std_logic_vector(to_unsigned(74,8) ,
30531	 => std_logic_vector(to_unsigned(41,8) ,
30532	 => std_logic_vector(to_unsigned(34,8) ,
30533	 => std_logic_vector(to_unsigned(30,8) ,
30534	 => std_logic_vector(to_unsigned(23,8) ,
30535	 => std_logic_vector(to_unsigned(20,8) ,
30536	 => std_logic_vector(to_unsigned(17,8) ,
30537	 => std_logic_vector(to_unsigned(10,8) ,
30538	 => std_logic_vector(to_unsigned(12,8) ,
30539	 => std_logic_vector(to_unsigned(12,8) ,
30540	 => std_logic_vector(to_unsigned(56,8) ,
30541	 => std_logic_vector(to_unsigned(170,8) ,
30542	 => std_logic_vector(to_unsigned(164,8) ,
30543	 => std_logic_vector(to_unsigned(36,8) ,
30544	 => std_logic_vector(to_unsigned(1,8) ,
30545	 => std_logic_vector(to_unsigned(8,8) ,
30546	 => std_logic_vector(to_unsigned(5,8) ,
30547	 => std_logic_vector(to_unsigned(2,8) ,
30548	 => std_logic_vector(to_unsigned(9,8) ,
30549	 => std_logic_vector(to_unsigned(13,8) ,
30550	 => std_logic_vector(to_unsigned(5,8) ,
30551	 => std_logic_vector(to_unsigned(8,8) ,
30552	 => std_logic_vector(to_unsigned(38,8) ,
30553	 => std_logic_vector(to_unsigned(78,8) ,
30554	 => std_logic_vector(to_unsigned(99,8) ,
30555	 => std_logic_vector(to_unsigned(103,8) ,
30556	 => std_logic_vector(to_unsigned(73,8) ,
30557	 => std_logic_vector(to_unsigned(29,8) ,
30558	 => std_logic_vector(to_unsigned(44,8) ,
30559	 => std_logic_vector(to_unsigned(63,8) ,
30560	 => std_logic_vector(to_unsigned(18,8) ,
30561	 => std_logic_vector(to_unsigned(0,8) ,
30562	 => std_logic_vector(to_unsigned(4,8) ,
30563	 => std_logic_vector(to_unsigned(33,8) ,
30564	 => std_logic_vector(to_unsigned(68,8) ,
30565	 => std_logic_vector(to_unsigned(82,8) ,
30566	 => std_logic_vector(to_unsigned(84,8) ,
30567	 => std_logic_vector(to_unsigned(78,8) ,
30568	 => std_logic_vector(to_unsigned(108,8) ,
30569	 => std_logic_vector(to_unsigned(57,8) ,
30570	 => std_logic_vector(to_unsigned(20,8) ,
30571	 => std_logic_vector(to_unsigned(2,8) ,
30572	 => std_logic_vector(to_unsigned(0,8) ,
30573	 => std_logic_vector(to_unsigned(1,8) ,
30574	 => std_logic_vector(to_unsigned(2,8) ,
30575	 => std_logic_vector(to_unsigned(9,8) ,
30576	 => std_logic_vector(to_unsigned(74,8) ,
30577	 => std_logic_vector(to_unsigned(35,8) ,
30578	 => std_logic_vector(to_unsigned(8,8) ,
30579	 => std_logic_vector(to_unsigned(8,8) ,
30580	 => std_logic_vector(to_unsigned(8,8) ,
30581	 => std_logic_vector(to_unsigned(4,8) ,
30582	 => std_logic_vector(to_unsigned(5,8) ,
30583	 => std_logic_vector(to_unsigned(16,8) ,
30584	 => std_logic_vector(to_unsigned(45,8) ,
30585	 => std_logic_vector(to_unsigned(84,8) ,
30586	 => std_logic_vector(to_unsigned(139,8) ,
30587	 => std_logic_vector(to_unsigned(154,8) ,
30588	 => std_logic_vector(to_unsigned(146,8) ,
30589	 => std_logic_vector(to_unsigned(136,8) ,
30590	 => std_logic_vector(to_unsigned(136,8) ,
30591	 => std_logic_vector(to_unsigned(99,8) ,
30592	 => std_logic_vector(to_unsigned(82,8) ,
30593	 => std_logic_vector(to_unsigned(14,8) ,
30594	 => std_logic_vector(to_unsigned(5,8) ,
30595	 => std_logic_vector(to_unsigned(76,8) ,
30596	 => std_logic_vector(to_unsigned(131,8) ,
30597	 => std_logic_vector(to_unsigned(147,8) ,
30598	 => std_logic_vector(to_unsigned(151,8) ,
30599	 => std_logic_vector(to_unsigned(134,8) ,
30600	 => std_logic_vector(to_unsigned(147,8) ,
30601	 => std_logic_vector(to_unsigned(154,8) ,
30602	 => std_logic_vector(to_unsigned(92,8) ,
30603	 => std_logic_vector(to_unsigned(40,8) ,
30604	 => std_logic_vector(to_unsigned(42,8) ,
30605	 => std_logic_vector(to_unsigned(45,8) ,
30606	 => std_logic_vector(to_unsigned(35,8) ,
30607	 => std_logic_vector(to_unsigned(8,8) ,
30608	 => std_logic_vector(to_unsigned(14,8) ,
30609	 => std_logic_vector(to_unsigned(85,8) ,
30610	 => std_logic_vector(to_unsigned(119,8) ,
30611	 => std_logic_vector(to_unsigned(154,8) ,
30612	 => std_logic_vector(to_unsigned(154,8) ,
30613	 => std_logic_vector(to_unsigned(156,8) ,
30614	 => std_logic_vector(to_unsigned(156,8) ,
30615	 => std_logic_vector(to_unsigned(152,8) ,
30616	 => std_logic_vector(to_unsigned(156,8) ,
30617	 => std_logic_vector(to_unsigned(151,8) ,
30618	 => std_logic_vector(to_unsigned(154,8) ,
30619	 => std_logic_vector(to_unsigned(163,8) ,
30620	 => std_logic_vector(to_unsigned(179,8) ,
30621	 => std_logic_vector(to_unsigned(173,8) ,
30622	 => std_logic_vector(to_unsigned(146,8) ,
30623	 => std_logic_vector(to_unsigned(139,8) ,
30624	 => std_logic_vector(to_unsigned(104,8) ,
30625	 => std_logic_vector(to_unsigned(96,8) ,
30626	 => std_logic_vector(to_unsigned(124,8) ,
30627	 => std_logic_vector(to_unsigned(131,8) ,
30628	 => std_logic_vector(to_unsigned(130,8) ,
30629	 => std_logic_vector(to_unsigned(127,8) ,
30630	 => std_logic_vector(to_unsigned(116,8) ,
30631	 => std_logic_vector(to_unsigned(95,8) ,
30632	 => std_logic_vector(to_unsigned(65,8) ,
30633	 => std_logic_vector(to_unsigned(37,8) ,
30634	 => std_logic_vector(to_unsigned(12,8) ,
30635	 => std_logic_vector(to_unsigned(20,8) ,
30636	 => std_logic_vector(to_unsigned(51,8) ,
30637	 => std_logic_vector(to_unsigned(59,8) ,
30638	 => std_logic_vector(to_unsigned(39,8) ,
30639	 => std_logic_vector(to_unsigned(4,8) ,
30640	 => std_logic_vector(to_unsigned(1,8) ,
30641	 => std_logic_vector(to_unsigned(11,8) ,
30642	 => std_logic_vector(to_unsigned(16,8) ,
30643	 => std_logic_vector(to_unsigned(25,8) ,
30644	 => std_logic_vector(to_unsigned(25,8) ,
30645	 => std_logic_vector(to_unsigned(17,8) ,
30646	 => std_logic_vector(to_unsigned(12,8) ,
30647	 => std_logic_vector(to_unsigned(5,8) ,
30648	 => std_logic_vector(to_unsigned(1,8) ,
30649	 => std_logic_vector(to_unsigned(2,8) ,
30650	 => std_logic_vector(to_unsigned(3,8) ,
30651	 => std_logic_vector(to_unsigned(2,8) ,
30652	 => std_logic_vector(to_unsigned(2,8) ,
30653	 => std_logic_vector(to_unsigned(2,8) ,
30654	 => std_logic_vector(to_unsigned(3,8) ,
30655	 => std_logic_vector(to_unsigned(3,8) ,
30656	 => std_logic_vector(to_unsigned(2,8) ,
30657	 => std_logic_vector(to_unsigned(9,8) ,
30658	 => std_logic_vector(to_unsigned(13,8) ,
30659	 => std_logic_vector(to_unsigned(6,8) ,
30660	 => std_logic_vector(to_unsigned(2,8) ,
30661	 => std_logic_vector(to_unsigned(4,8) ,
30662	 => std_logic_vector(to_unsigned(6,8) ,
30663	 => std_logic_vector(to_unsigned(14,8) ,
30664	 => std_logic_vector(to_unsigned(38,8) ,
30665	 => std_logic_vector(to_unsigned(49,8) ,
30666	 => std_logic_vector(to_unsigned(43,8) ,
30667	 => std_logic_vector(to_unsigned(48,8) ,
30668	 => std_logic_vector(to_unsigned(60,8) ,
30669	 => std_logic_vector(to_unsigned(27,8) ,
30670	 => std_logic_vector(to_unsigned(57,8) ,
30671	 => std_logic_vector(to_unsigned(109,8) ,
30672	 => std_logic_vector(to_unsigned(142,8) ,
30673	 => std_logic_vector(to_unsigned(131,8) ,
30674	 => std_logic_vector(to_unsigned(69,8) ,
30675	 => std_logic_vector(to_unsigned(7,8) ,
30676	 => std_logic_vector(to_unsigned(1,8) ,
30677	 => std_logic_vector(to_unsigned(3,8) ,
30678	 => std_logic_vector(to_unsigned(7,8) ,
30679	 => std_logic_vector(to_unsigned(8,8) ,
30680	 => std_logic_vector(to_unsigned(5,8) ,
30681	 => std_logic_vector(to_unsigned(4,8) ,
30682	 => std_logic_vector(to_unsigned(4,8) ,
30683	 => std_logic_vector(to_unsigned(4,8) ,
30684	 => std_logic_vector(to_unsigned(3,8) ,
30685	 => std_logic_vector(to_unsigned(3,8) ,
30686	 => std_logic_vector(to_unsigned(3,8) ,
30687	 => std_logic_vector(to_unsigned(1,8) ,
30688	 => std_logic_vector(to_unsigned(1,8) ,
30689	 => std_logic_vector(to_unsigned(1,8) ,
30690	 => std_logic_vector(to_unsigned(32,8) ,
30691	 => std_logic_vector(to_unsigned(17,8) ,
30692	 => std_logic_vector(to_unsigned(0,8) ,
30693	 => std_logic_vector(to_unsigned(34,8) ,
30694	 => std_logic_vector(to_unsigned(99,8) ,
30695	 => std_logic_vector(to_unsigned(51,8) ,
30696	 => std_logic_vector(to_unsigned(64,8) ,
30697	 => std_logic_vector(to_unsigned(71,8) ,
30698	 => std_logic_vector(to_unsigned(69,8) ,
30699	 => std_logic_vector(to_unsigned(91,8) ,
30700	 => std_logic_vector(to_unsigned(125,8) ,
30701	 => std_logic_vector(to_unsigned(170,8) ,
30702	 => std_logic_vector(to_unsigned(177,8) ,
30703	 => std_logic_vector(to_unsigned(159,8) ,
30704	 => std_logic_vector(to_unsigned(161,8) ,
30705	 => std_logic_vector(to_unsigned(161,8) ,
30706	 => std_logic_vector(to_unsigned(161,8) ,
30707	 => std_logic_vector(to_unsigned(156,8) ,
30708	 => std_logic_vector(to_unsigned(157,8) ,
30709	 => std_logic_vector(to_unsigned(161,8) ,
30710	 => std_logic_vector(to_unsigned(159,8) ,
30711	 => std_logic_vector(to_unsigned(156,8) ,
30712	 => std_logic_vector(to_unsigned(159,8) ,
30713	 => std_logic_vector(to_unsigned(157,8) ,
30714	 => std_logic_vector(to_unsigned(156,8) ,
30715	 => std_logic_vector(to_unsigned(156,8) ,
30716	 => std_logic_vector(to_unsigned(154,8) ,
30717	 => std_logic_vector(to_unsigned(151,8) ,
30718	 => std_logic_vector(to_unsigned(151,8) ,
30719	 => std_logic_vector(to_unsigned(156,8) ,
30720	 => std_logic_vector(to_unsigned(159,8) ,
30721	 => std_logic_vector(to_unsigned(1,8) ,
30722	 => std_logic_vector(to_unsigned(2,8) ,
30723	 => std_logic_vector(to_unsigned(2,8) ,
30724	 => std_logic_vector(to_unsigned(4,8) ,
30725	 => std_logic_vector(to_unsigned(8,8) ,
30726	 => std_logic_vector(to_unsigned(8,8) ,
30727	 => std_logic_vector(to_unsigned(9,8) ,
30728	 => std_logic_vector(to_unsigned(8,8) ,
30729	 => std_logic_vector(to_unsigned(6,8) ,
30730	 => std_logic_vector(to_unsigned(2,8) ,
30731	 => std_logic_vector(to_unsigned(2,8) ,
30732	 => std_logic_vector(to_unsigned(1,8) ,
30733	 => std_logic_vector(to_unsigned(0,8) ,
30734	 => std_logic_vector(to_unsigned(0,8) ,
30735	 => std_logic_vector(to_unsigned(0,8) ,
30736	 => std_logic_vector(to_unsigned(0,8) ,
30737	 => std_logic_vector(to_unsigned(1,8) ,
30738	 => std_logic_vector(to_unsigned(0,8) ,
30739	 => std_logic_vector(to_unsigned(0,8) ,
30740	 => std_logic_vector(to_unsigned(2,8) ,
30741	 => std_logic_vector(to_unsigned(8,8) ,
30742	 => std_logic_vector(to_unsigned(8,8) ,
30743	 => std_logic_vector(to_unsigned(9,8) ,
30744	 => std_logic_vector(to_unsigned(4,8) ,
30745	 => std_logic_vector(to_unsigned(2,8) ,
30746	 => std_logic_vector(to_unsigned(15,8) ,
30747	 => std_logic_vector(to_unsigned(38,8) ,
30748	 => std_logic_vector(to_unsigned(30,8) ,
30749	 => std_logic_vector(to_unsigned(17,8) ,
30750	 => std_logic_vector(to_unsigned(7,8) ,
30751	 => std_logic_vector(to_unsigned(8,8) ,
30752	 => std_logic_vector(to_unsigned(8,8) ,
30753	 => std_logic_vector(to_unsigned(8,8) ,
30754	 => std_logic_vector(to_unsigned(7,8) ,
30755	 => std_logic_vector(to_unsigned(5,8) ,
30756	 => std_logic_vector(to_unsigned(3,8) ,
30757	 => std_logic_vector(to_unsigned(1,8) ,
30758	 => std_logic_vector(to_unsigned(2,8) ,
30759	 => std_logic_vector(to_unsigned(19,8) ,
30760	 => std_logic_vector(to_unsigned(43,8) ,
30761	 => std_logic_vector(to_unsigned(36,8) ,
30762	 => std_logic_vector(to_unsigned(27,8) ,
30763	 => std_logic_vector(to_unsigned(18,8) ,
30764	 => std_logic_vector(to_unsigned(15,8) ,
30765	 => std_logic_vector(to_unsigned(14,8) ,
30766	 => std_logic_vector(to_unsigned(10,8) ,
30767	 => std_logic_vector(to_unsigned(3,8) ,
30768	 => std_logic_vector(to_unsigned(4,8) ,
30769	 => std_logic_vector(to_unsigned(4,8) ,
30770	 => std_logic_vector(to_unsigned(2,8) ,
30771	 => std_logic_vector(to_unsigned(2,8) ,
30772	 => std_logic_vector(to_unsigned(3,8) ,
30773	 => std_logic_vector(to_unsigned(2,8) ,
30774	 => std_logic_vector(to_unsigned(1,8) ,
30775	 => std_logic_vector(to_unsigned(29,8) ,
30776	 => std_logic_vector(to_unsigned(76,8) ,
30777	 => std_logic_vector(to_unsigned(23,8) ,
30778	 => std_logic_vector(to_unsigned(11,8) ,
30779	 => std_logic_vector(to_unsigned(29,8) ,
30780	 => std_logic_vector(to_unsigned(55,8) ,
30781	 => std_logic_vector(to_unsigned(39,8) ,
30782	 => std_logic_vector(to_unsigned(55,8) ,
30783	 => std_logic_vector(to_unsigned(90,8) ,
30784	 => std_logic_vector(to_unsigned(51,8) ,
30785	 => std_logic_vector(to_unsigned(103,8) ,
30786	 => std_logic_vector(to_unsigned(168,8) ,
30787	 => std_logic_vector(to_unsigned(70,8) ,
30788	 => std_logic_vector(to_unsigned(14,8) ,
30789	 => std_logic_vector(to_unsigned(27,8) ,
30790	 => std_logic_vector(to_unsigned(8,8) ,
30791	 => std_logic_vector(to_unsigned(3,8) ,
30792	 => std_logic_vector(to_unsigned(3,8) ,
30793	 => std_logic_vector(to_unsigned(4,8) ,
30794	 => std_logic_vector(to_unsigned(22,8) ,
30795	 => std_logic_vector(to_unsigned(38,8) ,
30796	 => std_logic_vector(to_unsigned(27,8) ,
30797	 => std_logic_vector(to_unsigned(16,8) ,
30798	 => std_logic_vector(to_unsigned(11,8) ,
30799	 => std_logic_vector(to_unsigned(7,8) ,
30800	 => std_logic_vector(to_unsigned(59,8) ,
30801	 => std_logic_vector(to_unsigned(119,8) ,
30802	 => std_logic_vector(to_unsigned(104,8) ,
30803	 => std_logic_vector(to_unsigned(69,8) ,
30804	 => std_logic_vector(to_unsigned(24,8) ,
30805	 => std_logic_vector(to_unsigned(37,8) ,
30806	 => std_logic_vector(to_unsigned(12,8) ,
30807	 => std_logic_vector(to_unsigned(16,8) ,
30808	 => std_logic_vector(to_unsigned(66,8) ,
30809	 => std_logic_vector(to_unsigned(71,8) ,
30810	 => std_logic_vector(to_unsigned(62,8) ,
30811	 => std_logic_vector(to_unsigned(124,8) ,
30812	 => std_logic_vector(to_unsigned(97,8) ,
30813	 => std_logic_vector(to_unsigned(29,8) ,
30814	 => std_logic_vector(to_unsigned(67,8) ,
30815	 => std_logic_vector(to_unsigned(76,8) ,
30816	 => std_logic_vector(to_unsigned(28,8) ,
30817	 => std_logic_vector(to_unsigned(15,8) ,
30818	 => std_logic_vector(to_unsigned(41,8) ,
30819	 => std_logic_vector(to_unsigned(37,8) ,
30820	 => std_logic_vector(to_unsigned(14,8) ,
30821	 => std_logic_vector(to_unsigned(14,8) ,
30822	 => std_logic_vector(to_unsigned(9,8) ,
30823	 => std_logic_vector(to_unsigned(1,8) ,
30824	 => std_logic_vector(to_unsigned(0,8) ,
30825	 => std_logic_vector(to_unsigned(0,8) ,
30826	 => std_logic_vector(to_unsigned(9,8) ,
30827	 => std_logic_vector(to_unsigned(53,8) ,
30828	 => std_logic_vector(to_unsigned(72,8) ,
30829	 => std_logic_vector(to_unsigned(55,8) ,
30830	 => std_logic_vector(to_unsigned(36,8) ,
30831	 => std_logic_vector(to_unsigned(12,8) ,
30832	 => std_logic_vector(to_unsigned(1,8) ,
30833	 => std_logic_vector(to_unsigned(1,8) ,
30834	 => std_logic_vector(to_unsigned(1,8) ,
30835	 => std_logic_vector(to_unsigned(1,8) ,
30836	 => std_logic_vector(to_unsigned(2,8) ,
30837	 => std_logic_vector(to_unsigned(1,8) ,
30838	 => std_logic_vector(to_unsigned(0,8) ,
30839	 => std_logic_vector(to_unsigned(1,8) ,
30840	 => std_logic_vector(to_unsigned(4,8) ,
30841	 => std_logic_vector(to_unsigned(4,8) ,
30842	 => std_logic_vector(to_unsigned(2,8) ,
30843	 => std_logic_vector(to_unsigned(2,8) ,
30844	 => std_logic_vector(to_unsigned(2,8) ,
30845	 => std_logic_vector(to_unsigned(1,8) ,
30846	 => std_logic_vector(to_unsigned(3,8) ,
30847	 => std_logic_vector(to_unsigned(9,8) ,
30848	 => std_logic_vector(to_unsigned(37,8) ,
30849	 => std_logic_vector(to_unsigned(78,8) ,
30850	 => std_logic_vector(to_unsigned(60,8) ,
30851	 => std_logic_vector(to_unsigned(51,8) ,
30852	 => std_logic_vector(to_unsigned(33,8) ,
30853	 => std_logic_vector(to_unsigned(15,8) ,
30854	 => std_logic_vector(to_unsigned(22,8) ,
30855	 => std_logic_vector(to_unsigned(18,8) ,
30856	 => std_logic_vector(to_unsigned(12,8) ,
30857	 => std_logic_vector(to_unsigned(28,8) ,
30858	 => std_logic_vector(to_unsigned(13,8) ,
30859	 => std_logic_vector(to_unsigned(7,8) ,
30860	 => std_logic_vector(to_unsigned(84,8) ,
30861	 => std_logic_vector(to_unsigned(184,8) ,
30862	 => std_logic_vector(to_unsigned(192,8) ,
30863	 => std_logic_vector(to_unsigned(138,8) ,
30864	 => std_logic_vector(to_unsigned(7,8) ,
30865	 => std_logic_vector(to_unsigned(3,8) ,
30866	 => std_logic_vector(to_unsigned(3,8) ,
30867	 => std_logic_vector(to_unsigned(1,8) ,
30868	 => std_logic_vector(to_unsigned(2,8) ,
30869	 => std_logic_vector(to_unsigned(3,8) ,
30870	 => std_logic_vector(to_unsigned(9,8) ,
30871	 => std_logic_vector(to_unsigned(34,8) ,
30872	 => std_logic_vector(to_unsigned(77,8) ,
30873	 => std_logic_vector(to_unsigned(81,8) ,
30874	 => std_logic_vector(to_unsigned(84,8) ,
30875	 => std_logic_vector(to_unsigned(72,8) ,
30876	 => std_logic_vector(to_unsigned(80,8) ,
30877	 => std_logic_vector(to_unsigned(97,8) ,
30878	 => std_logic_vector(to_unsigned(79,8) ,
30879	 => std_logic_vector(to_unsigned(71,8) ,
30880	 => std_logic_vector(to_unsigned(23,8) ,
30881	 => std_logic_vector(to_unsigned(2,8) ,
30882	 => std_logic_vector(to_unsigned(2,8) ,
30883	 => std_logic_vector(to_unsigned(28,8) ,
30884	 => std_logic_vector(to_unsigned(79,8) ,
30885	 => std_logic_vector(to_unsigned(95,8) ,
30886	 => std_logic_vector(to_unsigned(104,8) ,
30887	 => std_logic_vector(to_unsigned(104,8) ,
30888	 => std_logic_vector(to_unsigned(57,8) ,
30889	 => std_logic_vector(to_unsigned(3,8) ,
30890	 => std_logic_vector(to_unsigned(1,8) ,
30891	 => std_logic_vector(to_unsigned(16,8) ,
30892	 => std_logic_vector(to_unsigned(30,8) ,
30893	 => std_logic_vector(to_unsigned(8,8) ,
30894	 => std_logic_vector(to_unsigned(17,8) ,
30895	 => std_logic_vector(to_unsigned(59,8) ,
30896	 => std_logic_vector(to_unsigned(133,8) ,
30897	 => std_logic_vector(to_unsigned(107,8) ,
30898	 => std_logic_vector(to_unsigned(100,8) ,
30899	 => std_logic_vector(to_unsigned(51,8) ,
30900	 => std_logic_vector(to_unsigned(3,8) ,
30901	 => std_logic_vector(to_unsigned(4,8) ,
30902	 => std_logic_vector(to_unsigned(38,8) ,
30903	 => std_logic_vector(to_unsigned(91,8) ,
30904	 => std_logic_vector(to_unsigned(65,8) ,
30905	 => std_logic_vector(to_unsigned(68,8) ,
30906	 => std_logic_vector(to_unsigned(130,8) ,
30907	 => std_logic_vector(to_unsigned(130,8) ,
30908	 => std_logic_vector(to_unsigned(121,8) ,
30909	 => std_logic_vector(to_unsigned(124,8) ,
30910	 => std_logic_vector(to_unsigned(125,8) ,
30911	 => std_logic_vector(to_unsigned(72,8) ,
30912	 => std_logic_vector(to_unsigned(109,8) ,
30913	 => std_logic_vector(to_unsigned(58,8) ,
30914	 => std_logic_vector(to_unsigned(57,8) ,
30915	 => std_logic_vector(to_unsigned(157,8) ,
30916	 => std_logic_vector(to_unsigned(161,8) ,
30917	 => std_logic_vector(to_unsigned(157,8) ,
30918	 => std_logic_vector(to_unsigned(156,8) ,
30919	 => std_logic_vector(to_unsigned(142,8) ,
30920	 => std_logic_vector(to_unsigned(144,8) ,
30921	 => std_logic_vector(to_unsigned(147,8) ,
30922	 => std_logic_vector(to_unsigned(112,8) ,
30923	 => std_logic_vector(to_unsigned(58,8) ,
30924	 => std_logic_vector(to_unsigned(27,8) ,
30925	 => std_logic_vector(to_unsigned(23,8) ,
30926	 => std_logic_vector(to_unsigned(32,8) ,
30927	 => std_logic_vector(to_unsigned(13,8) ,
30928	 => std_logic_vector(to_unsigned(14,8) ,
30929	 => std_logic_vector(to_unsigned(101,8) ,
30930	 => std_logic_vector(to_unsigned(144,8) ,
30931	 => std_logic_vector(to_unsigned(159,8) ,
30932	 => std_logic_vector(to_unsigned(156,8) ,
30933	 => std_logic_vector(to_unsigned(152,8) ,
30934	 => std_logic_vector(to_unsigned(152,8) ,
30935	 => std_logic_vector(to_unsigned(157,8) ,
30936	 => std_logic_vector(to_unsigned(151,8) ,
30937	 => std_logic_vector(to_unsigned(152,8) ,
30938	 => std_logic_vector(to_unsigned(154,8) ,
30939	 => std_logic_vector(to_unsigned(154,8) ,
30940	 => std_logic_vector(to_unsigned(151,8) ,
30941	 => std_logic_vector(to_unsigned(154,8) ,
30942	 => std_logic_vector(to_unsigned(161,8) ,
30943	 => std_logic_vector(to_unsigned(159,8) ,
30944	 => std_logic_vector(to_unsigned(138,8) ,
30945	 => std_logic_vector(to_unsigned(115,8) ,
30946	 => std_logic_vector(to_unsigned(121,8) ,
30947	 => std_logic_vector(to_unsigned(128,8) ,
30948	 => std_logic_vector(to_unsigned(134,8) ,
30949	 => std_logic_vector(to_unsigned(128,8) ,
30950	 => std_logic_vector(to_unsigned(118,8) ,
30951	 => std_logic_vector(to_unsigned(96,8) ,
30952	 => std_logic_vector(to_unsigned(63,8) ,
30953	 => std_logic_vector(to_unsigned(44,8) ,
30954	 => std_logic_vector(to_unsigned(23,8) ,
30955	 => std_logic_vector(to_unsigned(24,8) ,
30956	 => std_logic_vector(to_unsigned(47,8) ,
30957	 => std_logic_vector(to_unsigned(47,8) ,
30958	 => std_logic_vector(to_unsigned(27,8) ,
30959	 => std_logic_vector(to_unsigned(4,8) ,
30960	 => std_logic_vector(to_unsigned(2,8) ,
30961	 => std_logic_vector(to_unsigned(10,8) ,
30962	 => std_logic_vector(to_unsigned(16,8) ,
30963	 => std_logic_vector(to_unsigned(27,8) ,
30964	 => std_logic_vector(to_unsigned(26,8) ,
30965	 => std_logic_vector(to_unsigned(17,8) ,
30966	 => std_logic_vector(to_unsigned(9,8) ,
30967	 => std_logic_vector(to_unsigned(3,8) ,
30968	 => std_logic_vector(to_unsigned(1,8) ,
30969	 => std_logic_vector(to_unsigned(2,8) ,
30970	 => std_logic_vector(to_unsigned(3,8) ,
30971	 => std_logic_vector(to_unsigned(2,8) ,
30972	 => std_logic_vector(to_unsigned(2,8) ,
30973	 => std_logic_vector(to_unsigned(2,8) ,
30974	 => std_logic_vector(to_unsigned(2,8) ,
30975	 => std_logic_vector(to_unsigned(3,8) ,
30976	 => std_logic_vector(to_unsigned(4,8) ,
30977	 => std_logic_vector(to_unsigned(3,8) ,
30978	 => std_logic_vector(to_unsigned(3,8) ,
30979	 => std_logic_vector(to_unsigned(6,8) ,
30980	 => std_logic_vector(to_unsigned(14,8) ,
30981	 => std_logic_vector(to_unsigned(14,8) ,
30982	 => std_logic_vector(to_unsigned(5,8) ,
30983	 => std_logic_vector(to_unsigned(21,8) ,
30984	 => std_logic_vector(to_unsigned(68,8) ,
30985	 => std_logic_vector(to_unsigned(51,8) ,
30986	 => std_logic_vector(to_unsigned(59,8) ,
30987	 => std_logic_vector(to_unsigned(92,8) ,
30988	 => std_logic_vector(to_unsigned(71,8) ,
30989	 => std_logic_vector(to_unsigned(53,8) ,
30990	 => std_logic_vector(to_unsigned(55,8) ,
30991	 => std_logic_vector(to_unsigned(108,8) ,
30992	 => std_logic_vector(to_unsigned(87,8) ,
30993	 => std_logic_vector(to_unsigned(25,8) ,
30994	 => std_logic_vector(to_unsigned(5,8) ,
30995	 => std_logic_vector(to_unsigned(2,8) ,
30996	 => std_logic_vector(to_unsigned(3,8) ,
30997	 => std_logic_vector(to_unsigned(5,8) ,
30998	 => std_logic_vector(to_unsigned(4,8) ,
30999	 => std_logic_vector(to_unsigned(2,8) ,
31000	 => std_logic_vector(to_unsigned(4,8) ,
31001	 => std_logic_vector(to_unsigned(6,8) ,
31002	 => std_logic_vector(to_unsigned(5,8) ,
31003	 => std_logic_vector(to_unsigned(4,8) ,
31004	 => std_logic_vector(to_unsigned(3,8) ,
31005	 => std_logic_vector(to_unsigned(4,8) ,
31006	 => std_logic_vector(to_unsigned(2,8) ,
31007	 => std_logic_vector(to_unsigned(1,8) ,
31008	 => std_logic_vector(to_unsigned(0,8) ,
31009	 => std_logic_vector(to_unsigned(0,8) ,
31010	 => std_logic_vector(to_unsigned(23,8) ,
31011	 => std_logic_vector(to_unsigned(19,8) ,
31012	 => std_logic_vector(to_unsigned(1,8) ,
31013	 => std_logic_vector(to_unsigned(6,8) ,
31014	 => std_logic_vector(to_unsigned(22,8) ,
31015	 => std_logic_vector(to_unsigned(29,8) ,
31016	 => std_logic_vector(to_unsigned(76,8) ,
31017	 => std_logic_vector(to_unsigned(99,8) ,
31018	 => std_logic_vector(to_unsigned(81,8) ,
31019	 => std_logic_vector(to_unsigned(109,8) ,
31020	 => std_logic_vector(to_unsigned(156,8) ,
31021	 => std_logic_vector(to_unsigned(161,8) ,
31022	 => std_logic_vector(to_unsigned(157,8) ,
31023	 => std_logic_vector(to_unsigned(161,8) ,
31024	 => std_logic_vector(to_unsigned(159,8) ,
31025	 => std_logic_vector(to_unsigned(159,8) ,
31026	 => std_logic_vector(to_unsigned(159,8) ,
31027	 => std_logic_vector(to_unsigned(156,8) ,
31028	 => std_logic_vector(to_unsigned(156,8) ,
31029	 => std_logic_vector(to_unsigned(156,8) ,
31030	 => std_logic_vector(to_unsigned(156,8) ,
31031	 => std_logic_vector(to_unsigned(156,8) ,
31032	 => std_logic_vector(to_unsigned(159,8) ,
31033	 => std_logic_vector(to_unsigned(157,8) ,
31034	 => std_logic_vector(to_unsigned(156,8) ,
31035	 => std_logic_vector(to_unsigned(156,8) ,
31036	 => std_logic_vector(to_unsigned(154,8) ,
31037	 => std_logic_vector(to_unsigned(149,8) ,
31038	 => std_logic_vector(to_unsigned(149,8) ,
31039	 => std_logic_vector(to_unsigned(149,8) ,
31040	 => std_logic_vector(to_unsigned(146,8) ,
31041	 => std_logic_vector(to_unsigned(1,8) ,
31042	 => std_logic_vector(to_unsigned(1,8) ,
31043	 => std_logic_vector(to_unsigned(1,8) ,
31044	 => std_logic_vector(to_unsigned(1,8) ,
31045	 => std_logic_vector(to_unsigned(9,8) ,
31046	 => std_logic_vector(to_unsigned(16,8) ,
31047	 => std_logic_vector(to_unsigned(10,8) ,
31048	 => std_logic_vector(to_unsigned(6,8) ,
31049	 => std_logic_vector(to_unsigned(4,8) ,
31050	 => std_logic_vector(to_unsigned(2,8) ,
31051	 => std_logic_vector(to_unsigned(1,8) ,
31052	 => std_logic_vector(to_unsigned(1,8) ,
31053	 => std_logic_vector(to_unsigned(0,8) ,
31054	 => std_logic_vector(to_unsigned(0,8) ,
31055	 => std_logic_vector(to_unsigned(0,8) ,
31056	 => std_logic_vector(to_unsigned(0,8) ,
31057	 => std_logic_vector(to_unsigned(0,8) ,
31058	 => std_logic_vector(to_unsigned(1,8) ,
31059	 => std_logic_vector(to_unsigned(2,8) ,
31060	 => std_logic_vector(to_unsigned(13,8) ,
31061	 => std_logic_vector(to_unsigned(15,8) ,
31062	 => std_logic_vector(to_unsigned(8,8) ,
31063	 => std_logic_vector(to_unsigned(12,8) ,
31064	 => std_logic_vector(to_unsigned(4,8) ,
31065	 => std_logic_vector(to_unsigned(10,8) ,
31066	 => std_logic_vector(to_unsigned(45,8) ,
31067	 => std_logic_vector(to_unsigned(29,8) ,
31068	 => std_logic_vector(to_unsigned(23,8) ,
31069	 => std_logic_vector(to_unsigned(28,8) ,
31070	 => std_logic_vector(to_unsigned(15,8) ,
31071	 => std_logic_vector(to_unsigned(17,8) ,
31072	 => std_logic_vector(to_unsigned(16,8) ,
31073	 => std_logic_vector(to_unsigned(14,8) ,
31074	 => std_logic_vector(to_unsigned(16,8) ,
31075	 => std_logic_vector(to_unsigned(12,8) ,
31076	 => std_logic_vector(to_unsigned(6,8) ,
31077	 => std_logic_vector(to_unsigned(2,8) ,
31078	 => std_logic_vector(to_unsigned(19,8) ,
31079	 => std_logic_vector(to_unsigned(52,8) ,
31080	 => std_logic_vector(to_unsigned(34,8) ,
31081	 => std_logic_vector(to_unsigned(19,8) ,
31082	 => std_logic_vector(to_unsigned(12,8) ,
31083	 => std_logic_vector(to_unsigned(8,8) ,
31084	 => std_logic_vector(to_unsigned(6,8) ,
31085	 => std_logic_vector(to_unsigned(5,8) ,
31086	 => std_logic_vector(to_unsigned(4,8) ,
31087	 => std_logic_vector(to_unsigned(6,8) ,
31088	 => std_logic_vector(to_unsigned(3,8) ,
31089	 => std_logic_vector(to_unsigned(2,8) ,
31090	 => std_logic_vector(to_unsigned(3,8) ,
31091	 => std_logic_vector(to_unsigned(1,8) ,
31092	 => std_logic_vector(to_unsigned(0,8) ,
31093	 => std_logic_vector(to_unsigned(0,8) ,
31094	 => std_logic_vector(to_unsigned(4,8) ,
31095	 => std_logic_vector(to_unsigned(58,8) ,
31096	 => std_logic_vector(to_unsigned(56,8) ,
31097	 => std_logic_vector(to_unsigned(37,8) ,
31098	 => std_logic_vector(to_unsigned(22,8) ,
31099	 => std_logic_vector(to_unsigned(17,8) ,
31100	 => std_logic_vector(to_unsigned(32,8) ,
31101	 => std_logic_vector(to_unsigned(61,8) ,
31102	 => std_logic_vector(to_unsigned(116,8) ,
31103	 => std_logic_vector(to_unsigned(32,8) ,
31104	 => std_logic_vector(to_unsigned(18,8) ,
31105	 => std_logic_vector(to_unsigned(112,8) ,
31106	 => std_logic_vector(to_unsigned(131,8) ,
31107	 => std_logic_vector(to_unsigned(101,8) ,
31108	 => std_logic_vector(to_unsigned(8,8) ,
31109	 => std_logic_vector(to_unsigned(6,8) ,
31110	 => std_logic_vector(to_unsigned(16,8) ,
31111	 => std_logic_vector(to_unsigned(9,8) ,
31112	 => std_logic_vector(to_unsigned(3,8) ,
31113	 => std_logic_vector(to_unsigned(7,8) ,
31114	 => std_logic_vector(to_unsigned(23,8) ,
31115	 => std_logic_vector(to_unsigned(29,8) ,
31116	 => std_logic_vector(to_unsigned(31,8) ,
31117	 => std_logic_vector(to_unsigned(18,8) ,
31118	 => std_logic_vector(to_unsigned(12,8) ,
31119	 => std_logic_vector(to_unsigned(5,8) ,
31120	 => std_logic_vector(to_unsigned(29,8) ,
31121	 => std_logic_vector(to_unsigned(142,8) ,
31122	 => std_logic_vector(to_unsigned(134,8) ,
31123	 => std_logic_vector(to_unsigned(136,8) ,
31124	 => std_logic_vector(to_unsigned(119,8) ,
31125	 => std_logic_vector(to_unsigned(107,8) ,
31126	 => std_logic_vector(to_unsigned(51,8) ,
31127	 => std_logic_vector(to_unsigned(40,8) ,
31128	 => std_logic_vector(to_unsigned(90,8) ,
31129	 => std_logic_vector(to_unsigned(51,8) ,
31130	 => std_logic_vector(to_unsigned(39,8) ,
31131	 => std_logic_vector(to_unsigned(47,8) ,
31132	 => std_logic_vector(to_unsigned(61,8) ,
31133	 => std_logic_vector(to_unsigned(70,8) ,
31134	 => std_logic_vector(to_unsigned(49,8) ,
31135	 => std_logic_vector(to_unsigned(21,8) ,
31136	 => std_logic_vector(to_unsigned(5,8) ,
31137	 => std_logic_vector(to_unsigned(9,8) ,
31138	 => std_logic_vector(to_unsigned(20,8) ,
31139	 => std_logic_vector(to_unsigned(6,8) ,
31140	 => std_logic_vector(to_unsigned(2,8) ,
31141	 => std_logic_vector(to_unsigned(5,8) ,
31142	 => std_logic_vector(to_unsigned(6,8) ,
31143	 => std_logic_vector(to_unsigned(1,8) ,
31144	 => std_logic_vector(to_unsigned(1,8) ,
31145	 => std_logic_vector(to_unsigned(1,8) ,
31146	 => std_logic_vector(to_unsigned(11,8) ,
31147	 => std_logic_vector(to_unsigned(57,8) ,
31148	 => std_logic_vector(to_unsigned(81,8) ,
31149	 => std_logic_vector(to_unsigned(71,8) ,
31150	 => std_logic_vector(to_unsigned(41,8) ,
31151	 => std_logic_vector(to_unsigned(16,8) ,
31152	 => std_logic_vector(to_unsigned(1,8) ,
31153	 => std_logic_vector(to_unsigned(1,8) ,
31154	 => std_logic_vector(to_unsigned(1,8) ,
31155	 => std_logic_vector(to_unsigned(1,8) ,
31156	 => std_logic_vector(to_unsigned(2,8) ,
31157	 => std_logic_vector(to_unsigned(3,8) ,
31158	 => std_logic_vector(to_unsigned(2,8) ,
31159	 => std_logic_vector(to_unsigned(1,8) ,
31160	 => std_logic_vector(to_unsigned(6,8) ,
31161	 => std_logic_vector(to_unsigned(6,8) ,
31162	 => std_logic_vector(to_unsigned(2,8) ,
31163	 => std_logic_vector(to_unsigned(2,8) ,
31164	 => std_logic_vector(to_unsigned(3,8) ,
31165	 => std_logic_vector(to_unsigned(14,8) ,
31166	 => std_logic_vector(to_unsigned(46,8) ,
31167	 => std_logic_vector(to_unsigned(76,8) ,
31168	 => std_logic_vector(to_unsigned(88,8) ,
31169	 => std_logic_vector(to_unsigned(65,8) ,
31170	 => std_logic_vector(to_unsigned(44,8) ,
31171	 => std_logic_vector(to_unsigned(32,8) ,
31172	 => std_logic_vector(to_unsigned(13,8) ,
31173	 => std_logic_vector(to_unsigned(6,8) ,
31174	 => std_logic_vector(to_unsigned(10,8) ,
31175	 => std_logic_vector(to_unsigned(15,8) ,
31176	 => std_logic_vector(to_unsigned(7,8) ,
31177	 => std_logic_vector(to_unsigned(19,8) ,
31178	 => std_logic_vector(to_unsigned(15,8) ,
31179	 => std_logic_vector(to_unsigned(2,8) ,
31180	 => std_logic_vector(to_unsigned(17,8) ,
31181	 => std_logic_vector(to_unsigned(45,8) ,
31182	 => std_logic_vector(to_unsigned(64,8) ,
31183	 => std_logic_vector(to_unsigned(112,8) ,
31184	 => std_logic_vector(to_unsigned(37,8) ,
31185	 => std_logic_vector(to_unsigned(0,8) ,
31186	 => std_logic_vector(to_unsigned(0,8) ,
31187	 => std_logic_vector(to_unsigned(1,8) ,
31188	 => std_logic_vector(to_unsigned(2,8) ,
31189	 => std_logic_vector(to_unsigned(5,8) ,
31190	 => std_logic_vector(to_unsigned(25,8) ,
31191	 => std_logic_vector(to_unsigned(59,8) ,
31192	 => std_logic_vector(to_unsigned(71,8) ,
31193	 => std_logic_vector(to_unsigned(67,8) ,
31194	 => std_logic_vector(to_unsigned(73,8) ,
31195	 => std_logic_vector(to_unsigned(60,8) ,
31196	 => std_logic_vector(to_unsigned(50,8) ,
31197	 => std_logic_vector(to_unsigned(51,8) ,
31198	 => std_logic_vector(to_unsigned(43,8) ,
31199	 => std_logic_vector(to_unsigned(32,8) ,
31200	 => std_logic_vector(to_unsigned(13,8) ,
31201	 => std_logic_vector(to_unsigned(3,8) ,
31202	 => std_logic_vector(to_unsigned(1,8) ,
31203	 => std_logic_vector(to_unsigned(16,8) ,
31204	 => std_logic_vector(to_unsigned(81,8) ,
31205	 => std_logic_vector(to_unsigned(93,8) ,
31206	 => std_logic_vector(to_unsigned(108,8) ,
31207	 => std_logic_vector(to_unsigned(133,8) ,
31208	 => std_logic_vector(to_unsigned(118,8) ,
31209	 => std_logic_vector(to_unsigned(72,8) ,
31210	 => std_logic_vector(to_unsigned(90,8) ,
31211	 => std_logic_vector(to_unsigned(134,8) ,
31212	 => std_logic_vector(to_unsigned(134,8) ,
31213	 => std_logic_vector(to_unsigned(118,8) ,
31214	 => std_logic_vector(to_unsigned(130,8) ,
31215	 => std_logic_vector(to_unsigned(96,8) ,
31216	 => std_logic_vector(to_unsigned(87,8) ,
31217	 => std_logic_vector(to_unsigned(67,8) ,
31218	 => std_logic_vector(to_unsigned(51,8) ,
31219	 => std_logic_vector(to_unsigned(81,8) ,
31220	 => std_logic_vector(to_unsigned(60,8) ,
31221	 => std_logic_vector(to_unsigned(67,8) ,
31222	 => std_logic_vector(to_unsigned(86,8) ,
31223	 => std_logic_vector(to_unsigned(73,8) ,
31224	 => std_logic_vector(to_unsigned(39,8) ,
31225	 => std_logic_vector(to_unsigned(12,8) ,
31226	 => std_logic_vector(to_unsigned(27,8) ,
31227	 => std_logic_vector(to_unsigned(63,8) ,
31228	 => std_logic_vector(to_unsigned(59,8) ,
31229	 => std_logic_vector(to_unsigned(52,8) ,
31230	 => std_logic_vector(to_unsigned(65,8) ,
31231	 => std_logic_vector(to_unsigned(71,8) ,
31232	 => std_logic_vector(to_unsigned(146,8) ,
31233	 => std_logic_vector(to_unsigned(173,8) ,
31234	 => std_logic_vector(to_unsigned(164,8) ,
31235	 => std_logic_vector(to_unsigned(168,8) ,
31236	 => std_logic_vector(to_unsigned(159,8) ,
31237	 => std_logic_vector(to_unsigned(161,8) ,
31238	 => std_logic_vector(to_unsigned(144,8) ,
31239	 => std_logic_vector(to_unsigned(81,8) ,
31240	 => std_logic_vector(to_unsigned(109,8) ,
31241	 => std_logic_vector(to_unsigned(116,8) ,
31242	 => std_logic_vector(to_unsigned(96,8) ,
31243	 => std_logic_vector(to_unsigned(82,8) ,
31244	 => std_logic_vector(to_unsigned(52,8) ,
31245	 => std_logic_vector(to_unsigned(29,8) ,
31246	 => std_logic_vector(to_unsigned(8,8) ,
31247	 => std_logic_vector(to_unsigned(11,8) ,
31248	 => std_logic_vector(to_unsigned(31,8) ,
31249	 => std_logic_vector(to_unsigned(115,8) ,
31250	 => std_logic_vector(to_unsigned(166,8) ,
31251	 => std_logic_vector(to_unsigned(152,8) ,
31252	 => std_logic_vector(to_unsigned(152,8) ,
31253	 => std_logic_vector(to_unsigned(154,8) ,
31254	 => std_logic_vector(to_unsigned(156,8) ,
31255	 => std_logic_vector(to_unsigned(152,8) ,
31256	 => std_logic_vector(to_unsigned(156,8) ,
31257	 => std_logic_vector(to_unsigned(156,8) ,
31258	 => std_logic_vector(to_unsigned(152,8) ,
31259	 => std_logic_vector(to_unsigned(157,8) ,
31260	 => std_logic_vector(to_unsigned(151,8) ,
31261	 => std_logic_vector(to_unsigned(152,8) ,
31262	 => std_logic_vector(to_unsigned(152,8) ,
31263	 => std_logic_vector(to_unsigned(156,8) ,
31264	 => std_logic_vector(to_unsigned(161,8) ,
31265	 => std_logic_vector(to_unsigned(147,8) ,
31266	 => std_logic_vector(to_unsigned(142,8) ,
31267	 => std_logic_vector(to_unsigned(142,8) ,
31268	 => std_logic_vector(to_unsigned(130,8) ,
31269	 => std_logic_vector(to_unsigned(134,8) ,
31270	 => std_logic_vector(to_unsigned(138,8) ,
31271	 => std_logic_vector(to_unsigned(116,8) ,
31272	 => std_logic_vector(to_unsigned(85,8) ,
31273	 => std_logic_vector(to_unsigned(64,8) ,
31274	 => std_logic_vector(to_unsigned(36,8) ,
31275	 => std_logic_vector(to_unsigned(22,8) ,
31276	 => std_logic_vector(to_unsigned(36,8) ,
31277	 => std_logic_vector(to_unsigned(48,8) ,
31278	 => std_logic_vector(to_unsigned(27,8) ,
31279	 => std_logic_vector(to_unsigned(5,8) ,
31280	 => std_logic_vector(to_unsigned(3,8) ,
31281	 => std_logic_vector(to_unsigned(12,8) ,
31282	 => std_logic_vector(to_unsigned(10,8) ,
31283	 => std_logic_vector(to_unsigned(9,8) ,
31284	 => std_logic_vector(to_unsigned(13,8) ,
31285	 => std_logic_vector(to_unsigned(15,8) ,
31286	 => std_logic_vector(to_unsigned(7,8) ,
31287	 => std_logic_vector(to_unsigned(1,8) ,
31288	 => std_logic_vector(to_unsigned(0,8) ,
31289	 => std_logic_vector(to_unsigned(1,8) ,
31290	 => std_logic_vector(to_unsigned(0,8) ,
31291	 => std_logic_vector(to_unsigned(1,8) ,
31292	 => std_logic_vector(to_unsigned(2,8) ,
31293	 => std_logic_vector(to_unsigned(2,8) ,
31294	 => std_logic_vector(to_unsigned(3,8) ,
31295	 => std_logic_vector(to_unsigned(3,8) ,
31296	 => std_logic_vector(to_unsigned(2,8) ,
31297	 => std_logic_vector(to_unsigned(3,8) ,
31298	 => std_logic_vector(to_unsigned(7,8) ,
31299	 => std_logic_vector(to_unsigned(9,8) ,
31300	 => std_logic_vector(to_unsigned(5,8) ,
31301	 => std_logic_vector(to_unsigned(4,8) ,
31302	 => std_logic_vector(to_unsigned(5,8) ,
31303	 => std_logic_vector(to_unsigned(16,8) ,
31304	 => std_logic_vector(to_unsigned(69,8) ,
31305	 => std_logic_vector(to_unsigned(62,8) ,
31306	 => std_logic_vector(to_unsigned(38,8) ,
31307	 => std_logic_vector(to_unsigned(60,8) ,
31308	 => std_logic_vector(to_unsigned(96,8) ,
31309	 => std_logic_vector(to_unsigned(90,8) ,
31310	 => std_logic_vector(to_unsigned(76,8) ,
31311	 => std_logic_vector(to_unsigned(104,8) ,
31312	 => std_logic_vector(to_unsigned(99,8) ,
31313	 => std_logic_vector(to_unsigned(54,8) ,
31314	 => std_logic_vector(to_unsigned(7,8) ,
31315	 => std_logic_vector(to_unsigned(3,8) ,
31316	 => std_logic_vector(to_unsigned(5,8) ,
31317	 => std_logic_vector(to_unsigned(3,8) ,
31318	 => std_logic_vector(to_unsigned(3,8) ,
31319	 => std_logic_vector(to_unsigned(4,8) ,
31320	 => std_logic_vector(to_unsigned(5,8) ,
31321	 => std_logic_vector(to_unsigned(7,8) ,
31322	 => std_logic_vector(to_unsigned(5,8) ,
31323	 => std_logic_vector(to_unsigned(4,8) ,
31324	 => std_logic_vector(to_unsigned(4,8) ,
31325	 => std_logic_vector(to_unsigned(4,8) ,
31326	 => std_logic_vector(to_unsigned(6,8) ,
31327	 => std_logic_vector(to_unsigned(3,8) ,
31328	 => std_logic_vector(to_unsigned(1,8) ,
31329	 => std_logic_vector(to_unsigned(0,8) ,
31330	 => std_logic_vector(to_unsigned(3,8) ,
31331	 => std_logic_vector(to_unsigned(23,8) ,
31332	 => std_logic_vector(to_unsigned(6,8) ,
31333	 => std_logic_vector(to_unsigned(1,8) ,
31334	 => std_logic_vector(to_unsigned(17,8) ,
31335	 => std_logic_vector(to_unsigned(46,8) ,
31336	 => std_logic_vector(to_unsigned(107,8) ,
31337	 => std_logic_vector(to_unsigned(171,8) ,
31338	 => std_logic_vector(to_unsigned(156,8) ,
31339	 => std_logic_vector(to_unsigned(121,8) ,
31340	 => std_logic_vector(to_unsigned(97,8) ,
31341	 => std_logic_vector(to_unsigned(124,8) ,
31342	 => std_logic_vector(to_unsigned(147,8) ,
31343	 => std_logic_vector(to_unsigned(156,8) ,
31344	 => std_logic_vector(to_unsigned(164,8) ,
31345	 => std_logic_vector(to_unsigned(159,8) ,
31346	 => std_logic_vector(to_unsigned(161,8) ,
31347	 => std_logic_vector(to_unsigned(159,8) ,
31348	 => std_logic_vector(to_unsigned(154,8) ,
31349	 => std_logic_vector(to_unsigned(149,8) ,
31350	 => std_logic_vector(to_unsigned(144,8) ,
31351	 => std_logic_vector(to_unsigned(146,8) ,
31352	 => std_logic_vector(to_unsigned(152,8) ,
31353	 => std_logic_vector(to_unsigned(152,8) ,
31354	 => std_logic_vector(to_unsigned(151,8) ,
31355	 => std_logic_vector(to_unsigned(152,8) ,
31356	 => std_logic_vector(to_unsigned(151,8) ,
31357	 => std_logic_vector(to_unsigned(146,8) ,
31358	 => std_logic_vector(to_unsigned(142,8) ,
31359	 => std_logic_vector(to_unsigned(141,8) ,
31360	 => std_logic_vector(to_unsigned(139,8) ,
31361	 => std_logic_vector(to_unsigned(3,8) ,
31362	 => std_logic_vector(to_unsigned(3,8) ,
31363	 => std_logic_vector(to_unsigned(1,8) ,
31364	 => std_logic_vector(to_unsigned(4,8) ,
31365	 => std_logic_vector(to_unsigned(12,8) ,
31366	 => std_logic_vector(to_unsigned(10,8) ,
31367	 => std_logic_vector(to_unsigned(6,8) ,
31368	 => std_logic_vector(to_unsigned(5,8) ,
31369	 => std_logic_vector(to_unsigned(4,8) ,
31370	 => std_logic_vector(to_unsigned(1,8) ,
31371	 => std_logic_vector(to_unsigned(1,8) ,
31372	 => std_logic_vector(to_unsigned(1,8) ,
31373	 => std_logic_vector(to_unsigned(1,8) ,
31374	 => std_logic_vector(to_unsigned(0,8) ,
31375	 => std_logic_vector(to_unsigned(0,8) ,
31376	 => std_logic_vector(to_unsigned(1,8) ,
31377	 => std_logic_vector(to_unsigned(1,8) ,
31378	 => std_logic_vector(to_unsigned(2,8) ,
31379	 => std_logic_vector(to_unsigned(4,8) ,
31380	 => std_logic_vector(to_unsigned(9,8) ,
31381	 => std_logic_vector(to_unsigned(9,8) ,
31382	 => std_logic_vector(to_unsigned(6,8) ,
31383	 => std_logic_vector(to_unsigned(7,8) ,
31384	 => std_logic_vector(to_unsigned(4,8) ,
31385	 => std_logic_vector(to_unsigned(20,8) ,
31386	 => std_logic_vector(to_unsigned(47,8) ,
31387	 => std_logic_vector(to_unsigned(24,8) ,
31388	 => std_logic_vector(to_unsigned(19,8) ,
31389	 => std_logic_vector(to_unsigned(17,8) ,
31390	 => std_logic_vector(to_unsigned(7,8) ,
31391	 => std_logic_vector(to_unsigned(6,8) ,
31392	 => std_logic_vector(to_unsigned(12,8) ,
31393	 => std_logic_vector(to_unsigned(9,8) ,
31394	 => std_logic_vector(to_unsigned(9,8) ,
31395	 => std_logic_vector(to_unsigned(3,8) ,
31396	 => std_logic_vector(to_unsigned(2,8) ,
31397	 => std_logic_vector(to_unsigned(16,8) ,
31398	 => std_logic_vector(to_unsigned(56,8) ,
31399	 => std_logic_vector(to_unsigned(48,8) ,
31400	 => std_logic_vector(to_unsigned(37,8) ,
31401	 => std_logic_vector(to_unsigned(26,8) ,
31402	 => std_logic_vector(to_unsigned(14,8) ,
31403	 => std_logic_vector(to_unsigned(9,8) ,
31404	 => std_logic_vector(to_unsigned(6,8) ,
31405	 => std_logic_vector(to_unsigned(7,8) ,
31406	 => std_logic_vector(to_unsigned(4,8) ,
31407	 => std_logic_vector(to_unsigned(2,8) ,
31408	 => std_logic_vector(to_unsigned(2,8) ,
31409	 => std_logic_vector(to_unsigned(2,8) ,
31410	 => std_logic_vector(to_unsigned(1,8) ,
31411	 => std_logic_vector(to_unsigned(4,8) ,
31412	 => std_logic_vector(to_unsigned(9,8) ,
31413	 => std_logic_vector(to_unsigned(22,8) ,
31414	 => std_logic_vector(to_unsigned(46,8) ,
31415	 => std_logic_vector(to_unsigned(55,8) ,
31416	 => std_logic_vector(to_unsigned(47,8) ,
31417	 => std_logic_vector(to_unsigned(40,8) ,
31418	 => std_logic_vector(to_unsigned(35,8) ,
31419	 => std_logic_vector(to_unsigned(17,8) ,
31420	 => std_logic_vector(to_unsigned(2,8) ,
31421	 => std_logic_vector(to_unsigned(3,8) ,
31422	 => std_logic_vector(to_unsigned(18,8) ,
31423	 => std_logic_vector(to_unsigned(4,8) ,
31424	 => std_logic_vector(to_unsigned(6,8) ,
31425	 => std_logic_vector(to_unsigned(91,8) ,
31426	 => std_logic_vector(to_unsigned(99,8) ,
31427	 => std_logic_vector(to_unsigned(51,8) ,
31428	 => std_logic_vector(to_unsigned(17,8) ,
31429	 => std_logic_vector(to_unsigned(4,8) ,
31430	 => std_logic_vector(to_unsigned(1,8) ,
31431	 => std_logic_vector(to_unsigned(3,8) ,
31432	 => std_logic_vector(to_unsigned(4,8) ,
31433	 => std_logic_vector(to_unsigned(6,8) ,
31434	 => std_logic_vector(to_unsigned(16,8) ,
31435	 => std_logic_vector(to_unsigned(24,8) ,
31436	 => std_logic_vector(to_unsigned(29,8) ,
31437	 => std_logic_vector(to_unsigned(18,8) ,
31438	 => std_logic_vector(to_unsigned(10,8) ,
31439	 => std_logic_vector(to_unsigned(5,8) ,
31440	 => std_logic_vector(to_unsigned(55,8) ,
31441	 => std_logic_vector(to_unsigned(157,8) ,
31442	 => std_logic_vector(to_unsigned(128,8) ,
31443	 => std_logic_vector(to_unsigned(154,8) ,
31444	 => std_logic_vector(to_unsigned(156,8) ,
31445	 => std_logic_vector(to_unsigned(152,8) ,
31446	 => std_logic_vector(to_unsigned(134,8) ,
31447	 => std_logic_vector(to_unsigned(131,8) ,
31448	 => std_logic_vector(to_unsigned(80,8) ,
31449	 => std_logic_vector(to_unsigned(17,8) ,
31450	 => std_logic_vector(to_unsigned(15,8) ,
31451	 => std_logic_vector(to_unsigned(22,8) ,
31452	 => std_logic_vector(to_unsigned(33,8) ,
31453	 => std_logic_vector(to_unsigned(35,8) ,
31454	 => std_logic_vector(to_unsigned(6,8) ,
31455	 => std_logic_vector(to_unsigned(2,8) ,
31456	 => std_logic_vector(to_unsigned(2,8) ,
31457	 => std_logic_vector(to_unsigned(8,8) ,
31458	 => std_logic_vector(to_unsigned(8,8) ,
31459	 => std_logic_vector(to_unsigned(3,8) ,
31460	 => std_logic_vector(to_unsigned(6,8) ,
31461	 => std_logic_vector(to_unsigned(5,8) ,
31462	 => std_logic_vector(to_unsigned(4,8) ,
31463	 => std_logic_vector(to_unsigned(2,8) ,
31464	 => std_logic_vector(to_unsigned(3,8) ,
31465	 => std_logic_vector(to_unsigned(8,8) ,
31466	 => std_logic_vector(to_unsigned(8,8) ,
31467	 => std_logic_vector(to_unsigned(51,8) ,
31468	 => std_logic_vector(to_unsigned(92,8) ,
31469	 => std_logic_vector(to_unsigned(77,8) ,
31470	 => std_logic_vector(to_unsigned(42,8) ,
31471	 => std_logic_vector(to_unsigned(13,8) ,
31472	 => std_logic_vector(to_unsigned(2,8) ,
31473	 => std_logic_vector(to_unsigned(2,8) ,
31474	 => std_logic_vector(to_unsigned(2,8) ,
31475	 => std_logic_vector(to_unsigned(0,8) ,
31476	 => std_logic_vector(to_unsigned(0,8) ,
31477	 => std_logic_vector(to_unsigned(2,8) ,
31478	 => std_logic_vector(to_unsigned(3,8) ,
31479	 => std_logic_vector(to_unsigned(2,8) ,
31480	 => std_logic_vector(to_unsigned(4,8) ,
31481	 => std_logic_vector(to_unsigned(4,8) ,
31482	 => std_logic_vector(to_unsigned(4,8) ,
31483	 => std_logic_vector(to_unsigned(15,8) ,
31484	 => std_logic_vector(to_unsigned(46,8) ,
31485	 => std_logic_vector(to_unsigned(82,8) ,
31486	 => std_logic_vector(to_unsigned(96,8) ,
31487	 => std_logic_vector(to_unsigned(105,8) ,
31488	 => std_logic_vector(to_unsigned(82,8) ,
31489	 => std_logic_vector(to_unsigned(30,8) ,
31490	 => std_logic_vector(to_unsigned(14,8) ,
31491	 => std_logic_vector(to_unsigned(11,8) ,
31492	 => std_logic_vector(to_unsigned(13,8) ,
31493	 => std_logic_vector(to_unsigned(8,8) ,
31494	 => std_logic_vector(to_unsigned(5,8) ,
31495	 => std_logic_vector(to_unsigned(12,8) ,
31496	 => std_logic_vector(to_unsigned(6,8) ,
31497	 => std_logic_vector(to_unsigned(11,8) ,
31498	 => std_logic_vector(to_unsigned(5,8) ,
31499	 => std_logic_vector(to_unsigned(1,8) ,
31500	 => std_logic_vector(to_unsigned(2,8) ,
31501	 => std_logic_vector(to_unsigned(2,8) ,
31502	 => std_logic_vector(to_unsigned(2,8) ,
31503	 => std_logic_vector(to_unsigned(4,8) ,
31504	 => std_logic_vector(to_unsigned(10,8) ,
31505	 => std_logic_vector(to_unsigned(8,8) ,
31506	 => std_logic_vector(to_unsigned(7,8) ,
31507	 => std_logic_vector(to_unsigned(12,8) ,
31508	 => std_logic_vector(to_unsigned(12,8) ,
31509	 => std_logic_vector(to_unsigned(14,8) ,
31510	 => std_logic_vector(to_unsigned(25,8) ,
31511	 => std_logic_vector(to_unsigned(23,8) ,
31512	 => std_logic_vector(to_unsigned(52,8) ,
31513	 => std_logic_vector(to_unsigned(64,8) ,
31514	 => std_logic_vector(to_unsigned(51,8) ,
31515	 => std_logic_vector(to_unsigned(48,8) ,
31516	 => std_logic_vector(to_unsigned(38,8) ,
31517	 => std_logic_vector(to_unsigned(26,8) ,
31518	 => std_logic_vector(to_unsigned(13,8) ,
31519	 => std_logic_vector(to_unsigned(10,8) ,
31520	 => std_logic_vector(to_unsigned(6,8) ,
31521	 => std_logic_vector(to_unsigned(1,8) ,
31522	 => std_logic_vector(to_unsigned(0,8) ,
31523	 => std_logic_vector(to_unsigned(2,8) ,
31524	 => std_logic_vector(to_unsigned(39,8) ,
31525	 => std_logic_vector(to_unsigned(100,8) ,
31526	 => std_logic_vector(to_unsigned(116,8) ,
31527	 => std_logic_vector(to_unsigned(104,8) ,
31528	 => std_logic_vector(to_unsigned(67,8) ,
31529	 => std_logic_vector(to_unsigned(78,8) ,
31530	 => std_logic_vector(to_unsigned(81,8) ,
31531	 => std_logic_vector(to_unsigned(80,8) ,
31532	 => std_logic_vector(to_unsigned(127,8) ,
31533	 => std_logic_vector(to_unsigned(103,8) ,
31534	 => std_logic_vector(to_unsigned(64,8) ,
31535	 => std_logic_vector(to_unsigned(52,8) ,
31536	 => std_logic_vector(to_unsigned(43,8) ,
31537	 => std_logic_vector(to_unsigned(29,8) ,
31538	 => std_logic_vector(to_unsigned(41,8) ,
31539	 => std_logic_vector(to_unsigned(96,8) ,
31540	 => std_logic_vector(to_unsigned(79,8) ,
31541	 => std_logic_vector(to_unsigned(54,8) ,
31542	 => std_logic_vector(to_unsigned(51,8) ,
31543	 => std_logic_vector(to_unsigned(40,8) ,
31544	 => std_logic_vector(to_unsigned(15,8) ,
31545	 => std_logic_vector(to_unsigned(2,8) ,
31546	 => std_logic_vector(to_unsigned(14,8) ,
31547	 => std_logic_vector(to_unsigned(54,8) ,
31548	 => std_logic_vector(to_unsigned(66,8) ,
31549	 => std_logic_vector(to_unsigned(61,8) ,
31550	 => std_logic_vector(to_unsigned(32,8) ,
31551	 => std_logic_vector(to_unsigned(35,8) ,
31552	 => std_logic_vector(to_unsigned(54,8) ,
31553	 => std_logic_vector(to_unsigned(90,8) ,
31554	 => std_logic_vector(to_unsigned(163,8) ,
31555	 => std_logic_vector(to_unsigned(156,8) ,
31556	 => std_logic_vector(to_unsigned(151,8) ,
31557	 => std_logic_vector(to_unsigned(164,8) ,
31558	 => std_logic_vector(to_unsigned(138,8) ,
31559	 => std_logic_vector(to_unsigned(51,8) ,
31560	 => std_logic_vector(to_unsigned(99,8) ,
31561	 => std_logic_vector(to_unsigned(118,8) ,
31562	 => std_logic_vector(to_unsigned(108,8) ,
31563	 => std_logic_vector(to_unsigned(96,8) ,
31564	 => std_logic_vector(to_unsigned(51,8) ,
31565	 => std_logic_vector(to_unsigned(20,8) ,
31566	 => std_logic_vector(to_unsigned(25,8) ,
31567	 => std_logic_vector(to_unsigned(72,8) ,
31568	 => std_logic_vector(to_unsigned(73,8) ,
31569	 => std_logic_vector(to_unsigned(92,8) ,
31570	 => std_logic_vector(to_unsigned(159,8) ,
31571	 => std_logic_vector(to_unsigned(156,8) ,
31572	 => std_logic_vector(to_unsigned(156,8) ,
31573	 => std_logic_vector(to_unsigned(154,8) ,
31574	 => std_logic_vector(to_unsigned(157,8) ,
31575	 => std_logic_vector(to_unsigned(152,8) ,
31576	 => std_logic_vector(to_unsigned(152,8) ,
31577	 => std_logic_vector(to_unsigned(156,8) ,
31578	 => std_logic_vector(to_unsigned(152,8) ,
31579	 => std_logic_vector(to_unsigned(156,8) ,
31580	 => std_logic_vector(to_unsigned(154,8) ,
31581	 => std_logic_vector(to_unsigned(144,8) ,
31582	 => std_logic_vector(to_unsigned(142,8) ,
31583	 => std_logic_vector(to_unsigned(141,8) ,
31584	 => std_logic_vector(to_unsigned(146,8) ,
31585	 => std_logic_vector(to_unsigned(163,8) ,
31586	 => std_logic_vector(to_unsigned(164,8) ,
31587	 => std_logic_vector(to_unsigned(154,8) ,
31588	 => std_logic_vector(to_unsigned(159,8) ,
31589	 => std_logic_vector(to_unsigned(127,8) ,
31590	 => std_logic_vector(to_unsigned(122,8) ,
31591	 => std_logic_vector(to_unsigned(130,8) ,
31592	 => std_logic_vector(to_unsigned(101,8) ,
31593	 => std_logic_vector(to_unsigned(82,8) ,
31594	 => std_logic_vector(to_unsigned(45,8) ,
31595	 => std_logic_vector(to_unsigned(17,8) ,
31596	 => std_logic_vector(to_unsigned(35,8) ,
31597	 => std_logic_vector(to_unsigned(39,8) ,
31598	 => std_logic_vector(to_unsigned(17,8) ,
31599	 => std_logic_vector(to_unsigned(4,8) ,
31600	 => std_logic_vector(to_unsigned(18,8) ,
31601	 => std_logic_vector(to_unsigned(51,8) ,
31602	 => std_logic_vector(to_unsigned(40,8) ,
31603	 => std_logic_vector(to_unsigned(30,8) ,
31604	 => std_logic_vector(to_unsigned(19,8) ,
31605	 => std_logic_vector(to_unsigned(8,8) ,
31606	 => std_logic_vector(to_unsigned(5,8) ,
31607	 => std_logic_vector(to_unsigned(2,8) ,
31608	 => std_logic_vector(to_unsigned(1,8) ,
31609	 => std_logic_vector(to_unsigned(2,8) ,
31610	 => std_logic_vector(to_unsigned(3,8) ,
31611	 => std_logic_vector(to_unsigned(3,8) ,
31612	 => std_logic_vector(to_unsigned(2,8) ,
31613	 => std_logic_vector(to_unsigned(2,8) ,
31614	 => std_logic_vector(to_unsigned(2,8) ,
31615	 => std_logic_vector(to_unsigned(0,8) ,
31616	 => std_logic_vector(to_unsigned(1,8) ,
31617	 => std_logic_vector(to_unsigned(2,8) ,
31618	 => std_logic_vector(to_unsigned(5,8) ,
31619	 => std_logic_vector(to_unsigned(14,8) ,
31620	 => std_logic_vector(to_unsigned(6,8) ,
31621	 => std_logic_vector(to_unsigned(6,8) ,
31622	 => std_logic_vector(to_unsigned(8,8) ,
31623	 => std_logic_vector(to_unsigned(19,8) ,
31624	 => std_logic_vector(to_unsigned(70,8) ,
31625	 => std_logic_vector(to_unsigned(82,8) ,
31626	 => std_logic_vector(to_unsigned(55,8) ,
31627	 => std_logic_vector(to_unsigned(29,8) ,
31628	 => std_logic_vector(to_unsigned(23,8) ,
31629	 => std_logic_vector(to_unsigned(45,8) ,
31630	 => std_logic_vector(to_unsigned(58,8) ,
31631	 => std_logic_vector(to_unsigned(59,8) ,
31632	 => std_logic_vector(to_unsigned(105,8) ,
31633	 => std_logic_vector(to_unsigned(63,8) ,
31634	 => std_logic_vector(to_unsigned(4,8) ,
31635	 => std_logic_vector(to_unsigned(4,8) ,
31636	 => std_logic_vector(to_unsigned(4,8) ,
31637	 => std_logic_vector(to_unsigned(3,8) ,
31638	 => std_logic_vector(to_unsigned(6,8) ,
31639	 => std_logic_vector(to_unsigned(9,8) ,
31640	 => std_logic_vector(to_unsigned(6,8) ,
31641	 => std_logic_vector(to_unsigned(6,8) ,
31642	 => std_logic_vector(to_unsigned(5,8) ,
31643	 => std_logic_vector(to_unsigned(5,8) ,
31644	 => std_logic_vector(to_unsigned(4,8) ,
31645	 => std_logic_vector(to_unsigned(3,8) ,
31646	 => std_logic_vector(to_unsigned(4,8) ,
31647	 => std_logic_vector(to_unsigned(4,8) ,
31648	 => std_logic_vector(to_unsigned(2,8) ,
31649	 => std_logic_vector(to_unsigned(0,8) ,
31650	 => std_logic_vector(to_unsigned(0,8) ,
31651	 => std_logic_vector(to_unsigned(10,8) ,
31652	 => std_logic_vector(to_unsigned(8,8) ,
31653	 => std_logic_vector(to_unsigned(1,8) ,
31654	 => std_logic_vector(to_unsigned(3,8) ,
31655	 => std_logic_vector(to_unsigned(9,8) ,
31656	 => std_logic_vector(to_unsigned(20,8) ,
31657	 => std_logic_vector(to_unsigned(51,8) ,
31658	 => std_logic_vector(to_unsigned(84,8) ,
31659	 => std_logic_vector(to_unsigned(90,8) ,
31660	 => std_logic_vector(to_unsigned(69,8) ,
31661	 => std_logic_vector(to_unsigned(115,8) ,
31662	 => std_logic_vector(to_unsigned(152,8) ,
31663	 => std_logic_vector(to_unsigned(146,8) ,
31664	 => std_logic_vector(to_unsigned(159,8) ,
31665	 => std_logic_vector(to_unsigned(154,8) ,
31666	 => std_logic_vector(to_unsigned(157,8) ,
31667	 => std_logic_vector(to_unsigned(157,8) ,
31668	 => std_logic_vector(to_unsigned(152,8) ,
31669	 => std_logic_vector(to_unsigned(141,8) ,
31670	 => std_logic_vector(to_unsigned(136,8) ,
31671	 => std_logic_vector(to_unsigned(138,8) ,
31672	 => std_logic_vector(to_unsigned(139,8) ,
31673	 => std_logic_vector(to_unsigned(141,8) ,
31674	 => std_logic_vector(to_unsigned(141,8) ,
31675	 => std_logic_vector(to_unsigned(146,8) ,
31676	 => std_logic_vector(to_unsigned(144,8) ,
31677	 => std_logic_vector(to_unsigned(138,8) ,
31678	 => std_logic_vector(to_unsigned(133,8) ,
31679	 => std_logic_vector(to_unsigned(130,8) ,
31680	 => std_logic_vector(to_unsigned(130,8) ,
31681	 => std_logic_vector(to_unsigned(3,8) ,
31682	 => std_logic_vector(to_unsigned(3,8) ,
31683	 => std_logic_vector(to_unsigned(2,8) ,
31684	 => std_logic_vector(to_unsigned(6,8) ,
31685	 => std_logic_vector(to_unsigned(7,8) ,
31686	 => std_logic_vector(to_unsigned(7,8) ,
31687	 => std_logic_vector(to_unsigned(6,8) ,
31688	 => std_logic_vector(to_unsigned(5,8) ,
31689	 => std_logic_vector(to_unsigned(3,8) ,
31690	 => std_logic_vector(to_unsigned(2,8) ,
31691	 => std_logic_vector(to_unsigned(0,8) ,
31692	 => std_logic_vector(to_unsigned(1,8) ,
31693	 => std_logic_vector(to_unsigned(1,8) ,
31694	 => std_logic_vector(to_unsigned(1,8) ,
31695	 => std_logic_vector(to_unsigned(1,8) ,
31696	 => std_logic_vector(to_unsigned(1,8) ,
31697	 => std_logic_vector(to_unsigned(1,8) ,
31698	 => std_logic_vector(to_unsigned(1,8) ,
31699	 => std_logic_vector(to_unsigned(1,8) ,
31700	 => std_logic_vector(to_unsigned(3,8) ,
31701	 => std_logic_vector(to_unsigned(7,8) ,
31702	 => std_logic_vector(to_unsigned(10,8) ,
31703	 => std_logic_vector(to_unsigned(7,8) ,
31704	 => std_logic_vector(to_unsigned(2,8) ,
31705	 => std_logic_vector(to_unsigned(16,8) ,
31706	 => std_logic_vector(to_unsigned(30,8) ,
31707	 => std_logic_vector(to_unsigned(19,8) ,
31708	 => std_logic_vector(to_unsigned(17,8) ,
31709	 => std_logic_vector(to_unsigned(8,8) ,
31710	 => std_logic_vector(to_unsigned(4,8) ,
31711	 => std_logic_vector(to_unsigned(3,8) ,
31712	 => std_logic_vector(to_unsigned(1,8) ,
31713	 => std_logic_vector(to_unsigned(1,8) ,
31714	 => std_logic_vector(to_unsigned(1,8) ,
31715	 => std_logic_vector(to_unsigned(1,8) ,
31716	 => std_logic_vector(to_unsigned(2,8) ,
31717	 => std_logic_vector(to_unsigned(28,8) ,
31718	 => std_logic_vector(to_unsigned(46,8) ,
31719	 => std_logic_vector(to_unsigned(35,8) ,
31720	 => std_logic_vector(to_unsigned(24,8) ,
31721	 => std_logic_vector(to_unsigned(13,8) ,
31722	 => std_logic_vector(to_unsigned(17,8) ,
31723	 => std_logic_vector(to_unsigned(14,8) ,
31724	 => std_logic_vector(to_unsigned(9,8) ,
31725	 => std_logic_vector(to_unsigned(8,8) ,
31726	 => std_logic_vector(to_unsigned(3,8) ,
31727	 => std_logic_vector(to_unsigned(1,8) ,
31728	 => std_logic_vector(to_unsigned(1,8) ,
31729	 => std_logic_vector(to_unsigned(0,8) ,
31730	 => std_logic_vector(to_unsigned(3,8) ,
31731	 => std_logic_vector(to_unsigned(24,8) ,
31732	 => std_logic_vector(to_unsigned(44,8) ,
31733	 => std_logic_vector(to_unsigned(55,8) ,
31734	 => std_logic_vector(to_unsigned(59,8) ,
31735	 => std_logic_vector(to_unsigned(44,8) ,
31736	 => std_logic_vector(to_unsigned(52,8) ,
31737	 => std_logic_vector(to_unsigned(49,8) ,
31738	 => std_logic_vector(to_unsigned(36,8) ,
31739	 => std_logic_vector(to_unsigned(19,8) ,
31740	 => std_logic_vector(to_unsigned(9,8) ,
31741	 => std_logic_vector(to_unsigned(4,8) ,
31742	 => std_logic_vector(to_unsigned(1,8) ,
31743	 => std_logic_vector(to_unsigned(0,8) ,
31744	 => std_logic_vector(to_unsigned(1,8) ,
31745	 => std_logic_vector(to_unsigned(49,8) ,
31746	 => std_logic_vector(to_unsigned(146,8) ,
31747	 => std_logic_vector(to_unsigned(27,8) ,
31748	 => std_logic_vector(to_unsigned(5,8) ,
31749	 => std_logic_vector(to_unsigned(12,8) ,
31750	 => std_logic_vector(to_unsigned(8,8) ,
31751	 => std_logic_vector(to_unsigned(5,8) ,
31752	 => std_logic_vector(to_unsigned(2,8) ,
31753	 => std_logic_vector(to_unsigned(4,8) ,
31754	 => std_logic_vector(to_unsigned(14,8) ,
31755	 => std_logic_vector(to_unsigned(20,8) ,
31756	 => std_logic_vector(to_unsigned(19,8) ,
31757	 => std_logic_vector(to_unsigned(16,8) ,
31758	 => std_logic_vector(to_unsigned(12,8) ,
31759	 => std_logic_vector(to_unsigned(4,8) ,
31760	 => std_logic_vector(to_unsigned(73,8) ,
31761	 => std_logic_vector(to_unsigned(154,8) ,
31762	 => std_logic_vector(to_unsigned(86,8) ,
31763	 => std_logic_vector(to_unsigned(104,8) ,
31764	 => std_logic_vector(to_unsigned(99,8) ,
31765	 => std_logic_vector(to_unsigned(84,8) ,
31766	 => std_logic_vector(to_unsigned(81,8) ,
31767	 => std_logic_vector(to_unsigned(114,8) ,
31768	 => std_logic_vector(to_unsigned(26,8) ,
31769	 => std_logic_vector(to_unsigned(0,8) ,
31770	 => std_logic_vector(to_unsigned(1,8) ,
31771	 => std_logic_vector(to_unsigned(2,8) ,
31772	 => std_logic_vector(to_unsigned(5,8) ,
31773	 => std_logic_vector(to_unsigned(3,8) ,
31774	 => std_logic_vector(to_unsigned(1,8) ,
31775	 => std_logic_vector(to_unsigned(2,8) ,
31776	 => std_logic_vector(to_unsigned(1,8) ,
31777	 => std_logic_vector(to_unsigned(2,8) ,
31778	 => std_logic_vector(to_unsigned(2,8) ,
31779	 => std_logic_vector(to_unsigned(3,8) ,
31780	 => std_logic_vector(to_unsigned(3,8) ,
31781	 => std_logic_vector(to_unsigned(1,8) ,
31782	 => std_logic_vector(to_unsigned(1,8) ,
31783	 => std_logic_vector(to_unsigned(6,8) ,
31784	 => std_logic_vector(to_unsigned(17,8) ,
31785	 => std_logic_vector(to_unsigned(13,8) ,
31786	 => std_logic_vector(to_unsigned(5,8) ,
31787	 => std_logic_vector(to_unsigned(42,8) ,
31788	 => std_logic_vector(to_unsigned(100,8) ,
31789	 => std_logic_vector(to_unsigned(84,8) ,
31790	 => std_logic_vector(to_unsigned(39,8) ,
31791	 => std_logic_vector(to_unsigned(7,8) ,
31792	 => std_logic_vector(to_unsigned(2,8) ,
31793	 => std_logic_vector(to_unsigned(3,8) ,
31794	 => std_logic_vector(to_unsigned(2,8) ,
31795	 => std_logic_vector(to_unsigned(1,8) ,
31796	 => std_logic_vector(to_unsigned(1,8) ,
31797	 => std_logic_vector(to_unsigned(2,8) ,
31798	 => std_logic_vector(to_unsigned(6,8) ,
31799	 => std_logic_vector(to_unsigned(9,8) ,
31800	 => std_logic_vector(to_unsigned(27,8) ,
31801	 => std_logic_vector(to_unsigned(41,8) ,
31802	 => std_logic_vector(to_unsigned(45,8) ,
31803	 => std_logic_vector(to_unsigned(90,8) ,
31804	 => std_logic_vector(to_unsigned(108,8) ,
31805	 => std_logic_vector(to_unsigned(105,8) ,
31806	 => std_logic_vector(to_unsigned(84,8) ,
31807	 => std_logic_vector(to_unsigned(46,8) ,
31808	 => std_logic_vector(to_unsigned(21,8) ,
31809	 => std_logic_vector(to_unsigned(5,8) ,
31810	 => std_logic_vector(to_unsigned(6,8) ,
31811	 => std_logic_vector(to_unsigned(12,8) ,
31812	 => std_logic_vector(to_unsigned(14,8) ,
31813	 => std_logic_vector(to_unsigned(12,8) ,
31814	 => std_logic_vector(to_unsigned(6,8) ,
31815	 => std_logic_vector(to_unsigned(7,8) ,
31816	 => std_logic_vector(to_unsigned(3,8) ,
31817	 => std_logic_vector(to_unsigned(3,8) ,
31818	 => std_logic_vector(to_unsigned(3,8) ,
31819	 => std_logic_vector(to_unsigned(4,8) ,
31820	 => std_logic_vector(to_unsigned(5,8) ,
31821	 => std_logic_vector(to_unsigned(4,8) ,
31822	 => std_logic_vector(to_unsigned(3,8) ,
31823	 => std_logic_vector(to_unsigned(1,8) ,
31824	 => std_logic_vector(to_unsigned(5,8) ,
31825	 => std_logic_vector(to_unsigned(21,8) ,
31826	 => std_logic_vector(to_unsigned(18,8) ,
31827	 => std_logic_vector(to_unsigned(11,8) ,
31828	 => std_logic_vector(to_unsigned(15,8) ,
31829	 => std_logic_vector(to_unsigned(20,8) ,
31830	 => std_logic_vector(to_unsigned(13,8) ,
31831	 => std_logic_vector(to_unsigned(12,8) ,
31832	 => std_logic_vector(to_unsigned(16,8) ,
31833	 => std_logic_vector(to_unsigned(27,8) ,
31834	 => std_logic_vector(to_unsigned(25,8) ,
31835	 => std_logic_vector(to_unsigned(22,8) ,
31836	 => std_logic_vector(to_unsigned(22,8) ,
31837	 => std_logic_vector(to_unsigned(12,8) ,
31838	 => std_logic_vector(to_unsigned(5,8) ,
31839	 => std_logic_vector(to_unsigned(3,8) ,
31840	 => std_logic_vector(to_unsigned(2,8) ,
31841	 => std_logic_vector(to_unsigned(1,8) ,
31842	 => std_logic_vector(to_unsigned(6,8) ,
31843	 => std_logic_vector(to_unsigned(9,8) ,
31844	 => std_logic_vector(to_unsigned(7,8) ,
31845	 => std_logic_vector(to_unsigned(41,8) ,
31846	 => std_logic_vector(to_unsigned(85,8) ,
31847	 => std_logic_vector(to_unsigned(80,8) ,
31848	 => std_logic_vector(to_unsigned(69,8) ,
31849	 => std_logic_vector(to_unsigned(45,8) ,
31850	 => std_logic_vector(to_unsigned(11,8) ,
31851	 => std_logic_vector(to_unsigned(16,8) ,
31852	 => std_logic_vector(to_unsigned(39,8) ,
31853	 => std_logic_vector(to_unsigned(17,8) ,
31854	 => std_logic_vector(to_unsigned(35,8) ,
31855	 => std_logic_vector(to_unsigned(66,8) ,
31856	 => std_logic_vector(to_unsigned(64,8) ,
31857	 => std_logic_vector(to_unsigned(77,8) ,
31858	 => std_logic_vector(to_unsigned(91,8) ,
31859	 => std_logic_vector(to_unsigned(100,8) ,
31860	 => std_logic_vector(to_unsigned(44,8) ,
31861	 => std_logic_vector(to_unsigned(45,8) ,
31862	 => std_logic_vector(to_unsigned(62,8) ,
31863	 => std_logic_vector(to_unsigned(17,8) ,
31864	 => std_logic_vector(to_unsigned(1,8) ,
31865	 => std_logic_vector(to_unsigned(1,8) ,
31866	 => std_logic_vector(to_unsigned(18,8) ,
31867	 => std_logic_vector(to_unsigned(54,8) ,
31868	 => std_logic_vector(to_unsigned(76,8) ,
31869	 => std_logic_vector(to_unsigned(62,8) ,
31870	 => std_logic_vector(to_unsigned(41,8) ,
31871	 => std_logic_vector(to_unsigned(14,8) ,
31872	 => std_logic_vector(to_unsigned(0,8) ,
31873	 => std_logic_vector(to_unsigned(7,8) ,
31874	 => std_logic_vector(to_unsigned(125,8) ,
31875	 => std_logic_vector(to_unsigned(168,8) ,
31876	 => std_logic_vector(to_unsigned(146,8) ,
31877	 => std_logic_vector(to_unsigned(161,8) ,
31878	 => std_logic_vector(to_unsigned(151,8) ,
31879	 => std_logic_vector(to_unsigned(88,8) ,
31880	 => std_logic_vector(to_unsigned(92,8) ,
31881	 => std_logic_vector(to_unsigned(127,8) ,
31882	 => std_logic_vector(to_unsigned(72,8) ,
31883	 => std_logic_vector(to_unsigned(29,8) ,
31884	 => std_logic_vector(to_unsigned(25,8) ,
31885	 => std_logic_vector(to_unsigned(51,8) ,
31886	 => std_logic_vector(to_unsigned(90,8) ,
31887	 => std_logic_vector(to_unsigned(91,8) ,
31888	 => std_logic_vector(to_unsigned(72,8) ,
31889	 => std_logic_vector(to_unsigned(125,8) ,
31890	 => std_logic_vector(to_unsigned(164,8) ,
31891	 => std_logic_vector(to_unsigned(152,8) ,
31892	 => std_logic_vector(to_unsigned(154,8) ,
31893	 => std_logic_vector(to_unsigned(157,8) ,
31894	 => std_logic_vector(to_unsigned(156,8) ,
31895	 => std_logic_vector(to_unsigned(157,8) ,
31896	 => std_logic_vector(to_unsigned(154,8) ,
31897	 => std_logic_vector(to_unsigned(156,8) ,
31898	 => std_logic_vector(to_unsigned(157,8) ,
31899	 => std_logic_vector(to_unsigned(156,8) ,
31900	 => std_logic_vector(to_unsigned(154,8) ,
31901	 => std_logic_vector(to_unsigned(154,8) ,
31902	 => std_logic_vector(to_unsigned(139,8) ,
31903	 => std_logic_vector(to_unsigned(134,8) ,
31904	 => std_logic_vector(to_unsigned(136,8) ,
31905	 => std_logic_vector(to_unsigned(119,8) ,
31906	 => std_logic_vector(to_unsigned(33,8) ,
31907	 => std_logic_vector(to_unsigned(12,8) ,
31908	 => std_logic_vector(to_unsigned(63,8) ,
31909	 => std_logic_vector(to_unsigned(37,8) ,
31910	 => std_logic_vector(to_unsigned(17,8) ,
31911	 => std_logic_vector(to_unsigned(104,8) ,
31912	 => std_logic_vector(to_unsigned(122,8) ,
31913	 => std_logic_vector(to_unsigned(88,8) ,
31914	 => std_logic_vector(to_unsigned(51,8) ,
31915	 => std_logic_vector(to_unsigned(13,8) ,
31916	 => std_logic_vector(to_unsigned(23,8) ,
31917	 => std_logic_vector(to_unsigned(32,8) ,
31918	 => std_logic_vector(to_unsigned(8,8) ,
31919	 => std_logic_vector(to_unsigned(27,8) ,
31920	 => std_logic_vector(to_unsigned(154,8) ,
31921	 => std_logic_vector(to_unsigned(154,8) ,
31922	 => std_logic_vector(to_unsigned(144,8) ,
31923	 => std_logic_vector(to_unsigned(166,8) ,
31924	 => std_logic_vector(to_unsigned(86,8) ,
31925	 => std_logic_vector(to_unsigned(4,8) ,
31926	 => std_logic_vector(to_unsigned(6,8) ,
31927	 => std_logic_vector(to_unsigned(60,8) ,
31928	 => std_logic_vector(to_unsigned(91,8) ,
31929	 => std_logic_vector(to_unsigned(97,8) ,
31930	 => std_logic_vector(to_unsigned(112,8) ,
31931	 => std_logic_vector(to_unsigned(109,8) ,
31932	 => std_logic_vector(to_unsigned(91,8) ,
31933	 => std_logic_vector(to_unsigned(80,8) ,
31934	 => std_logic_vector(to_unsigned(74,8) ,
31935	 => std_logic_vector(to_unsigned(30,8) ,
31936	 => std_logic_vector(to_unsigned(2,8) ,
31937	 => std_logic_vector(to_unsigned(2,8) ,
31938	 => std_logic_vector(to_unsigned(4,8) ,
31939	 => std_logic_vector(to_unsigned(15,8) ,
31940	 => std_logic_vector(to_unsigned(13,8) ,
31941	 => std_logic_vector(to_unsigned(6,8) ,
31942	 => std_logic_vector(to_unsigned(9,8) ,
31943	 => std_logic_vector(to_unsigned(17,8) ,
31944	 => std_logic_vector(to_unsigned(42,8) ,
31945	 => std_logic_vector(to_unsigned(47,8) ,
31946	 => std_logic_vector(to_unsigned(45,8) ,
31947	 => std_logic_vector(to_unsigned(47,8) ,
31948	 => std_logic_vector(to_unsigned(9,8) ,
31949	 => std_logic_vector(to_unsigned(2,8) ,
31950	 => std_logic_vector(to_unsigned(49,8) ,
31951	 => std_logic_vector(to_unsigned(107,8) ,
31952	 => std_logic_vector(to_unsigned(49,8) ,
31953	 => std_logic_vector(to_unsigned(6,8) ,
31954	 => std_logic_vector(to_unsigned(0,8) ,
31955	 => std_logic_vector(to_unsigned(4,8) ,
31956	 => std_logic_vector(to_unsigned(10,8) ,
31957	 => std_logic_vector(to_unsigned(8,8) ,
31958	 => std_logic_vector(to_unsigned(10,8) ,
31959	 => std_logic_vector(to_unsigned(6,8) ,
31960	 => std_logic_vector(to_unsigned(5,8) ,
31961	 => std_logic_vector(to_unsigned(5,8) ,
31962	 => std_logic_vector(to_unsigned(6,8) ,
31963	 => std_logic_vector(to_unsigned(5,8) ,
31964	 => std_logic_vector(to_unsigned(5,8) ,
31965	 => std_logic_vector(to_unsigned(3,8) ,
31966	 => std_logic_vector(to_unsigned(4,8) ,
31967	 => std_logic_vector(to_unsigned(7,8) ,
31968	 => std_logic_vector(to_unsigned(5,8) ,
31969	 => std_logic_vector(to_unsigned(3,8) ,
31970	 => std_logic_vector(to_unsigned(1,8) ,
31971	 => std_logic_vector(to_unsigned(1,8) ,
31972	 => std_logic_vector(to_unsigned(4,8) ,
31973	 => std_logic_vector(to_unsigned(2,8) ,
31974	 => std_logic_vector(to_unsigned(1,8) ,
31975	 => std_logic_vector(to_unsigned(2,8) ,
31976	 => std_logic_vector(to_unsigned(7,8) ,
31977	 => std_logic_vector(to_unsigned(23,8) ,
31978	 => std_logic_vector(to_unsigned(101,8) ,
31979	 => std_logic_vector(to_unsigned(168,8) ,
31980	 => std_logic_vector(to_unsigned(152,8) ,
31981	 => std_logic_vector(to_unsigned(159,8) ,
31982	 => std_logic_vector(to_unsigned(154,8) ,
31983	 => std_logic_vector(to_unsigned(156,8) ,
31984	 => std_logic_vector(to_unsigned(161,8) ,
31985	 => std_logic_vector(to_unsigned(154,8) ,
31986	 => std_logic_vector(to_unsigned(154,8) ,
31987	 => std_logic_vector(to_unsigned(154,8) ,
31988	 => std_logic_vector(to_unsigned(149,8) ,
31989	 => std_logic_vector(to_unsigned(139,8) ,
31990	 => std_logic_vector(to_unsigned(136,8) ,
31991	 => std_logic_vector(to_unsigned(136,8) ,
31992	 => std_logic_vector(to_unsigned(138,8) ,
31993	 => std_logic_vector(to_unsigned(136,8) ,
31994	 => std_logic_vector(to_unsigned(139,8) ,
31995	 => std_logic_vector(to_unsigned(142,8) ,
31996	 => std_logic_vector(to_unsigned(138,8) ,
31997	 => std_logic_vector(to_unsigned(124,8) ,
31998	 => std_logic_vector(to_unsigned(122,8) ,
31999	 => std_logic_vector(to_unsigned(125,8) ,
32000	 => std_logic_vector(to_unsigned(124,8) ,
32001	 => std_logic_vector(to_unsigned(4,8) ,
32002	 => std_logic_vector(to_unsigned(4,8) ,
32003	 => std_logic_vector(to_unsigned(3,8) ,
32004	 => std_logic_vector(to_unsigned(2,8) ,
32005	 => std_logic_vector(to_unsigned(4,8) ,
32006	 => std_logic_vector(to_unsigned(8,8) ,
32007	 => std_logic_vector(to_unsigned(8,8) ,
32008	 => std_logic_vector(to_unsigned(5,8) ,
32009	 => std_logic_vector(to_unsigned(4,8) ,
32010	 => std_logic_vector(to_unsigned(1,8) ,
32011	 => std_logic_vector(to_unsigned(0,8) ,
32012	 => std_logic_vector(to_unsigned(1,8) ,
32013	 => std_logic_vector(to_unsigned(0,8) ,
32014	 => std_logic_vector(to_unsigned(1,8) ,
32015	 => std_logic_vector(to_unsigned(2,8) ,
32016	 => std_logic_vector(to_unsigned(1,8) ,
32017	 => std_logic_vector(to_unsigned(1,8) ,
32018	 => std_logic_vector(to_unsigned(1,8) ,
32019	 => std_logic_vector(to_unsigned(2,8) ,
32020	 => std_logic_vector(to_unsigned(4,8) ,
32021	 => std_logic_vector(to_unsigned(10,8) ,
32022	 => std_logic_vector(to_unsigned(8,8) ,
32023	 => std_logic_vector(to_unsigned(5,8) ,
32024	 => std_logic_vector(to_unsigned(1,8) ,
32025	 => std_logic_vector(to_unsigned(5,8) ,
32026	 => std_logic_vector(to_unsigned(22,8) ,
32027	 => std_logic_vector(to_unsigned(13,8) ,
32028	 => std_logic_vector(to_unsigned(7,8) ,
32029	 => std_logic_vector(to_unsigned(8,8) ,
32030	 => std_logic_vector(to_unsigned(7,8) ,
32031	 => std_logic_vector(to_unsigned(7,8) ,
32032	 => std_logic_vector(to_unsigned(6,8) ,
32033	 => std_logic_vector(to_unsigned(5,8) ,
32034	 => std_logic_vector(to_unsigned(8,8) ,
32035	 => std_logic_vector(to_unsigned(6,8) ,
32036	 => std_logic_vector(to_unsigned(6,8) ,
32037	 => std_logic_vector(to_unsigned(32,8) ,
32038	 => std_logic_vector(to_unsigned(35,8) ,
32039	 => std_logic_vector(to_unsigned(32,8) ,
32040	 => std_logic_vector(to_unsigned(17,8) ,
32041	 => std_logic_vector(to_unsigned(6,8) ,
32042	 => std_logic_vector(to_unsigned(5,8) ,
32043	 => std_logic_vector(to_unsigned(2,8) ,
32044	 => std_logic_vector(to_unsigned(2,8) ,
32045	 => std_logic_vector(to_unsigned(1,8) ,
32046	 => std_logic_vector(to_unsigned(0,8) ,
32047	 => std_logic_vector(to_unsigned(1,8) ,
32048	 => std_logic_vector(to_unsigned(1,8) ,
32049	 => std_logic_vector(to_unsigned(2,8) ,
32050	 => std_logic_vector(to_unsigned(3,8) ,
32051	 => std_logic_vector(to_unsigned(5,8) ,
32052	 => std_logic_vector(to_unsigned(5,8) ,
32053	 => std_logic_vector(to_unsigned(10,8) ,
32054	 => std_logic_vector(to_unsigned(42,8) ,
32055	 => std_logic_vector(to_unsigned(60,8) ,
32056	 => std_logic_vector(to_unsigned(57,8) ,
32057	 => std_logic_vector(to_unsigned(52,8) ,
32058	 => std_logic_vector(to_unsigned(36,8) ,
32059	 => std_logic_vector(to_unsigned(14,8) ,
32060	 => std_logic_vector(to_unsigned(9,8) ,
32061	 => std_logic_vector(to_unsigned(8,8) ,
32062	 => std_logic_vector(to_unsigned(3,8) ,
32063	 => std_logic_vector(to_unsigned(2,8) ,
32064	 => std_logic_vector(to_unsigned(1,8) ,
32065	 => std_logic_vector(to_unsigned(4,8) ,
32066	 => std_logic_vector(to_unsigned(35,8) ,
32067	 => std_logic_vector(to_unsigned(13,8) ,
32068	 => std_logic_vector(to_unsigned(4,8) ,
32069	 => std_logic_vector(to_unsigned(3,8) ,
32070	 => std_logic_vector(to_unsigned(6,8) ,
32071	 => std_logic_vector(to_unsigned(8,8) ,
32072	 => std_logic_vector(to_unsigned(4,8) ,
32073	 => std_logic_vector(to_unsigned(3,8) ,
32074	 => std_logic_vector(to_unsigned(6,8) ,
32075	 => std_logic_vector(to_unsigned(10,8) ,
32076	 => std_logic_vector(to_unsigned(9,8) ,
32077	 => std_logic_vector(to_unsigned(12,8) ,
32078	 => std_logic_vector(to_unsigned(12,8) ,
32079	 => std_logic_vector(to_unsigned(12,8) ,
32080	 => std_logic_vector(to_unsigned(95,8) ,
32081	 => std_logic_vector(to_unsigned(179,8) ,
32082	 => std_logic_vector(to_unsigned(64,8) ,
32083	 => std_logic_vector(to_unsigned(68,8) ,
32084	 => std_logic_vector(to_unsigned(88,8) ,
32085	 => std_logic_vector(to_unsigned(52,8) ,
32086	 => std_logic_vector(to_unsigned(77,8) ,
32087	 => std_logic_vector(to_unsigned(48,8) ,
32088	 => std_logic_vector(to_unsigned(17,8) ,
32089	 => std_logic_vector(to_unsigned(1,8) ,
32090	 => std_logic_vector(to_unsigned(2,8) ,
32091	 => std_logic_vector(to_unsigned(2,8) ,
32092	 => std_logic_vector(to_unsigned(1,8) ,
32093	 => std_logic_vector(to_unsigned(0,8) ,
32094	 => std_logic_vector(to_unsigned(1,8) ,
32095	 => std_logic_vector(to_unsigned(1,8) ,
32096	 => std_logic_vector(to_unsigned(0,8) ,
32097	 => std_logic_vector(to_unsigned(1,8) ,
32098	 => std_logic_vector(to_unsigned(2,8) ,
32099	 => std_logic_vector(to_unsigned(3,8) ,
32100	 => std_logic_vector(to_unsigned(2,8) ,
32101	 => std_logic_vector(to_unsigned(2,8) ,
32102	 => std_logic_vector(to_unsigned(6,8) ,
32103	 => std_logic_vector(to_unsigned(18,8) ,
32104	 => std_logic_vector(to_unsigned(20,8) ,
32105	 => std_logic_vector(to_unsigned(11,8) ,
32106	 => std_logic_vector(to_unsigned(4,8) ,
32107	 => std_logic_vector(to_unsigned(29,8) ,
32108	 => std_logic_vector(to_unsigned(101,8) ,
32109	 => std_logic_vector(to_unsigned(77,8) ,
32110	 => std_logic_vector(to_unsigned(35,8) ,
32111	 => std_logic_vector(to_unsigned(5,8) ,
32112	 => std_logic_vector(to_unsigned(2,8) ,
32113	 => std_logic_vector(to_unsigned(4,8) ,
32114	 => std_logic_vector(to_unsigned(5,8) ,
32115	 => std_logic_vector(to_unsigned(9,8) ,
32116	 => std_logic_vector(to_unsigned(27,8) ,
32117	 => std_logic_vector(to_unsigned(24,8) ,
32118	 => std_logic_vector(to_unsigned(22,8) ,
32119	 => std_logic_vector(to_unsigned(31,8) ,
32120	 => std_logic_vector(to_unsigned(57,8) ,
32121	 => std_logic_vector(to_unsigned(86,8) ,
32122	 => std_logic_vector(to_unsigned(68,8) ,
32123	 => std_logic_vector(to_unsigned(76,8) ,
32124	 => std_logic_vector(to_unsigned(88,8) ,
32125	 => std_logic_vector(to_unsigned(66,8) ,
32126	 => std_logic_vector(to_unsigned(22,8) ,
32127	 => std_logic_vector(to_unsigned(3,8) ,
32128	 => std_logic_vector(to_unsigned(1,8) ,
32129	 => std_logic_vector(to_unsigned(3,8) ,
32130	 => std_logic_vector(to_unsigned(11,8) ,
32131	 => std_logic_vector(to_unsigned(9,8) ,
32132	 => std_logic_vector(to_unsigned(8,8) ,
32133	 => std_logic_vector(to_unsigned(26,8) ,
32134	 => std_logic_vector(to_unsigned(7,8) ,
32135	 => std_logic_vector(to_unsigned(0,8) ,
32136	 => std_logic_vector(to_unsigned(0,8) ,
32137	 => std_logic_vector(to_unsigned(1,8) ,
32138	 => std_logic_vector(to_unsigned(3,8) ,
32139	 => std_logic_vector(to_unsigned(5,8) ,
32140	 => std_logic_vector(to_unsigned(5,8) ,
32141	 => std_logic_vector(to_unsigned(10,8) ,
32142	 => std_logic_vector(to_unsigned(15,8) ,
32143	 => std_logic_vector(to_unsigned(17,8) ,
32144	 => std_logic_vector(to_unsigned(25,8) ,
32145	 => std_logic_vector(to_unsigned(43,8) ,
32146	 => std_logic_vector(to_unsigned(54,8) ,
32147	 => std_logic_vector(to_unsigned(14,8) ,
32148	 => std_logic_vector(to_unsigned(8,8) ,
32149	 => std_logic_vector(to_unsigned(16,8) ,
32150	 => std_logic_vector(to_unsigned(9,8) ,
32151	 => std_logic_vector(to_unsigned(9,8) ,
32152	 => std_logic_vector(to_unsigned(7,8) ,
32153	 => std_logic_vector(to_unsigned(3,8) ,
32154	 => std_logic_vector(to_unsigned(5,8) ,
32155	 => std_logic_vector(to_unsigned(11,8) ,
32156	 => std_logic_vector(to_unsigned(9,8) ,
32157	 => std_logic_vector(to_unsigned(2,8) ,
32158	 => std_logic_vector(to_unsigned(2,8) ,
32159	 => std_logic_vector(to_unsigned(5,8) ,
32160	 => std_logic_vector(to_unsigned(13,8) ,
32161	 => std_logic_vector(to_unsigned(29,8) ,
32162	 => std_logic_vector(to_unsigned(25,8) ,
32163	 => std_logic_vector(to_unsigned(22,8) ,
32164	 => std_logic_vector(to_unsigned(8,8) ,
32165	 => std_logic_vector(to_unsigned(14,8) ,
32166	 => std_logic_vector(to_unsigned(79,8) ,
32167	 => std_logic_vector(to_unsigned(58,8) ,
32168	 => std_logic_vector(to_unsigned(35,8) ,
32169	 => std_logic_vector(to_unsigned(35,8) ,
32170	 => std_logic_vector(to_unsigned(35,8) ,
32171	 => std_logic_vector(to_unsigned(20,8) ,
32172	 => std_logic_vector(to_unsigned(2,8) ,
32173	 => std_logic_vector(to_unsigned(0,8) ,
32174	 => std_logic_vector(to_unsigned(2,8) ,
32175	 => std_logic_vector(to_unsigned(19,8) ,
32176	 => std_logic_vector(to_unsigned(62,8) ,
32177	 => std_logic_vector(to_unsigned(82,8) ,
32178	 => std_logic_vector(to_unsigned(84,8) ,
32179	 => std_logic_vector(to_unsigned(74,8) ,
32180	 => std_logic_vector(to_unsigned(25,8) ,
32181	 => std_logic_vector(to_unsigned(33,8) ,
32182	 => std_logic_vector(to_unsigned(19,8) ,
32183	 => std_logic_vector(to_unsigned(1,8) ,
32184	 => std_logic_vector(to_unsigned(0,8) ,
32185	 => std_logic_vector(to_unsigned(0,8) ,
32186	 => std_logic_vector(to_unsigned(8,8) ,
32187	 => std_logic_vector(to_unsigned(35,8) ,
32188	 => std_logic_vector(to_unsigned(76,8) ,
32189	 => std_logic_vector(to_unsigned(82,8) ,
32190	 => std_logic_vector(to_unsigned(47,8) ,
32191	 => std_logic_vector(to_unsigned(31,8) ,
32192	 => std_logic_vector(to_unsigned(19,8) ,
32193	 => std_logic_vector(to_unsigned(4,8) ,
32194	 => std_logic_vector(to_unsigned(64,8) ,
32195	 => std_logic_vector(to_unsigned(168,8) ,
32196	 => std_logic_vector(to_unsigned(144,8) ,
32197	 => std_logic_vector(to_unsigned(156,8) ,
32198	 => std_logic_vector(to_unsigned(168,8) ,
32199	 => std_logic_vector(to_unsigned(50,8) ,
32200	 => std_logic_vector(to_unsigned(8,8) ,
32201	 => std_logic_vector(to_unsigned(24,8) ,
32202	 => std_logic_vector(to_unsigned(22,8) ,
32203	 => std_logic_vector(to_unsigned(45,8) ,
32204	 => std_logic_vector(to_unsigned(81,8) ,
32205	 => std_logic_vector(to_unsigned(88,8) ,
32206	 => std_logic_vector(to_unsigned(81,8) ,
32207	 => std_logic_vector(to_unsigned(63,8) ,
32208	 => std_logic_vector(to_unsigned(71,8) ,
32209	 => std_logic_vector(to_unsigned(149,8) ,
32210	 => std_logic_vector(to_unsigned(156,8) ,
32211	 => std_logic_vector(to_unsigned(152,8) ,
32212	 => std_logic_vector(to_unsigned(154,8) ,
32213	 => std_logic_vector(to_unsigned(159,8) ,
32214	 => std_logic_vector(to_unsigned(159,8) ,
32215	 => std_logic_vector(to_unsigned(157,8) ,
32216	 => std_logic_vector(to_unsigned(156,8) ,
32217	 => std_logic_vector(to_unsigned(157,8) ,
32218	 => std_logic_vector(to_unsigned(156,8) ,
32219	 => std_logic_vector(to_unsigned(156,8) ,
32220	 => std_logic_vector(to_unsigned(154,8) ,
32221	 => std_logic_vector(to_unsigned(154,8) ,
32222	 => std_logic_vector(to_unsigned(147,8) ,
32223	 => std_logic_vector(to_unsigned(152,8) ,
32224	 => std_logic_vector(to_unsigned(73,8) ,
32225	 => std_logic_vector(to_unsigned(7,8) ,
32226	 => std_logic_vector(to_unsigned(6,8) ,
32227	 => std_logic_vector(to_unsigned(2,8) ,
32228	 => std_logic_vector(to_unsigned(1,8) ,
32229	 => std_logic_vector(to_unsigned(6,8) ,
32230	 => std_logic_vector(to_unsigned(5,8) ,
32231	 => std_logic_vector(to_unsigned(19,8) ,
32232	 => std_logic_vector(to_unsigned(45,8) ,
32233	 => std_logic_vector(to_unsigned(53,8) ,
32234	 => std_logic_vector(to_unsigned(25,8) ,
32235	 => std_logic_vector(to_unsigned(8,8) ,
32236	 => std_logic_vector(to_unsigned(24,8) ,
32237	 => std_logic_vector(to_unsigned(41,8) ,
32238	 => std_logic_vector(to_unsigned(15,8) ,
32239	 => std_logic_vector(to_unsigned(92,8) ,
32240	 => std_logic_vector(to_unsigned(188,8) ,
32241	 => std_logic_vector(to_unsigned(147,8) ,
32242	 => std_logic_vector(to_unsigned(149,8) ,
32243	 => std_logic_vector(to_unsigned(171,8) ,
32244	 => std_logic_vector(to_unsigned(66,8) ,
32245	 => std_logic_vector(to_unsigned(2,8) ,
32246	 => std_logic_vector(to_unsigned(8,8) ,
32247	 => std_logic_vector(to_unsigned(119,8) ,
32248	 => std_logic_vector(to_unsigned(183,8) ,
32249	 => std_logic_vector(to_unsigned(166,8) ,
32250	 => std_logic_vector(to_unsigned(177,8) ,
32251	 => std_logic_vector(to_unsigned(171,8) ,
32252	 => std_logic_vector(to_unsigned(181,8) ,
32253	 => std_logic_vector(to_unsigned(183,8) ,
32254	 => std_logic_vector(to_unsigned(200,8) ,
32255	 => std_logic_vector(to_unsigned(136,8) ,
32256	 => std_logic_vector(to_unsigned(4,8) ,
32257	 => std_logic_vector(to_unsigned(1,8) ,
32258	 => std_logic_vector(to_unsigned(3,8) ,
32259	 => std_logic_vector(to_unsigned(10,8) ,
32260	 => std_logic_vector(to_unsigned(12,8) ,
32261	 => std_logic_vector(to_unsigned(6,8) ,
32262	 => std_logic_vector(to_unsigned(13,8) ,
32263	 => std_logic_vector(to_unsigned(15,8) ,
32264	 => std_logic_vector(to_unsigned(27,8) ,
32265	 => std_logic_vector(to_unsigned(92,8) ,
32266	 => std_logic_vector(to_unsigned(130,8) ,
32267	 => std_logic_vector(to_unsigned(125,8) ,
32268	 => std_logic_vector(to_unsigned(32,8) ,
32269	 => std_logic_vector(to_unsigned(8,8) ,
32270	 => std_logic_vector(to_unsigned(101,8) ,
32271	 => std_logic_vector(to_unsigned(154,8) ,
32272	 => std_logic_vector(to_unsigned(72,8) ,
32273	 => std_logic_vector(to_unsigned(11,8) ,
32274	 => std_logic_vector(to_unsigned(3,8) ,
32275	 => std_logic_vector(to_unsigned(1,8) ,
32276	 => std_logic_vector(to_unsigned(6,8) ,
32277	 => std_logic_vector(to_unsigned(7,8) ,
32278	 => std_logic_vector(to_unsigned(4,8) ,
32279	 => std_logic_vector(to_unsigned(5,8) ,
32280	 => std_logic_vector(to_unsigned(5,8) ,
32281	 => std_logic_vector(to_unsigned(6,8) ,
32282	 => std_logic_vector(to_unsigned(5,8) ,
32283	 => std_logic_vector(to_unsigned(5,8) ,
32284	 => std_logic_vector(to_unsigned(6,8) ,
32285	 => std_logic_vector(to_unsigned(4,8) ,
32286	 => std_logic_vector(to_unsigned(5,8) ,
32287	 => std_logic_vector(to_unsigned(5,8) ,
32288	 => std_logic_vector(to_unsigned(4,8) ,
32289	 => std_logic_vector(to_unsigned(4,8) ,
32290	 => std_logic_vector(to_unsigned(3,8) ,
32291	 => std_logic_vector(to_unsigned(1,8) ,
32292	 => std_logic_vector(to_unsigned(2,8) ,
32293	 => std_logic_vector(to_unsigned(7,8) ,
32294	 => std_logic_vector(to_unsigned(7,8) ,
32295	 => std_logic_vector(to_unsigned(5,8) ,
32296	 => std_logic_vector(to_unsigned(30,8) ,
32297	 => std_logic_vector(to_unsigned(90,8) ,
32298	 => std_logic_vector(to_unsigned(119,8) ,
32299	 => std_logic_vector(to_unsigned(134,8) ,
32300	 => std_logic_vector(to_unsigned(152,8) ,
32301	 => std_logic_vector(to_unsigned(151,8) ,
32302	 => std_logic_vector(to_unsigned(164,8) ,
32303	 => std_logic_vector(to_unsigned(159,8) ,
32304	 => std_logic_vector(to_unsigned(157,8) ,
32305	 => std_logic_vector(to_unsigned(151,8) ,
32306	 => std_logic_vector(to_unsigned(146,8) ,
32307	 => std_logic_vector(to_unsigned(149,8) ,
32308	 => std_logic_vector(to_unsigned(146,8) ,
32309	 => std_logic_vector(to_unsigned(133,8) ,
32310	 => std_logic_vector(to_unsigned(134,8) ,
32311	 => std_logic_vector(to_unsigned(139,8) ,
32312	 => std_logic_vector(to_unsigned(141,8) ,
32313	 => std_logic_vector(to_unsigned(136,8) ,
32314	 => std_logic_vector(to_unsigned(139,8) ,
32315	 => std_logic_vector(to_unsigned(139,8) ,
32316	 => std_logic_vector(to_unsigned(128,8) ,
32317	 => std_logic_vector(to_unsigned(128,8) ,
32318	 => std_logic_vector(to_unsigned(128,8) ,
32319	 => std_logic_vector(to_unsigned(131,8) ,
32320	 => std_logic_vector(to_unsigned(134,8) ,
32321	 => std_logic_vector(to_unsigned(6,8) ,
32322	 => std_logic_vector(to_unsigned(4,8) ,
32323	 => std_logic_vector(to_unsigned(4,8) ,
32324	 => std_logic_vector(to_unsigned(2,8) ,
32325	 => std_logic_vector(to_unsigned(4,8) ,
32326	 => std_logic_vector(to_unsigned(7,8) ,
32327	 => std_logic_vector(to_unsigned(6,8) ,
32328	 => std_logic_vector(to_unsigned(3,8) ,
32329	 => std_logic_vector(to_unsigned(3,8) ,
32330	 => std_logic_vector(to_unsigned(2,8) ,
32331	 => std_logic_vector(to_unsigned(1,8) ,
32332	 => std_logic_vector(to_unsigned(1,8) ,
32333	 => std_logic_vector(to_unsigned(1,8) ,
32334	 => std_logic_vector(to_unsigned(1,8) ,
32335	 => std_logic_vector(to_unsigned(1,8) ,
32336	 => std_logic_vector(to_unsigned(1,8) ,
32337	 => std_logic_vector(to_unsigned(1,8) ,
32338	 => std_logic_vector(to_unsigned(1,8) ,
32339	 => std_logic_vector(to_unsigned(2,8) ,
32340	 => std_logic_vector(to_unsigned(8,8) ,
32341	 => std_logic_vector(to_unsigned(13,8) ,
32342	 => std_logic_vector(to_unsigned(6,8) ,
32343	 => std_logic_vector(to_unsigned(2,8) ,
32344	 => std_logic_vector(to_unsigned(1,8) ,
32345	 => std_logic_vector(to_unsigned(1,8) ,
32346	 => std_logic_vector(to_unsigned(13,8) ,
32347	 => std_logic_vector(to_unsigned(6,8) ,
32348	 => std_logic_vector(to_unsigned(4,8) ,
32349	 => std_logic_vector(to_unsigned(4,8) ,
32350	 => std_logic_vector(to_unsigned(4,8) ,
32351	 => std_logic_vector(to_unsigned(4,8) ,
32352	 => std_logic_vector(to_unsigned(6,8) ,
32353	 => std_logic_vector(to_unsigned(12,8) ,
32354	 => std_logic_vector(to_unsigned(19,8) ,
32355	 => std_logic_vector(to_unsigned(7,8) ,
32356	 => std_logic_vector(to_unsigned(10,8) ,
32357	 => std_logic_vector(to_unsigned(37,8) ,
32358	 => std_logic_vector(to_unsigned(30,8) ,
32359	 => std_logic_vector(to_unsigned(31,8) ,
32360	 => std_logic_vector(to_unsigned(20,8) ,
32361	 => std_logic_vector(to_unsigned(14,8) ,
32362	 => std_logic_vector(to_unsigned(8,8) ,
32363	 => std_logic_vector(to_unsigned(4,8) ,
32364	 => std_logic_vector(to_unsigned(1,8) ,
32365	 => std_logic_vector(to_unsigned(0,8) ,
32366	 => std_logic_vector(to_unsigned(1,8) ,
32367	 => std_logic_vector(to_unsigned(3,8) ,
32368	 => std_logic_vector(to_unsigned(2,8) ,
32369	 => std_logic_vector(to_unsigned(1,8) ,
32370	 => std_logic_vector(to_unsigned(0,8) ,
32371	 => std_logic_vector(to_unsigned(0,8) ,
32372	 => std_logic_vector(to_unsigned(0,8) ,
32373	 => std_logic_vector(to_unsigned(4,8) ,
32374	 => std_logic_vector(to_unsigned(61,8) ,
32375	 => std_logic_vector(to_unsigned(81,8) ,
32376	 => std_logic_vector(to_unsigned(64,8) ,
32377	 => std_logic_vector(to_unsigned(51,8) ,
32378	 => std_logic_vector(to_unsigned(40,8) ,
32379	 => std_logic_vector(to_unsigned(23,8) ,
32380	 => std_logic_vector(to_unsigned(8,8) ,
32381	 => std_logic_vector(to_unsigned(3,8) ,
32382	 => std_logic_vector(to_unsigned(3,8) ,
32383	 => std_logic_vector(to_unsigned(2,8) ,
32384	 => std_logic_vector(to_unsigned(1,8) ,
32385	 => std_logic_vector(to_unsigned(0,8) ,
32386	 => std_logic_vector(to_unsigned(1,8) ,
32387	 => std_logic_vector(to_unsigned(7,8) ,
32388	 => std_logic_vector(to_unsigned(8,8) ,
32389	 => std_logic_vector(to_unsigned(3,8) ,
32390	 => std_logic_vector(to_unsigned(1,8) ,
32391	 => std_logic_vector(to_unsigned(1,8) ,
32392	 => std_logic_vector(to_unsigned(1,8) ,
32393	 => std_logic_vector(to_unsigned(3,8) ,
32394	 => std_logic_vector(to_unsigned(11,8) ,
32395	 => std_logic_vector(to_unsigned(10,8) ,
32396	 => std_logic_vector(to_unsigned(6,8) ,
32397	 => std_logic_vector(to_unsigned(10,8) ,
32398	 => std_logic_vector(to_unsigned(10,8) ,
32399	 => std_logic_vector(to_unsigned(17,8) ,
32400	 => std_logic_vector(to_unsigned(99,8) ,
32401	 => std_logic_vector(to_unsigned(157,8) ,
32402	 => std_logic_vector(to_unsigned(82,8) ,
32403	 => std_logic_vector(to_unsigned(109,8) ,
32404	 => std_logic_vector(to_unsigned(127,8) ,
32405	 => std_logic_vector(to_unsigned(62,8) ,
32406	 => std_logic_vector(to_unsigned(56,8) ,
32407	 => std_logic_vector(to_unsigned(65,8) ,
32408	 => std_logic_vector(to_unsigned(24,8) ,
32409	 => std_logic_vector(to_unsigned(0,8) ,
32410	 => std_logic_vector(to_unsigned(2,8) ,
32411	 => std_logic_vector(to_unsigned(2,8) ,
32412	 => std_logic_vector(to_unsigned(1,8) ,
32413	 => std_logic_vector(to_unsigned(1,8) ,
32414	 => std_logic_vector(to_unsigned(1,8) ,
32415	 => std_logic_vector(to_unsigned(0,8) ,
32416	 => std_logic_vector(to_unsigned(2,8) ,
32417	 => std_logic_vector(to_unsigned(4,8) ,
32418	 => std_logic_vector(to_unsigned(6,8) ,
32419	 => std_logic_vector(to_unsigned(5,8) ,
32420	 => std_logic_vector(to_unsigned(4,8) ,
32421	 => std_logic_vector(to_unsigned(12,8) ,
32422	 => std_logic_vector(to_unsigned(20,8) ,
32423	 => std_logic_vector(to_unsigned(22,8) ,
32424	 => std_logic_vector(to_unsigned(24,8) ,
32425	 => std_logic_vector(to_unsigned(13,8) ,
32426	 => std_logic_vector(to_unsigned(7,8) ,
32427	 => std_logic_vector(to_unsigned(31,8) ,
32428	 => std_logic_vector(to_unsigned(79,8) ,
32429	 => std_logic_vector(to_unsigned(60,8) ,
32430	 => std_logic_vector(to_unsigned(20,8) ,
32431	 => std_logic_vector(to_unsigned(10,8) ,
32432	 => std_logic_vector(to_unsigned(13,8) ,
32433	 => std_logic_vector(to_unsigned(15,8) ,
32434	 => std_logic_vector(to_unsigned(18,8) ,
32435	 => std_logic_vector(to_unsigned(13,8) ,
32436	 => std_logic_vector(to_unsigned(35,8) ,
32437	 => std_logic_vector(to_unsigned(38,8) ,
32438	 => std_logic_vector(to_unsigned(20,8) ,
32439	 => std_logic_vector(to_unsigned(35,8) ,
32440	 => std_logic_vector(to_unsigned(45,8) ,
32441	 => std_logic_vector(to_unsigned(90,8) ,
32442	 => std_logic_vector(to_unsigned(57,8) ,
32443	 => std_logic_vector(to_unsigned(10,8) ,
32444	 => std_logic_vector(to_unsigned(10,8) ,
32445	 => std_logic_vector(to_unsigned(4,8) ,
32446	 => std_logic_vector(to_unsigned(1,8) ,
32447	 => std_logic_vector(to_unsigned(1,8) ,
32448	 => std_logic_vector(to_unsigned(1,8) ,
32449	 => std_logic_vector(to_unsigned(4,8) ,
32450	 => std_logic_vector(to_unsigned(17,8) ,
32451	 => std_logic_vector(to_unsigned(10,8) ,
32452	 => std_logic_vector(to_unsigned(7,8) ,
32453	 => std_logic_vector(to_unsigned(26,8) ,
32454	 => std_logic_vector(to_unsigned(22,8) ,
32455	 => std_logic_vector(to_unsigned(17,8) ,
32456	 => std_logic_vector(to_unsigned(33,8) ,
32457	 => std_logic_vector(to_unsigned(47,8) ,
32458	 => std_logic_vector(to_unsigned(65,8) ,
32459	 => std_logic_vector(to_unsigned(85,8) ,
32460	 => std_logic_vector(to_unsigned(104,8) ,
32461	 => std_logic_vector(to_unsigned(125,8) ,
32462	 => std_logic_vector(to_unsigned(139,8) ,
32463	 => std_logic_vector(to_unsigned(147,8) ,
32464	 => std_logic_vector(to_unsigned(156,8) ,
32465	 => std_logic_vector(to_unsigned(147,8) ,
32466	 => std_logic_vector(to_unsigned(146,8) ,
32467	 => std_logic_vector(to_unsigned(50,8) ,
32468	 => std_logic_vector(to_unsigned(12,8) ,
32469	 => std_logic_vector(to_unsigned(8,8) ,
32470	 => std_logic_vector(to_unsigned(4,8) ,
32471	 => std_logic_vector(to_unsigned(6,8) ,
32472	 => std_logic_vector(to_unsigned(5,8) ,
32473	 => std_logic_vector(to_unsigned(3,8) ,
32474	 => std_logic_vector(to_unsigned(1,8) ,
32475	 => std_logic_vector(to_unsigned(2,8) ,
32476	 => std_logic_vector(to_unsigned(2,8) ,
32477	 => std_logic_vector(to_unsigned(2,8) ,
32478	 => std_logic_vector(to_unsigned(5,8) ,
32479	 => std_logic_vector(to_unsigned(24,8) ,
32480	 => std_logic_vector(to_unsigned(48,8) ,
32481	 => std_logic_vector(to_unsigned(32,8) ,
32482	 => std_logic_vector(to_unsigned(13,8) ,
32483	 => std_logic_vector(to_unsigned(10,8) ,
32484	 => std_logic_vector(to_unsigned(6,8) ,
32485	 => std_logic_vector(to_unsigned(5,8) ,
32486	 => std_logic_vector(to_unsigned(51,8) ,
32487	 => std_logic_vector(to_unsigned(60,8) ,
32488	 => std_logic_vector(to_unsigned(42,8) ,
32489	 => std_logic_vector(to_unsigned(54,8) ,
32490	 => std_logic_vector(to_unsigned(33,8) ,
32491	 => std_logic_vector(to_unsigned(5,8) ,
32492	 => std_logic_vector(to_unsigned(1,8) ,
32493	 => std_logic_vector(to_unsigned(2,8) ,
32494	 => std_logic_vector(to_unsigned(1,8) ,
32495	 => std_logic_vector(to_unsigned(5,8) ,
32496	 => std_logic_vector(to_unsigned(24,8) ,
32497	 => std_logic_vector(to_unsigned(32,8) ,
32498	 => std_logic_vector(to_unsigned(36,8) ,
32499	 => std_logic_vector(to_unsigned(20,8) ,
32500	 => std_logic_vector(to_unsigned(8,8) ,
32501	 => std_logic_vector(to_unsigned(3,8) ,
32502	 => std_logic_vector(to_unsigned(1,8) ,
32503	 => std_logic_vector(to_unsigned(0,8) ,
32504	 => std_logic_vector(to_unsigned(1,8) ,
32505	 => std_logic_vector(to_unsigned(1,8) ,
32506	 => std_logic_vector(to_unsigned(2,8) ,
32507	 => std_logic_vector(to_unsigned(37,8) ,
32508	 => std_logic_vector(to_unsigned(91,8) ,
32509	 => std_logic_vector(to_unsigned(88,8) ,
32510	 => std_logic_vector(to_unsigned(101,8) ,
32511	 => std_logic_vector(to_unsigned(47,8) ,
32512	 => std_logic_vector(to_unsigned(18,8) ,
32513	 => std_logic_vector(to_unsigned(5,8) ,
32514	 => std_logic_vector(to_unsigned(32,8) ,
32515	 => std_logic_vector(to_unsigned(152,8) ,
32516	 => std_logic_vector(to_unsigned(144,8) ,
32517	 => std_logic_vector(to_unsigned(144,8) ,
32518	 => std_logic_vector(to_unsigned(166,8) ,
32519	 => std_logic_vector(to_unsigned(29,8) ,
32520	 => std_logic_vector(to_unsigned(1,8) ,
32521	 => std_logic_vector(to_unsigned(6,8) ,
32522	 => std_logic_vector(to_unsigned(15,8) ,
32523	 => std_logic_vector(to_unsigned(68,8) ,
32524	 => std_logic_vector(to_unsigned(99,8) ,
32525	 => std_logic_vector(to_unsigned(70,8) ,
32526	 => std_logic_vector(to_unsigned(61,8) ,
32527	 => std_logic_vector(to_unsigned(45,8) ,
32528	 => std_logic_vector(to_unsigned(30,8) ,
32529	 => std_logic_vector(to_unsigned(112,8) ,
32530	 => std_logic_vector(to_unsigned(170,8) ,
32531	 => std_logic_vector(to_unsigned(152,8) ,
32532	 => std_logic_vector(to_unsigned(152,8) ,
32533	 => std_logic_vector(to_unsigned(156,8) ,
32534	 => std_logic_vector(to_unsigned(161,8) ,
32535	 => std_logic_vector(to_unsigned(157,8) ,
32536	 => std_logic_vector(to_unsigned(152,8) ,
32537	 => std_logic_vector(to_unsigned(154,8) ,
32538	 => std_logic_vector(to_unsigned(154,8) ,
32539	 => std_logic_vector(to_unsigned(154,8) ,
32540	 => std_logic_vector(to_unsigned(154,8) ,
32541	 => std_logic_vector(to_unsigned(156,8) ,
32542	 => std_logic_vector(to_unsigned(159,8) ,
32543	 => std_logic_vector(to_unsigned(142,8) ,
32544	 => std_logic_vector(to_unsigned(25,8) ,
32545	 => std_logic_vector(to_unsigned(0,8) ,
32546	 => std_logic_vector(to_unsigned(16,8) ,
32547	 => std_logic_vector(to_unsigned(24,8) ,
32548	 => std_logic_vector(to_unsigned(1,8) ,
32549	 => std_logic_vector(to_unsigned(3,8) ,
32550	 => std_logic_vector(to_unsigned(4,8) ,
32551	 => std_logic_vector(to_unsigned(2,8) ,
32552	 => std_logic_vector(to_unsigned(8,8) ,
32553	 => std_logic_vector(to_unsigned(49,8) ,
32554	 => std_logic_vector(to_unsigned(41,8) ,
32555	 => std_logic_vector(to_unsigned(19,8) ,
32556	 => std_logic_vector(to_unsigned(35,8) ,
32557	 => std_logic_vector(to_unsigned(35,8) ,
32558	 => std_logic_vector(to_unsigned(24,8) ,
32559	 => std_logic_vector(to_unsigned(125,8) ,
32560	 => std_logic_vector(to_unsigned(159,8) ,
32561	 => std_logic_vector(to_unsigned(149,8) ,
32562	 => std_logic_vector(to_unsigned(146,8) ,
32563	 => std_logic_vector(to_unsigned(164,8) ,
32564	 => std_logic_vector(to_unsigned(60,8) ,
32565	 => std_logic_vector(to_unsigned(3,8) ,
32566	 => std_logic_vector(to_unsigned(12,8) ,
32567	 => std_logic_vector(to_unsigned(114,8) ,
32568	 => std_logic_vector(to_unsigned(156,8) ,
32569	 => std_logic_vector(to_unsigned(146,8) ,
32570	 => std_logic_vector(to_unsigned(152,8) ,
32571	 => std_logic_vector(to_unsigned(146,8) ,
32572	 => std_logic_vector(to_unsigned(154,8) ,
32573	 => std_logic_vector(to_unsigned(151,8) ,
32574	 => std_logic_vector(to_unsigned(166,8) ,
32575	 => std_logic_vector(to_unsigned(124,8) ,
32576	 => std_logic_vector(to_unsigned(8,8) ,
32577	 => std_logic_vector(to_unsigned(0,8) ,
32578	 => std_logic_vector(to_unsigned(1,8) ,
32579	 => std_logic_vector(to_unsigned(7,8) ,
32580	 => std_logic_vector(to_unsigned(13,8) ,
32581	 => std_logic_vector(to_unsigned(9,8) ,
32582	 => std_logic_vector(to_unsigned(9,8) ,
32583	 => std_logic_vector(to_unsigned(9,8) ,
32584	 => std_logic_vector(to_unsigned(21,8) ,
32585	 => std_logic_vector(to_unsigned(118,8) ,
32586	 => std_logic_vector(to_unsigned(186,8) ,
32587	 => std_logic_vector(to_unsigned(131,8) ,
32588	 => std_logic_vector(to_unsigned(39,8) ,
32589	 => std_logic_vector(to_unsigned(69,8) ,
32590	 => std_logic_vector(to_unsigned(147,8) ,
32591	 => std_logic_vector(to_unsigned(138,8) ,
32592	 => std_logic_vector(to_unsigned(111,8) ,
32593	 => std_logic_vector(to_unsigned(24,8) ,
32594	 => std_logic_vector(to_unsigned(1,8) ,
32595	 => std_logic_vector(to_unsigned(1,8) ,
32596	 => std_logic_vector(to_unsigned(2,8) ,
32597	 => std_logic_vector(to_unsigned(3,8) ,
32598	 => std_logic_vector(to_unsigned(5,8) ,
32599	 => std_logic_vector(to_unsigned(4,8) ,
32600	 => std_logic_vector(to_unsigned(4,8) ,
32601	 => std_logic_vector(to_unsigned(6,8) ,
32602	 => std_logic_vector(to_unsigned(5,8) ,
32603	 => std_logic_vector(to_unsigned(4,8) ,
32604	 => std_logic_vector(to_unsigned(6,8) ,
32605	 => std_logic_vector(to_unsigned(8,8) ,
32606	 => std_logic_vector(to_unsigned(5,8) ,
32607	 => std_logic_vector(to_unsigned(4,8) ,
32608	 => std_logic_vector(to_unsigned(5,8) ,
32609	 => std_logic_vector(to_unsigned(5,8) ,
32610	 => std_logic_vector(to_unsigned(4,8) ,
32611	 => std_logic_vector(to_unsigned(5,8) ,
32612	 => std_logic_vector(to_unsigned(2,8) ,
32613	 => std_logic_vector(to_unsigned(3,8) ,
32614	 => std_logic_vector(to_unsigned(3,8) ,
32615	 => std_logic_vector(to_unsigned(6,8) ,
32616	 => std_logic_vector(to_unsigned(51,8) ,
32617	 => std_logic_vector(to_unsigned(122,8) ,
32618	 => std_logic_vector(to_unsigned(130,8) ,
32619	 => std_logic_vector(to_unsigned(131,8) ,
32620	 => std_logic_vector(to_unsigned(147,8) ,
32621	 => std_logic_vector(to_unsigned(154,8) ,
32622	 => std_logic_vector(to_unsigned(163,8) ,
32623	 => std_logic_vector(to_unsigned(152,8) ,
32624	 => std_logic_vector(to_unsigned(141,8) ,
32625	 => std_logic_vector(to_unsigned(131,8) ,
32626	 => std_logic_vector(to_unsigned(127,8) ,
32627	 => std_logic_vector(to_unsigned(131,8) ,
32628	 => std_logic_vector(to_unsigned(138,8) ,
32629	 => std_logic_vector(to_unsigned(130,8) ,
32630	 => std_logic_vector(to_unsigned(146,8) ,
32631	 => std_logic_vector(to_unsigned(159,8) ,
32632	 => std_logic_vector(to_unsigned(159,8) ,
32633	 => std_logic_vector(to_unsigned(154,8) ,
32634	 => std_logic_vector(to_unsigned(156,8) ,
32635	 => std_logic_vector(to_unsigned(154,8) ,
32636	 => std_logic_vector(to_unsigned(142,8) ,
32637	 => std_logic_vector(to_unsigned(151,8) ,
32638	 => std_logic_vector(to_unsigned(144,8) ,
32639	 => std_logic_vector(to_unsigned(144,8) ,
32640	 => std_logic_vector(to_unsigned(152,8) ,
32641	 => std_logic_vector(to_unsigned(6,8) ,
32642	 => std_logic_vector(to_unsigned(4,8) ,
32643	 => std_logic_vector(to_unsigned(3,8) ,
32644	 => std_logic_vector(to_unsigned(4,8) ,
32645	 => std_logic_vector(to_unsigned(4,8) ,
32646	 => std_logic_vector(to_unsigned(4,8) ,
32647	 => std_logic_vector(to_unsigned(4,8) ,
32648	 => std_logic_vector(to_unsigned(1,8) ,
32649	 => std_logic_vector(to_unsigned(1,8) ,
32650	 => std_logic_vector(to_unsigned(2,8) ,
32651	 => std_logic_vector(to_unsigned(2,8) ,
32652	 => std_logic_vector(to_unsigned(2,8) ,
32653	 => std_logic_vector(to_unsigned(1,8) ,
32654	 => std_logic_vector(to_unsigned(1,8) ,
32655	 => std_logic_vector(to_unsigned(1,8) ,
32656	 => std_logic_vector(to_unsigned(1,8) ,
32657	 => std_logic_vector(to_unsigned(1,8) ,
32658	 => std_logic_vector(to_unsigned(2,8) ,
32659	 => std_logic_vector(to_unsigned(4,8) ,
32660	 => std_logic_vector(to_unsigned(5,8) ,
32661	 => std_logic_vector(to_unsigned(9,8) ,
32662	 => std_logic_vector(to_unsigned(5,8) ,
32663	 => std_logic_vector(to_unsigned(2,8) ,
32664	 => std_logic_vector(to_unsigned(1,8) ,
32665	 => std_logic_vector(to_unsigned(0,8) ,
32666	 => std_logic_vector(to_unsigned(6,8) ,
32667	 => std_logic_vector(to_unsigned(9,8) ,
32668	 => std_logic_vector(to_unsigned(5,8) ,
32669	 => std_logic_vector(to_unsigned(4,8) ,
32670	 => std_logic_vector(to_unsigned(4,8) ,
32671	 => std_logic_vector(to_unsigned(3,8) ,
32672	 => std_logic_vector(to_unsigned(1,8) ,
32673	 => std_logic_vector(to_unsigned(2,8) ,
32674	 => std_logic_vector(to_unsigned(3,8) ,
32675	 => std_logic_vector(to_unsigned(2,8) ,
32676	 => std_logic_vector(to_unsigned(20,8) ,
32677	 => std_logic_vector(to_unsigned(44,8) ,
32678	 => std_logic_vector(to_unsigned(34,8) ,
32679	 => std_logic_vector(to_unsigned(37,8) ,
32680	 => std_logic_vector(to_unsigned(30,8) ,
32681	 => std_logic_vector(to_unsigned(14,8) ,
32682	 => std_logic_vector(to_unsigned(12,8) ,
32683	 => std_logic_vector(to_unsigned(8,8) ,
32684	 => std_logic_vector(to_unsigned(2,8) ,
32685	 => std_logic_vector(to_unsigned(1,8) ,
32686	 => std_logic_vector(to_unsigned(7,8) ,
32687	 => std_logic_vector(to_unsigned(6,8) ,
32688	 => std_logic_vector(to_unsigned(1,8) ,
32689	 => std_logic_vector(to_unsigned(0,8) ,
32690	 => std_logic_vector(to_unsigned(0,8) ,
32691	 => std_logic_vector(to_unsigned(0,8) ,
32692	 => std_logic_vector(to_unsigned(2,8) ,
32693	 => std_logic_vector(to_unsigned(14,8) ,
32694	 => std_logic_vector(to_unsigned(55,8) ,
32695	 => std_logic_vector(to_unsigned(71,8) ,
32696	 => std_logic_vector(to_unsigned(59,8) ,
32697	 => std_logic_vector(to_unsigned(51,8) ,
32698	 => std_logic_vector(to_unsigned(48,8) ,
32699	 => std_logic_vector(to_unsigned(32,8) ,
32700	 => std_logic_vector(to_unsigned(16,8) ,
32701	 => std_logic_vector(to_unsigned(11,8) ,
32702	 => std_logic_vector(to_unsigned(3,8) ,
32703	 => std_logic_vector(to_unsigned(1,8) ,
32704	 => std_logic_vector(to_unsigned(0,8) ,
32705	 => std_logic_vector(to_unsigned(1,8) ,
32706	 => std_logic_vector(to_unsigned(0,8) ,
32707	 => std_logic_vector(to_unsigned(1,8) ,
32708	 => std_logic_vector(to_unsigned(4,8) ,
32709	 => std_logic_vector(to_unsigned(9,8) ,
32710	 => std_logic_vector(to_unsigned(3,8) ,
32711	 => std_logic_vector(to_unsigned(2,8) ,
32712	 => std_logic_vector(to_unsigned(4,8) ,
32713	 => std_logic_vector(to_unsigned(10,8) ,
32714	 => std_logic_vector(to_unsigned(10,8) ,
32715	 => std_logic_vector(to_unsigned(5,8) ,
32716	 => std_logic_vector(to_unsigned(8,8) ,
32717	 => std_logic_vector(to_unsigned(9,8) ,
32718	 => std_logic_vector(to_unsigned(10,8) ,
32719	 => std_logic_vector(to_unsigned(14,8) ,
32720	 => std_logic_vector(to_unsigned(14,8) ,
32721	 => std_logic_vector(to_unsigned(16,8) ,
32722	 => std_logic_vector(to_unsigned(20,8) ,
32723	 => std_logic_vector(to_unsigned(30,8) ,
32724	 => std_logic_vector(to_unsigned(41,8) ,
32725	 => std_logic_vector(to_unsigned(37,8) ,
32726	 => std_logic_vector(to_unsigned(41,8) ,
32727	 => std_logic_vector(to_unsigned(80,8) ,
32728	 => std_logic_vector(to_unsigned(52,8) ,
32729	 => std_logic_vector(to_unsigned(8,8) ,
32730	 => std_logic_vector(to_unsigned(1,8) ,
32731	 => std_logic_vector(to_unsigned(1,8) ,
32732	 => std_logic_vector(to_unsigned(1,8) ,
32733	 => std_logic_vector(to_unsigned(1,8) ,
32734	 => std_logic_vector(to_unsigned(0,8) ,
32735	 => std_logic_vector(to_unsigned(1,8) ,
32736	 => std_logic_vector(to_unsigned(7,8) ,
32737	 => std_logic_vector(to_unsigned(7,8) ,
32738	 => std_logic_vector(to_unsigned(3,8) ,
32739	 => std_logic_vector(to_unsigned(2,8) ,
32740	 => std_logic_vector(to_unsigned(10,8) ,
32741	 => std_logic_vector(to_unsigned(21,8) ,
32742	 => std_logic_vector(to_unsigned(18,8) ,
32743	 => std_logic_vector(to_unsigned(21,8) ,
32744	 => std_logic_vector(to_unsigned(17,8) ,
32745	 => std_logic_vector(to_unsigned(9,8) ,
32746	 => std_logic_vector(to_unsigned(20,8) ,
32747	 => std_logic_vector(to_unsigned(77,8) ,
32748	 => std_logic_vector(to_unsigned(81,8) ,
32749	 => std_logic_vector(to_unsigned(44,8) ,
32750	 => std_logic_vector(to_unsigned(13,8) ,
32751	 => std_logic_vector(to_unsigned(13,8) ,
32752	 => std_logic_vector(to_unsigned(24,8) ,
32753	 => std_logic_vector(to_unsigned(24,8) ,
32754	 => std_logic_vector(to_unsigned(27,8) ,
32755	 => std_logic_vector(to_unsigned(16,8) ,
32756	 => std_logic_vector(to_unsigned(24,8) ,
32757	 => std_logic_vector(to_unsigned(37,8) ,
32758	 => std_logic_vector(to_unsigned(10,8) ,
32759	 => std_logic_vector(to_unsigned(30,8) ,
32760	 => std_logic_vector(to_unsigned(51,8) ,
32761	 => std_logic_vector(to_unsigned(90,8) ,
32762	 => std_logic_vector(to_unsigned(50,8) ,
32763	 => std_logic_vector(to_unsigned(1,8) ,
32764	 => std_logic_vector(to_unsigned(0,8) ,
32765	 => std_logic_vector(to_unsigned(1,8) ,
32766	 => std_logic_vector(to_unsigned(6,8) ,
32767	 => std_logic_vector(to_unsigned(9,8) ,
32768	 => std_logic_vector(to_unsigned(8,8) ,
32769	 => std_logic_vector(to_unsigned(10,8) ,
32770	 => std_logic_vector(to_unsigned(48,8) ,
32771	 => std_logic_vector(to_unsigned(111,8) ,
32772	 => std_logic_vector(to_unsigned(108,8) ,
32773	 => std_logic_vector(to_unsigned(122,8) ,
32774	 => std_logic_vector(to_unsigned(142,8) ,
32775	 => std_logic_vector(to_unsigned(161,8) ,
32776	 => std_logic_vector(to_unsigned(171,8) ,
32777	 => std_logic_vector(to_unsigned(179,8) ,
32778	 => std_logic_vector(to_unsigned(181,8) ,
32779	 => std_logic_vector(to_unsigned(179,8) ,
32780	 => std_logic_vector(to_unsigned(171,8) ,
32781	 => std_logic_vector(to_unsigned(170,8) ,
32782	 => std_logic_vector(to_unsigned(164,8) ,
32783	 => std_logic_vector(to_unsigned(161,8) ,
32784	 => std_logic_vector(to_unsigned(159,8) ,
32785	 => std_logic_vector(to_unsigned(124,8) ,
32786	 => std_logic_vector(to_unsigned(103,8) ,
32787	 => std_logic_vector(to_unsigned(44,8) ,
32788	 => std_logic_vector(to_unsigned(13,8) ,
32789	 => std_logic_vector(to_unsigned(4,8) ,
32790	 => std_logic_vector(to_unsigned(3,8) ,
32791	 => std_logic_vector(to_unsigned(6,8) ,
32792	 => std_logic_vector(to_unsigned(4,8) ,
32793	 => std_logic_vector(to_unsigned(4,8) ,
32794	 => std_logic_vector(to_unsigned(1,8) ,
32795	 => std_logic_vector(to_unsigned(1,8) ,
32796	 => std_logic_vector(to_unsigned(6,8) ,
32797	 => std_logic_vector(to_unsigned(7,8) ,
32798	 => std_logic_vector(to_unsigned(11,8) ,
32799	 => std_logic_vector(to_unsigned(26,8) ,
32800	 => std_logic_vector(to_unsigned(32,8) ,
32801	 => std_logic_vector(to_unsigned(19,8) ,
32802	 => std_logic_vector(to_unsigned(11,8) ,
32803	 => std_logic_vector(to_unsigned(7,8) ,
32804	 => std_logic_vector(to_unsigned(4,8) ,
32805	 => std_logic_vector(to_unsigned(1,8) ,
32806	 => std_logic_vector(to_unsigned(10,8) ,
32807	 => std_logic_vector(to_unsigned(45,8) ,
32808	 => std_logic_vector(to_unsigned(30,8) ,
32809	 => std_logic_vector(to_unsigned(21,8) ,
32810	 => std_logic_vector(to_unsigned(12,8) ,
32811	 => std_logic_vector(to_unsigned(3,8) ,
32812	 => std_logic_vector(to_unsigned(2,8) ,
32813	 => std_logic_vector(to_unsigned(2,8) ,
32814	 => std_logic_vector(to_unsigned(0,8) ,
32815	 => std_logic_vector(to_unsigned(2,8) ,
32816	 => std_logic_vector(to_unsigned(10,8) ,
32817	 => std_logic_vector(to_unsigned(10,8) ,
32818	 => std_logic_vector(to_unsigned(8,8) ,
32819	 => std_logic_vector(to_unsigned(7,8) ,
32820	 => std_logic_vector(to_unsigned(5,8) ,
32821	 => std_logic_vector(to_unsigned(3,8) ,
32822	 => std_logic_vector(to_unsigned(4,8) ,
32823	 => std_logic_vector(to_unsigned(3,8) ,
32824	 => std_logic_vector(to_unsigned(6,8) ,
32825	 => std_logic_vector(to_unsigned(5,8) ,
32826	 => std_logic_vector(to_unsigned(3,8) ,
32827	 => std_logic_vector(to_unsigned(47,8) ,
32828	 => std_logic_vector(to_unsigned(84,8) ,
32829	 => std_logic_vector(to_unsigned(70,8) ,
32830	 => std_logic_vector(to_unsigned(69,8) ,
32831	 => std_logic_vector(to_unsigned(14,8) ,
32832	 => std_logic_vector(to_unsigned(7,8) ,
32833	 => std_logic_vector(to_unsigned(3,8) ,
32834	 => std_logic_vector(to_unsigned(12,8) ,
32835	 => std_logic_vector(to_unsigned(119,8) ,
32836	 => std_logic_vector(to_unsigned(166,8) ,
32837	 => std_logic_vector(to_unsigned(184,8) ,
32838	 => std_logic_vector(to_unsigned(112,8) ,
32839	 => std_logic_vector(to_unsigned(10,8) ,
32840	 => std_logic_vector(to_unsigned(4,8) ,
32841	 => std_logic_vector(to_unsigned(6,8) ,
32842	 => std_logic_vector(to_unsigned(6,8) ,
32843	 => std_logic_vector(to_unsigned(23,8) ,
32844	 => std_logic_vector(to_unsigned(51,8) ,
32845	 => std_logic_vector(to_unsigned(37,8) ,
32846	 => std_logic_vector(to_unsigned(32,8) ,
32847	 => std_logic_vector(to_unsigned(37,8) ,
32848	 => std_logic_vector(to_unsigned(13,8) ,
32849	 => std_logic_vector(to_unsigned(27,8) ,
32850	 => std_logic_vector(to_unsigned(142,8) ,
32851	 => std_logic_vector(to_unsigned(163,8) ,
32852	 => std_logic_vector(to_unsigned(152,8) ,
32853	 => std_logic_vector(to_unsigned(154,8) ,
32854	 => std_logic_vector(to_unsigned(159,8) ,
32855	 => std_logic_vector(to_unsigned(157,8) ,
32856	 => std_logic_vector(to_unsigned(156,8) ,
32857	 => std_logic_vector(to_unsigned(154,8) ,
32858	 => std_logic_vector(to_unsigned(156,8) ,
32859	 => std_logic_vector(to_unsigned(156,8) ,
32860	 => std_logic_vector(to_unsigned(154,8) ,
32861	 => std_logic_vector(to_unsigned(149,8) ,
32862	 => std_logic_vector(to_unsigned(152,8) ,
32863	 => std_logic_vector(to_unsigned(128,8) ,
32864	 => std_logic_vector(to_unsigned(15,8) ,
32865	 => std_logic_vector(to_unsigned(2,8) ,
32866	 => std_logic_vector(to_unsigned(2,8) ,
32867	 => std_logic_vector(to_unsigned(4,8) ,
32868	 => std_logic_vector(to_unsigned(3,8) ,
32869	 => std_logic_vector(to_unsigned(4,8) ,
32870	 => std_logic_vector(to_unsigned(3,8) ,
32871	 => std_logic_vector(to_unsigned(2,8) ,
32872	 => std_logic_vector(to_unsigned(4,8) ,
32873	 => std_logic_vector(to_unsigned(30,8) ,
32874	 => std_logic_vector(to_unsigned(95,8) ,
32875	 => std_logic_vector(to_unsigned(66,8) ,
32876	 => std_logic_vector(to_unsigned(23,8) ,
32877	 => std_logic_vector(to_unsigned(11,8) ,
32878	 => std_logic_vector(to_unsigned(17,8) ,
32879	 => std_logic_vector(to_unsigned(124,8) ,
32880	 => std_logic_vector(to_unsigned(163,8) ,
32881	 => std_logic_vector(to_unsigned(147,8) ,
32882	 => std_logic_vector(to_unsigned(149,8) ,
32883	 => std_logic_vector(to_unsigned(157,8) ,
32884	 => std_logic_vector(to_unsigned(45,8) ,
32885	 => std_logic_vector(to_unsigned(2,8) ,
32886	 => std_logic_vector(to_unsigned(16,8) ,
32887	 => std_logic_vector(to_unsigned(131,8) ,
32888	 => std_logic_vector(to_unsigned(168,8) ,
32889	 => std_logic_vector(to_unsigned(147,8) ,
32890	 => std_logic_vector(to_unsigned(156,8) ,
32891	 => std_logic_vector(to_unsigned(157,8) ,
32892	 => std_logic_vector(to_unsigned(157,8) ,
32893	 => std_logic_vector(to_unsigned(159,8) ,
32894	 => std_logic_vector(to_unsigned(156,8) ,
32895	 => std_logic_vector(to_unsigned(151,8) ,
32896	 => std_logic_vector(to_unsigned(115,8) ,
32897	 => std_logic_vector(to_unsigned(23,8) ,
32898	 => std_logic_vector(to_unsigned(0,8) ,
32899	 => std_logic_vector(to_unsigned(3,8) ,
32900	 => std_logic_vector(to_unsigned(16,8) ,
32901	 => std_logic_vector(to_unsigned(11,8) ,
32902	 => std_logic_vector(to_unsigned(7,8) ,
32903	 => std_logic_vector(to_unsigned(9,8) ,
32904	 => std_logic_vector(to_unsigned(16,8) ,
32905	 => std_logic_vector(to_unsigned(71,8) ,
32906	 => std_logic_vector(to_unsigned(177,8) ,
32907	 => std_logic_vector(to_unsigned(115,8) ,
32908	 => std_logic_vector(to_unsigned(45,8) ,
32909	 => std_logic_vector(to_unsigned(127,8) ,
32910	 => std_logic_vector(to_unsigned(166,8) ,
32911	 => std_logic_vector(to_unsigned(146,8) ,
32912	 => std_logic_vector(to_unsigned(119,8) ,
32913	 => std_logic_vector(to_unsigned(38,8) ,
32914	 => std_logic_vector(to_unsigned(1,8) ,
32915	 => std_logic_vector(to_unsigned(1,8) ,
32916	 => std_logic_vector(to_unsigned(1,8) ,
32917	 => std_logic_vector(to_unsigned(2,8) ,
32918	 => std_logic_vector(to_unsigned(5,8) ,
32919	 => std_logic_vector(to_unsigned(5,8) ,
32920	 => std_logic_vector(to_unsigned(4,8) ,
32921	 => std_logic_vector(to_unsigned(6,8) ,
32922	 => std_logic_vector(to_unsigned(6,8) ,
32923	 => std_logic_vector(to_unsigned(5,8) ,
32924	 => std_logic_vector(to_unsigned(6,8) ,
32925	 => std_logic_vector(to_unsigned(7,8) ,
32926	 => std_logic_vector(to_unsigned(5,8) ,
32927	 => std_logic_vector(to_unsigned(4,8) ,
32928	 => std_logic_vector(to_unsigned(4,8) ,
32929	 => std_logic_vector(to_unsigned(4,8) ,
32930	 => std_logic_vector(to_unsigned(2,8) ,
32931	 => std_logic_vector(to_unsigned(2,8) ,
32932	 => std_logic_vector(to_unsigned(2,8) ,
32933	 => std_logic_vector(to_unsigned(1,8) ,
32934	 => std_logic_vector(to_unsigned(1,8) ,
32935	 => std_logic_vector(to_unsigned(13,8) ,
32936	 => std_logic_vector(to_unsigned(109,8) ,
32937	 => std_logic_vector(to_unsigned(149,8) ,
32938	 => std_logic_vector(to_unsigned(154,8) ,
32939	 => std_logic_vector(to_unsigned(168,8) ,
32940	 => std_logic_vector(to_unsigned(142,8) ,
32941	 => std_logic_vector(to_unsigned(136,8) ,
32942	 => std_logic_vector(to_unsigned(161,8) ,
32943	 => std_logic_vector(to_unsigned(151,8) ,
32944	 => std_logic_vector(to_unsigned(133,8) ,
32945	 => std_logic_vector(to_unsigned(124,8) ,
32946	 => std_logic_vector(to_unsigned(128,8) ,
32947	 => std_logic_vector(to_unsigned(134,8) ,
32948	 => std_logic_vector(to_unsigned(125,8) ,
32949	 => std_logic_vector(to_unsigned(147,8) ,
32950	 => std_logic_vector(to_unsigned(163,8) ,
32951	 => std_logic_vector(to_unsigned(159,8) ,
32952	 => std_logic_vector(to_unsigned(164,8) ,
32953	 => std_logic_vector(to_unsigned(161,8) ,
32954	 => std_logic_vector(to_unsigned(164,8) ,
32955	 => std_logic_vector(to_unsigned(163,8) ,
32956	 => std_logic_vector(to_unsigned(159,8) ,
32957	 => std_logic_vector(to_unsigned(157,8) ,
32958	 => std_logic_vector(to_unsigned(156,8) ,
32959	 => std_logic_vector(to_unsigned(159,8) ,
32960	 => std_logic_vector(to_unsigned(157,8) ,
32961	 => std_logic_vector(to_unsigned(8,8) ,
32962	 => std_logic_vector(to_unsigned(6,8) ,
32963	 => std_logic_vector(to_unsigned(5,8) ,
32964	 => std_logic_vector(to_unsigned(5,8) ,
32965	 => std_logic_vector(to_unsigned(4,8) ,
32966	 => std_logic_vector(to_unsigned(2,8) ,
32967	 => std_logic_vector(to_unsigned(3,8) ,
32968	 => std_logic_vector(to_unsigned(2,8) ,
32969	 => std_logic_vector(to_unsigned(1,8) ,
32970	 => std_logic_vector(to_unsigned(1,8) ,
32971	 => std_logic_vector(to_unsigned(1,8) ,
32972	 => std_logic_vector(to_unsigned(1,8) ,
32973	 => std_logic_vector(to_unsigned(1,8) ,
32974	 => std_logic_vector(to_unsigned(1,8) ,
32975	 => std_logic_vector(to_unsigned(2,8) ,
32976	 => std_logic_vector(to_unsigned(1,8) ,
32977	 => std_logic_vector(to_unsigned(1,8) ,
32978	 => std_logic_vector(to_unsigned(3,8) ,
32979	 => std_logic_vector(to_unsigned(2,8) ,
32980	 => std_logic_vector(to_unsigned(2,8) ,
32981	 => std_logic_vector(to_unsigned(3,8) ,
32982	 => std_logic_vector(to_unsigned(2,8) ,
32983	 => std_logic_vector(to_unsigned(1,8) ,
32984	 => std_logic_vector(to_unsigned(1,8) ,
32985	 => std_logic_vector(to_unsigned(0,8) ,
32986	 => std_logic_vector(to_unsigned(2,8) ,
32987	 => std_logic_vector(to_unsigned(12,8) ,
32988	 => std_logic_vector(to_unsigned(9,8) ,
32989	 => std_logic_vector(to_unsigned(8,8) ,
32990	 => std_logic_vector(to_unsigned(7,8) ,
32991	 => std_logic_vector(to_unsigned(6,8) ,
32992	 => std_logic_vector(to_unsigned(10,8) ,
32993	 => std_logic_vector(to_unsigned(14,8) ,
32994	 => std_logic_vector(to_unsigned(6,8) ,
32995	 => std_logic_vector(to_unsigned(14,8) ,
32996	 => std_logic_vector(to_unsigned(53,8) ,
32997	 => std_logic_vector(to_unsigned(39,8) ,
32998	 => std_logic_vector(to_unsigned(35,8) ,
32999	 => std_logic_vector(to_unsigned(34,8) ,
33000	 => std_logic_vector(to_unsigned(19,8) ,
33001	 => std_logic_vector(to_unsigned(5,8) ,
33002	 => std_logic_vector(to_unsigned(4,8) ,
33003	 => std_logic_vector(to_unsigned(2,8) ,
33004	 => std_logic_vector(to_unsigned(1,8) ,
33005	 => std_logic_vector(to_unsigned(3,8) ,
33006	 => std_logic_vector(to_unsigned(13,8) ,
33007	 => std_logic_vector(to_unsigned(2,8) ,
33008	 => std_logic_vector(to_unsigned(0,8) ,
33009	 => std_logic_vector(to_unsigned(1,8) ,
33010	 => std_logic_vector(to_unsigned(0,8) ,
33011	 => std_logic_vector(to_unsigned(0,8) ,
33012	 => std_logic_vector(to_unsigned(13,8) ,
33013	 => std_logic_vector(to_unsigned(50,8) ,
33014	 => std_logic_vector(to_unsigned(41,8) ,
33015	 => std_logic_vector(to_unsigned(46,8) ,
33016	 => std_logic_vector(to_unsigned(47,8) ,
33017	 => std_logic_vector(to_unsigned(31,8) ,
33018	 => std_logic_vector(to_unsigned(13,8) ,
33019	 => std_logic_vector(to_unsigned(16,8) ,
33020	 => std_logic_vector(to_unsigned(17,8) ,
33021	 => std_logic_vector(to_unsigned(14,8) ,
33022	 => std_logic_vector(to_unsigned(13,8) ,
33023	 => std_logic_vector(to_unsigned(5,8) ,
33024	 => std_logic_vector(to_unsigned(1,8) ,
33025	 => std_logic_vector(to_unsigned(0,8) ,
33026	 => std_logic_vector(to_unsigned(0,8) ,
33027	 => std_logic_vector(to_unsigned(0,8) ,
33028	 => std_logic_vector(to_unsigned(0,8) ,
33029	 => std_logic_vector(to_unsigned(1,8) ,
33030	 => std_logic_vector(to_unsigned(2,8) ,
33031	 => std_logic_vector(to_unsigned(2,8) ,
33032	 => std_logic_vector(to_unsigned(8,8) ,
33033	 => std_logic_vector(to_unsigned(8,8) ,
33034	 => std_logic_vector(to_unsigned(5,8) ,
33035	 => std_logic_vector(to_unsigned(5,8) ,
33036	 => std_logic_vector(to_unsigned(9,8) ,
33037	 => std_logic_vector(to_unsigned(6,8) ,
33038	 => std_logic_vector(to_unsigned(9,8) ,
33039	 => std_logic_vector(to_unsigned(11,8) ,
33040	 => std_logic_vector(to_unsigned(5,8) ,
33041	 => std_logic_vector(to_unsigned(3,8) ,
33042	 => std_logic_vector(to_unsigned(1,8) ,
33043	 => std_logic_vector(to_unsigned(1,8) ,
33044	 => std_logic_vector(to_unsigned(1,8) ,
33045	 => std_logic_vector(to_unsigned(2,8) ,
33046	 => std_logic_vector(to_unsigned(3,8) ,
33047	 => std_logic_vector(to_unsigned(4,8) ,
33048	 => std_logic_vector(to_unsigned(6,8) ,
33049	 => std_logic_vector(to_unsigned(13,8) ,
33050	 => std_logic_vector(to_unsigned(6,8) ,
33051	 => std_logic_vector(to_unsigned(3,8) ,
33052	 => std_logic_vector(to_unsigned(1,8) ,
33053	 => std_logic_vector(to_unsigned(1,8) ,
33054	 => std_logic_vector(to_unsigned(3,8) ,
33055	 => std_logic_vector(to_unsigned(8,8) ,
33056	 => std_logic_vector(to_unsigned(5,8) ,
33057	 => std_logic_vector(to_unsigned(2,8) ,
33058	 => std_logic_vector(to_unsigned(3,8) ,
33059	 => std_logic_vector(to_unsigned(4,8) ,
33060	 => std_logic_vector(to_unsigned(17,8) ,
33061	 => std_logic_vector(to_unsigned(23,8) ,
33062	 => std_logic_vector(to_unsigned(17,8) ,
33063	 => std_logic_vector(to_unsigned(17,8) ,
33064	 => std_logic_vector(to_unsigned(15,8) ,
33065	 => std_logic_vector(to_unsigned(5,8) ,
33066	 => std_logic_vector(to_unsigned(13,8) ,
33067	 => std_logic_vector(to_unsigned(64,8) ,
33068	 => std_logic_vector(to_unsigned(63,8) ,
33069	 => std_logic_vector(to_unsigned(16,8) ,
33070	 => std_logic_vector(to_unsigned(8,8) ,
33071	 => std_logic_vector(to_unsigned(10,8) ,
33072	 => std_logic_vector(to_unsigned(20,8) ,
33073	 => std_logic_vector(to_unsigned(17,8) ,
33074	 => std_logic_vector(to_unsigned(31,8) ,
33075	 => std_logic_vector(to_unsigned(38,8) ,
33076	 => std_logic_vector(to_unsigned(15,8) ,
33077	 => std_logic_vector(to_unsigned(35,8) ,
33078	 => std_logic_vector(to_unsigned(23,8) ,
33079	 => std_logic_vector(to_unsigned(32,8) ,
33080	 => std_logic_vector(to_unsigned(32,8) ,
33081	 => std_logic_vector(to_unsigned(24,8) ,
33082	 => std_logic_vector(to_unsigned(26,8) ,
33083	 => std_logic_vector(to_unsigned(3,8) ,
33084	 => std_logic_vector(to_unsigned(1,8) ,
33085	 => std_logic_vector(to_unsigned(10,8) ,
33086	 => std_logic_vector(to_unsigned(17,8) ,
33087	 => std_logic_vector(to_unsigned(11,8) ,
33088	 => std_logic_vector(to_unsigned(14,8) ,
33089	 => std_logic_vector(to_unsigned(19,8) ,
33090	 => std_logic_vector(to_unsigned(31,8) ,
33091	 => std_logic_vector(to_unsigned(161,8) ,
33092	 => std_logic_vector(to_unsigned(177,8) ,
33093	 => std_logic_vector(to_unsigned(166,8) ,
33094	 => std_logic_vector(to_unsigned(159,8) ,
33095	 => std_logic_vector(to_unsigned(156,8) ,
33096	 => std_logic_vector(to_unsigned(157,8) ,
33097	 => std_logic_vector(to_unsigned(152,8) ,
33098	 => std_logic_vector(to_unsigned(146,8) ,
33099	 => std_logic_vector(to_unsigned(147,8) ,
33100	 => std_logic_vector(to_unsigned(147,8) ,
33101	 => std_logic_vector(to_unsigned(147,8) ,
33102	 => std_logic_vector(to_unsigned(151,8) ,
33103	 => std_logic_vector(to_unsigned(144,8) ,
33104	 => std_logic_vector(to_unsigned(151,8) ,
33105	 => std_logic_vector(to_unsigned(133,8) ,
33106	 => std_logic_vector(to_unsigned(80,8) ,
33107	 => std_logic_vector(to_unsigned(25,8) ,
33108	 => std_logic_vector(to_unsigned(9,8) ,
33109	 => std_logic_vector(to_unsigned(5,8) ,
33110	 => std_logic_vector(to_unsigned(3,8) ,
33111	 => std_logic_vector(to_unsigned(3,8) ,
33112	 => std_logic_vector(to_unsigned(3,8) ,
33113	 => std_logic_vector(to_unsigned(1,8) ,
33114	 => std_logic_vector(to_unsigned(2,8) ,
33115	 => std_logic_vector(to_unsigned(6,8) ,
33116	 => std_logic_vector(to_unsigned(9,8) ,
33117	 => std_logic_vector(to_unsigned(6,8) ,
33118	 => std_logic_vector(to_unsigned(8,8) ,
33119	 => std_logic_vector(to_unsigned(15,8) ,
33120	 => std_logic_vector(to_unsigned(16,8) ,
33121	 => std_logic_vector(to_unsigned(14,8) ,
33122	 => std_logic_vector(to_unsigned(11,8) ,
33123	 => std_logic_vector(to_unsigned(8,8) ,
33124	 => std_logic_vector(to_unsigned(4,8) ,
33125	 => std_logic_vector(to_unsigned(1,8) ,
33126	 => std_logic_vector(to_unsigned(1,8) ,
33127	 => std_logic_vector(to_unsigned(7,8) ,
33128	 => std_logic_vector(to_unsigned(9,8) ,
33129	 => std_logic_vector(to_unsigned(3,8) ,
33130	 => std_logic_vector(to_unsigned(1,8) ,
33131	 => std_logic_vector(to_unsigned(1,8) ,
33132	 => std_logic_vector(to_unsigned(2,8) ,
33133	 => std_logic_vector(to_unsigned(1,8) ,
33134	 => std_logic_vector(to_unsigned(2,8) ,
33135	 => std_logic_vector(to_unsigned(15,8) ,
33136	 => std_logic_vector(to_unsigned(25,8) ,
33137	 => std_logic_vector(to_unsigned(16,8) ,
33138	 => std_logic_vector(to_unsigned(9,8) ,
33139	 => std_logic_vector(to_unsigned(9,8) ,
33140	 => std_logic_vector(to_unsigned(5,8) ,
33141	 => std_logic_vector(to_unsigned(5,8) ,
33142	 => std_logic_vector(to_unsigned(4,8) ,
33143	 => std_logic_vector(to_unsigned(8,8) ,
33144	 => std_logic_vector(to_unsigned(12,8) ,
33145	 => std_logic_vector(to_unsigned(6,8) ,
33146	 => std_logic_vector(to_unsigned(11,8) ,
33147	 => std_logic_vector(to_unsigned(52,8) ,
33148	 => std_logic_vector(to_unsigned(58,8) ,
33149	 => std_logic_vector(to_unsigned(67,8) ,
33150	 => std_logic_vector(to_unsigned(34,8) ,
33151	 => std_logic_vector(to_unsigned(6,8) ,
33152	 => std_logic_vector(to_unsigned(5,8) ,
33153	 => std_logic_vector(to_unsigned(5,8) ,
33154	 => std_logic_vector(to_unsigned(7,8) ,
33155	 => std_logic_vector(to_unsigned(20,8) ,
33156	 => std_logic_vector(to_unsigned(46,8) ,
33157	 => std_logic_vector(to_unsigned(103,8) ,
33158	 => std_logic_vector(to_unsigned(40,8) ,
33159	 => std_logic_vector(to_unsigned(2,8) ,
33160	 => std_logic_vector(to_unsigned(3,8) ,
33161	 => std_logic_vector(to_unsigned(6,8) ,
33162	 => std_logic_vector(to_unsigned(8,8) ,
33163	 => std_logic_vector(to_unsigned(12,8) ,
33164	 => std_logic_vector(to_unsigned(20,8) ,
33165	 => std_logic_vector(to_unsigned(13,8) ,
33166	 => std_logic_vector(to_unsigned(24,8) ,
33167	 => std_logic_vector(to_unsigned(30,8) ,
33168	 => std_logic_vector(to_unsigned(14,8) ,
33169	 => std_logic_vector(to_unsigned(3,8) ,
33170	 => std_logic_vector(to_unsigned(60,8) ,
33171	 => std_logic_vector(to_unsigned(175,8) ,
33172	 => std_logic_vector(to_unsigned(154,8) ,
33173	 => std_logic_vector(to_unsigned(156,8) ,
33174	 => std_logic_vector(to_unsigned(156,8) ,
33175	 => std_logic_vector(to_unsigned(157,8) ,
33176	 => std_logic_vector(to_unsigned(156,8) ,
33177	 => std_logic_vector(to_unsigned(157,8) ,
33178	 => std_logic_vector(to_unsigned(157,8) ,
33179	 => std_logic_vector(to_unsigned(151,8) ,
33180	 => std_logic_vector(to_unsigned(152,8) ,
33181	 => std_logic_vector(to_unsigned(149,8) ,
33182	 => std_logic_vector(to_unsigned(149,8) ,
33183	 => std_logic_vector(to_unsigned(146,8) ,
33184	 => std_logic_vector(to_unsigned(30,8) ,
33185	 => std_logic_vector(to_unsigned(1,8) ,
33186	 => std_logic_vector(to_unsigned(2,8) ,
33187	 => std_logic_vector(to_unsigned(1,8) ,
33188	 => std_logic_vector(to_unsigned(2,8) ,
33189	 => std_logic_vector(to_unsigned(3,8) ,
33190	 => std_logic_vector(to_unsigned(2,8) ,
33191	 => std_logic_vector(to_unsigned(3,8) ,
33192	 => std_logic_vector(to_unsigned(3,8) ,
33193	 => std_logic_vector(to_unsigned(5,8) ,
33194	 => std_logic_vector(to_unsigned(35,8) ,
33195	 => std_logic_vector(to_unsigned(74,8) ,
33196	 => std_logic_vector(to_unsigned(25,8) ,
33197	 => std_logic_vector(to_unsigned(0,8) ,
33198	 => std_logic_vector(to_unsigned(7,8) ,
33199	 => std_logic_vector(to_unsigned(131,8) ,
33200	 => std_logic_vector(to_unsigned(156,8) ,
33201	 => std_logic_vector(to_unsigned(146,8) ,
33202	 => std_logic_vector(to_unsigned(151,8) ,
33203	 => std_logic_vector(to_unsigned(159,8) ,
33204	 => std_logic_vector(to_unsigned(45,8) ,
33205	 => std_logic_vector(to_unsigned(2,8) ,
33206	 => std_logic_vector(to_unsigned(18,8) ,
33207	 => std_logic_vector(to_unsigned(136,8) ,
33208	 => std_logic_vector(to_unsigned(161,8) ,
33209	 => std_logic_vector(to_unsigned(149,8) ,
33210	 => std_logic_vector(to_unsigned(159,8) ,
33211	 => std_logic_vector(to_unsigned(161,8) ,
33212	 => std_logic_vector(to_unsigned(161,8) ,
33213	 => std_logic_vector(to_unsigned(157,8) ,
33214	 => std_logic_vector(to_unsigned(157,8) ,
33215	 => std_logic_vector(to_unsigned(154,8) ,
33216	 => std_logic_vector(to_unsigned(208,8) ,
33217	 => std_logic_vector(to_unsigned(96,8) ,
33218	 => std_logic_vector(to_unsigned(2,8) ,
33219	 => std_logic_vector(to_unsigned(1,8) ,
33220	 => std_logic_vector(to_unsigned(9,8) ,
33221	 => std_logic_vector(to_unsigned(13,8) ,
33222	 => std_logic_vector(to_unsigned(8,8) ,
33223	 => std_logic_vector(to_unsigned(14,8) ,
33224	 => std_logic_vector(to_unsigned(12,8) ,
33225	 => std_logic_vector(to_unsigned(41,8) ,
33226	 => std_logic_vector(to_unsigned(163,8) ,
33227	 => std_logic_vector(to_unsigned(108,8) ,
33228	 => std_logic_vector(to_unsigned(57,8) ,
33229	 => std_logic_vector(to_unsigned(146,8) ,
33230	 => std_logic_vector(to_unsigned(164,8) ,
33231	 => std_logic_vector(to_unsigned(157,8) ,
33232	 => std_logic_vector(to_unsigned(115,8) ,
33233	 => std_logic_vector(to_unsigned(33,8) ,
33234	 => std_logic_vector(to_unsigned(2,8) ,
33235	 => std_logic_vector(to_unsigned(1,8) ,
33236	 => std_logic_vector(to_unsigned(2,8) ,
33237	 => std_logic_vector(to_unsigned(1,8) ,
33238	 => std_logic_vector(to_unsigned(2,8) ,
33239	 => std_logic_vector(to_unsigned(4,8) ,
33240	 => std_logic_vector(to_unsigned(4,8) ,
33241	 => std_logic_vector(to_unsigned(4,8) ,
33242	 => std_logic_vector(to_unsigned(6,8) ,
33243	 => std_logic_vector(to_unsigned(5,8) ,
33244	 => std_logic_vector(to_unsigned(5,8) ,
33245	 => std_logic_vector(to_unsigned(5,8) ,
33246	 => std_logic_vector(to_unsigned(5,8) ,
33247	 => std_logic_vector(to_unsigned(4,8) ,
33248	 => std_logic_vector(to_unsigned(2,8) ,
33249	 => std_logic_vector(to_unsigned(1,8) ,
33250	 => std_logic_vector(to_unsigned(1,8) ,
33251	 => std_logic_vector(to_unsigned(1,8) ,
33252	 => std_logic_vector(to_unsigned(1,8) ,
33253	 => std_logic_vector(to_unsigned(1,8) ,
33254	 => std_logic_vector(to_unsigned(2,8) ,
33255	 => std_logic_vector(to_unsigned(13,8) ,
33256	 => std_logic_vector(to_unsigned(62,8) ,
33257	 => std_logic_vector(to_unsigned(101,8) ,
33258	 => std_logic_vector(to_unsigned(144,8) ,
33259	 => std_logic_vector(to_unsigned(156,8) ,
33260	 => std_logic_vector(to_unsigned(128,8) ,
33261	 => std_logic_vector(to_unsigned(119,8) ,
33262	 => std_logic_vector(to_unsigned(164,8) ,
33263	 => std_logic_vector(to_unsigned(152,8) ,
33264	 => std_logic_vector(to_unsigned(142,8) ,
33265	 => std_logic_vector(to_unsigned(147,8) ,
33266	 => std_logic_vector(to_unsigned(127,8) ,
33267	 => std_logic_vector(to_unsigned(116,8) ,
33268	 => std_logic_vector(to_unsigned(121,8) ,
33269	 => std_logic_vector(to_unsigned(139,8) ,
33270	 => std_logic_vector(to_unsigned(151,8) ,
33271	 => std_logic_vector(to_unsigned(151,8) ,
33272	 => std_logic_vector(to_unsigned(156,8) ,
33273	 => std_logic_vector(to_unsigned(152,8) ,
33274	 => std_logic_vector(to_unsigned(154,8) ,
33275	 => std_logic_vector(to_unsigned(156,8) ,
33276	 => std_logic_vector(to_unsigned(159,8) ,
33277	 => std_logic_vector(to_unsigned(152,8) ,
33278	 => std_logic_vector(to_unsigned(159,8) ,
33279	 => std_logic_vector(to_unsigned(159,8) ,
33280	 => std_logic_vector(to_unsigned(149,8) ,
33281	 => std_logic_vector(to_unsigned(5,8) ,
33282	 => std_logic_vector(to_unsigned(5,8) ,
33283	 => std_logic_vector(to_unsigned(6,8) ,
33284	 => std_logic_vector(to_unsigned(5,8) ,
33285	 => std_logic_vector(to_unsigned(5,8) ,
33286	 => std_logic_vector(to_unsigned(4,8) ,
33287	 => std_logic_vector(to_unsigned(2,8) ,
33288	 => std_logic_vector(to_unsigned(3,8) ,
33289	 => std_logic_vector(to_unsigned(1,8) ,
33290	 => std_logic_vector(to_unsigned(1,8) ,
33291	 => std_logic_vector(to_unsigned(2,8) ,
33292	 => std_logic_vector(to_unsigned(2,8) ,
33293	 => std_logic_vector(to_unsigned(1,8) ,
33294	 => std_logic_vector(to_unsigned(1,8) ,
33295	 => std_logic_vector(to_unsigned(2,8) ,
33296	 => std_logic_vector(to_unsigned(1,8) ,
33297	 => std_logic_vector(to_unsigned(1,8) ,
33298	 => std_logic_vector(to_unsigned(1,8) ,
33299	 => std_logic_vector(to_unsigned(1,8) ,
33300	 => std_logic_vector(to_unsigned(3,8) ,
33301	 => std_logic_vector(to_unsigned(1,8) ,
33302	 => std_logic_vector(to_unsigned(1,8) ,
33303	 => std_logic_vector(to_unsigned(0,8) ,
33304	 => std_logic_vector(to_unsigned(0,8) ,
33305	 => std_logic_vector(to_unsigned(0,8) ,
33306	 => std_logic_vector(to_unsigned(0,8) ,
33307	 => std_logic_vector(to_unsigned(9,8) ,
33308	 => std_logic_vector(to_unsigned(17,8) ,
33309	 => std_logic_vector(to_unsigned(12,8) ,
33310	 => std_logic_vector(to_unsigned(8,8) ,
33311	 => std_logic_vector(to_unsigned(13,8) ,
33312	 => std_logic_vector(to_unsigned(19,8) ,
33313	 => std_logic_vector(to_unsigned(22,8) ,
33314	 => std_logic_vector(to_unsigned(17,8) ,
33315	 => std_logic_vector(to_unsigned(40,8) ,
33316	 => std_logic_vector(to_unsigned(45,8) ,
33317	 => std_logic_vector(to_unsigned(28,8) ,
33318	 => std_logic_vector(to_unsigned(34,8) ,
33319	 => std_logic_vector(to_unsigned(24,8) ,
33320	 => std_logic_vector(to_unsigned(10,8) ,
33321	 => std_logic_vector(to_unsigned(6,8) ,
33322	 => std_logic_vector(to_unsigned(4,8) ,
33323	 => std_logic_vector(to_unsigned(1,8) ,
33324	 => std_logic_vector(to_unsigned(1,8) ,
33325	 => std_logic_vector(to_unsigned(12,8) ,
33326	 => std_logic_vector(to_unsigned(14,8) ,
33327	 => std_logic_vector(to_unsigned(2,8) ,
33328	 => std_logic_vector(to_unsigned(0,8) ,
33329	 => std_logic_vector(to_unsigned(0,8) ,
33330	 => std_logic_vector(to_unsigned(1,8) ,
33331	 => std_logic_vector(to_unsigned(1,8) ,
33332	 => std_logic_vector(to_unsigned(2,8) ,
33333	 => std_logic_vector(to_unsigned(16,8) ,
33334	 => std_logic_vector(to_unsigned(22,8) ,
33335	 => std_logic_vector(to_unsigned(25,8) ,
33336	 => std_logic_vector(to_unsigned(24,8) ,
33337	 => std_logic_vector(to_unsigned(16,8) ,
33338	 => std_logic_vector(to_unsigned(6,8) ,
33339	 => std_logic_vector(to_unsigned(3,8) ,
33340	 => std_logic_vector(to_unsigned(7,8) ,
33341	 => std_logic_vector(to_unsigned(12,8) ,
33342	 => std_logic_vector(to_unsigned(17,8) ,
33343	 => std_logic_vector(to_unsigned(17,8) ,
33344	 => std_logic_vector(to_unsigned(8,8) ,
33345	 => std_logic_vector(to_unsigned(2,8) ,
33346	 => std_logic_vector(to_unsigned(0,8) ,
33347	 => std_logic_vector(to_unsigned(1,8) ,
33348	 => std_logic_vector(to_unsigned(1,8) ,
33349	 => std_logic_vector(to_unsigned(0,8) ,
33350	 => std_logic_vector(to_unsigned(1,8) ,
33351	 => std_logic_vector(to_unsigned(2,8) ,
33352	 => std_logic_vector(to_unsigned(4,8) ,
33353	 => std_logic_vector(to_unsigned(3,8) ,
33354	 => std_logic_vector(to_unsigned(4,8) ,
33355	 => std_logic_vector(to_unsigned(7,8) ,
33356	 => std_logic_vector(to_unsigned(10,8) ,
33357	 => std_logic_vector(to_unsigned(2,8) ,
33358	 => std_logic_vector(to_unsigned(5,8) ,
33359	 => std_logic_vector(to_unsigned(8,8) ,
33360	 => std_logic_vector(to_unsigned(8,8) ,
33361	 => std_logic_vector(to_unsigned(4,8) ,
33362	 => std_logic_vector(to_unsigned(1,8) ,
33363	 => std_logic_vector(to_unsigned(2,8) ,
33364	 => std_logic_vector(to_unsigned(2,8) ,
33365	 => std_logic_vector(to_unsigned(0,8) ,
33366	 => std_logic_vector(to_unsigned(0,8) ,
33367	 => std_logic_vector(to_unsigned(0,8) ,
33368	 => std_logic_vector(to_unsigned(0,8) ,
33369	 => std_logic_vector(to_unsigned(0,8) ,
33370	 => std_logic_vector(to_unsigned(2,8) ,
33371	 => std_logic_vector(to_unsigned(2,8) ,
33372	 => std_logic_vector(to_unsigned(2,8) ,
33373	 => std_logic_vector(to_unsigned(5,8) ,
33374	 => std_logic_vector(to_unsigned(8,8) ,
33375	 => std_logic_vector(to_unsigned(8,8) ,
33376	 => std_logic_vector(to_unsigned(5,8) ,
33377	 => std_logic_vector(to_unsigned(3,8) ,
33378	 => std_logic_vector(to_unsigned(1,8) ,
33379	 => std_logic_vector(to_unsigned(6,8) ,
33380	 => std_logic_vector(to_unsigned(19,8) ,
33381	 => std_logic_vector(to_unsigned(14,8) ,
33382	 => std_logic_vector(to_unsigned(16,8) ,
33383	 => std_logic_vector(to_unsigned(12,8) ,
33384	 => std_logic_vector(to_unsigned(8,8) ,
33385	 => std_logic_vector(to_unsigned(2,8) ,
33386	 => std_logic_vector(to_unsigned(9,8) ,
33387	 => std_logic_vector(to_unsigned(51,8) ,
33388	 => std_logic_vector(to_unsigned(45,8) ,
33389	 => std_logic_vector(to_unsigned(7,8) ,
33390	 => std_logic_vector(to_unsigned(4,8) ,
33391	 => std_logic_vector(to_unsigned(8,8) ,
33392	 => std_logic_vector(to_unsigned(15,8) ,
33393	 => std_logic_vector(to_unsigned(30,8) ,
33394	 => std_logic_vector(to_unsigned(29,8) ,
33395	 => std_logic_vector(to_unsigned(42,8) ,
33396	 => std_logic_vector(to_unsigned(10,8) ,
33397	 => std_logic_vector(to_unsigned(19,8) ,
33398	 => std_logic_vector(to_unsigned(24,8) ,
33399	 => std_logic_vector(to_unsigned(25,8) ,
33400	 => std_logic_vector(to_unsigned(27,8) ,
33401	 => std_logic_vector(to_unsigned(13,8) ,
33402	 => std_logic_vector(to_unsigned(15,8) ,
33403	 => std_logic_vector(to_unsigned(3,8) ,
33404	 => std_logic_vector(to_unsigned(2,8) ,
33405	 => std_logic_vector(to_unsigned(12,8) ,
33406	 => std_logic_vector(to_unsigned(15,8) ,
33407	 => std_logic_vector(to_unsigned(10,8) ,
33408	 => std_logic_vector(to_unsigned(9,8) ,
33409	 => std_logic_vector(to_unsigned(19,8) ,
33410	 => std_logic_vector(to_unsigned(23,8) ,
33411	 => std_logic_vector(to_unsigned(125,8) ,
33412	 => std_logic_vector(to_unsigned(161,8) ,
33413	 => std_logic_vector(to_unsigned(149,8) ,
33414	 => std_logic_vector(to_unsigned(152,8) ,
33415	 => std_logic_vector(to_unsigned(149,8) ,
33416	 => std_logic_vector(to_unsigned(149,8) ,
33417	 => std_logic_vector(to_unsigned(147,8) ,
33418	 => std_logic_vector(to_unsigned(151,8) ,
33419	 => std_logic_vector(to_unsigned(147,8) ,
33420	 => std_logic_vector(to_unsigned(149,8) ,
33421	 => std_logic_vector(to_unsigned(149,8) ,
33422	 => std_logic_vector(to_unsigned(152,8) ,
33423	 => std_logic_vector(to_unsigned(146,8) ,
33424	 => std_logic_vector(to_unsigned(144,8) ,
33425	 => std_logic_vector(to_unsigned(149,8) ,
33426	 => std_logic_vector(to_unsigned(49,8) ,
33427	 => std_logic_vector(to_unsigned(6,8) ,
33428	 => std_logic_vector(to_unsigned(4,8) ,
33429	 => std_logic_vector(to_unsigned(5,8) ,
33430	 => std_logic_vector(to_unsigned(4,8) ,
33431	 => std_logic_vector(to_unsigned(3,8) ,
33432	 => std_logic_vector(to_unsigned(2,8) ,
33433	 => std_logic_vector(to_unsigned(1,8) ,
33434	 => std_logic_vector(to_unsigned(3,8) ,
33435	 => std_logic_vector(to_unsigned(6,8) ,
33436	 => std_logic_vector(to_unsigned(8,8) ,
33437	 => std_logic_vector(to_unsigned(3,8) ,
33438	 => std_logic_vector(to_unsigned(5,8) ,
33439	 => std_logic_vector(to_unsigned(10,8) ,
33440	 => std_logic_vector(to_unsigned(14,8) ,
33441	 => std_logic_vector(to_unsigned(10,8) ,
33442	 => std_logic_vector(to_unsigned(6,8) ,
33443	 => std_logic_vector(to_unsigned(6,8) ,
33444	 => std_logic_vector(to_unsigned(3,8) ,
33445	 => std_logic_vector(to_unsigned(1,8) ,
33446	 => std_logic_vector(to_unsigned(1,8) ,
33447	 => std_logic_vector(to_unsigned(1,8) ,
33448	 => std_logic_vector(to_unsigned(0,8) ,
33449	 => std_logic_vector(to_unsigned(0,8) ,
33450	 => std_logic_vector(to_unsigned(1,8) ,
33451	 => std_logic_vector(to_unsigned(0,8) ,
33452	 => std_logic_vector(to_unsigned(1,8) ,
33453	 => std_logic_vector(to_unsigned(1,8) ,
33454	 => std_logic_vector(to_unsigned(4,8) ,
33455	 => std_logic_vector(to_unsigned(17,8) ,
33456	 => std_logic_vector(to_unsigned(22,8) ,
33457	 => std_logic_vector(to_unsigned(13,8) ,
33458	 => std_logic_vector(to_unsigned(8,8) ,
33459	 => std_logic_vector(to_unsigned(6,8) ,
33460	 => std_logic_vector(to_unsigned(4,8) ,
33461	 => std_logic_vector(to_unsigned(3,8) ,
33462	 => std_logic_vector(to_unsigned(6,8) ,
33463	 => std_logic_vector(to_unsigned(10,8) ,
33464	 => std_logic_vector(to_unsigned(8,8) ,
33465	 => std_logic_vector(to_unsigned(6,8) ,
33466	 => std_logic_vector(to_unsigned(15,8) ,
33467	 => std_logic_vector(to_unsigned(44,8) ,
33468	 => std_logic_vector(to_unsigned(38,8) ,
33469	 => std_logic_vector(to_unsigned(29,8) ,
33470	 => std_logic_vector(to_unsigned(12,8) ,
33471	 => std_logic_vector(to_unsigned(4,8) ,
33472	 => std_logic_vector(to_unsigned(4,8) ,
33473	 => std_logic_vector(to_unsigned(3,8) ,
33474	 => std_logic_vector(to_unsigned(4,8) ,
33475	 => std_logic_vector(to_unsigned(2,8) ,
33476	 => std_logic_vector(to_unsigned(2,8) ,
33477	 => std_logic_vector(to_unsigned(7,8) ,
33478	 => std_logic_vector(to_unsigned(11,8) ,
33479	 => std_logic_vector(to_unsigned(3,8) ,
33480	 => std_logic_vector(to_unsigned(4,8) ,
33481	 => std_logic_vector(to_unsigned(9,8) ,
33482	 => std_logic_vector(to_unsigned(5,8) ,
33483	 => std_logic_vector(to_unsigned(12,8) ,
33484	 => std_logic_vector(to_unsigned(28,8) ,
33485	 => std_logic_vector(to_unsigned(17,8) ,
33486	 => std_logic_vector(to_unsigned(17,8) ,
33487	 => std_logic_vector(to_unsigned(16,8) ,
33488	 => std_logic_vector(to_unsigned(8,8) ,
33489	 => std_logic_vector(to_unsigned(3,8) ,
33490	 => std_logic_vector(to_unsigned(78,8) ,
33491	 => std_logic_vector(to_unsigned(175,8) ,
33492	 => std_logic_vector(to_unsigned(154,8) ,
33493	 => std_logic_vector(to_unsigned(156,8) ,
33494	 => std_logic_vector(to_unsigned(156,8) ,
33495	 => std_logic_vector(to_unsigned(156,8) ,
33496	 => std_logic_vector(to_unsigned(157,8) ,
33497	 => std_logic_vector(to_unsigned(159,8) ,
33498	 => std_logic_vector(to_unsigned(157,8) ,
33499	 => std_logic_vector(to_unsigned(156,8) ,
33500	 => std_logic_vector(to_unsigned(146,8) ,
33501	 => std_logic_vector(to_unsigned(144,8) ,
33502	 => std_logic_vector(to_unsigned(147,8) ,
33503	 => std_logic_vector(to_unsigned(157,8) ,
33504	 => std_logic_vector(to_unsigned(84,8) ,
33505	 => std_logic_vector(to_unsigned(2,8) ,
33506	 => std_logic_vector(to_unsigned(2,8) ,
33507	 => std_logic_vector(to_unsigned(4,8) ,
33508	 => std_logic_vector(to_unsigned(2,8) ,
33509	 => std_logic_vector(to_unsigned(2,8) ,
33510	 => std_logic_vector(to_unsigned(2,8) ,
33511	 => std_logic_vector(to_unsigned(1,8) ,
33512	 => std_logic_vector(to_unsigned(2,8) ,
33513	 => std_logic_vector(to_unsigned(10,8) ,
33514	 => std_logic_vector(to_unsigned(30,8) ,
33515	 => std_logic_vector(to_unsigned(40,8) ,
33516	 => std_logic_vector(to_unsigned(18,8) ,
33517	 => std_logic_vector(to_unsigned(5,8) ,
33518	 => std_logic_vector(to_unsigned(9,8) ,
33519	 => std_logic_vector(to_unsigned(111,8) ,
33520	 => std_logic_vector(to_unsigned(159,8) ,
33521	 => std_logic_vector(to_unsigned(144,8) ,
33522	 => std_logic_vector(to_unsigned(152,8) ,
33523	 => std_logic_vector(to_unsigned(154,8) ,
33524	 => std_logic_vector(to_unsigned(30,8) ,
33525	 => std_logic_vector(to_unsigned(1,8) ,
33526	 => std_logic_vector(to_unsigned(19,8) ,
33527	 => std_logic_vector(to_unsigned(138,8) ,
33528	 => std_logic_vector(to_unsigned(159,8) ,
33529	 => std_logic_vector(to_unsigned(151,8) ,
33530	 => std_logic_vector(to_unsigned(156,8) ,
33531	 => std_logic_vector(to_unsigned(159,8) ,
33532	 => std_logic_vector(to_unsigned(157,8) ,
33533	 => std_logic_vector(to_unsigned(159,8) ,
33534	 => std_logic_vector(to_unsigned(161,8) ,
33535	 => std_logic_vector(to_unsigned(164,8) ,
33536	 => std_logic_vector(to_unsigned(101,8) ,
33537	 => std_logic_vector(to_unsigned(27,8) ,
33538	 => std_logic_vector(to_unsigned(12,8) ,
33539	 => std_logic_vector(to_unsigned(1,8) ,
33540	 => std_logic_vector(to_unsigned(2,8) ,
33541	 => std_logic_vector(to_unsigned(15,8) ,
33542	 => std_logic_vector(to_unsigned(11,8) ,
33543	 => std_logic_vector(to_unsigned(9,8) ,
33544	 => std_logic_vector(to_unsigned(11,8) ,
33545	 => std_logic_vector(to_unsigned(26,8) ,
33546	 => std_logic_vector(to_unsigned(128,8) ,
33547	 => std_logic_vector(to_unsigned(108,8) ,
33548	 => std_logic_vector(to_unsigned(51,8) ,
33549	 => std_logic_vector(to_unsigned(141,8) ,
33550	 => std_logic_vector(to_unsigned(166,8) ,
33551	 => std_logic_vector(to_unsigned(142,8) ,
33552	 => std_logic_vector(to_unsigned(101,8) ,
33553	 => std_logic_vector(to_unsigned(25,8) ,
33554	 => std_logic_vector(to_unsigned(4,8) ,
33555	 => std_logic_vector(to_unsigned(7,8) ,
33556	 => std_logic_vector(to_unsigned(4,8) ,
33557	 => std_logic_vector(to_unsigned(1,8) ,
33558	 => std_logic_vector(to_unsigned(1,8) ,
33559	 => std_logic_vector(to_unsigned(4,8) ,
33560	 => std_logic_vector(to_unsigned(4,8) ,
33561	 => std_logic_vector(to_unsigned(4,8) ,
33562	 => std_logic_vector(to_unsigned(6,8) ,
33563	 => std_logic_vector(to_unsigned(7,8) ,
33564	 => std_logic_vector(to_unsigned(6,8) ,
33565	 => std_logic_vector(to_unsigned(7,8) ,
33566	 => std_logic_vector(to_unsigned(7,8) ,
33567	 => std_logic_vector(to_unsigned(6,8) ,
33568	 => std_logic_vector(to_unsigned(2,8) ,
33569	 => std_logic_vector(to_unsigned(2,8) ,
33570	 => std_logic_vector(to_unsigned(1,8) ,
33571	 => std_logic_vector(to_unsigned(6,8) ,
33572	 => std_logic_vector(to_unsigned(30,8) ,
33573	 => std_logic_vector(to_unsigned(7,8) ,
33574	 => std_logic_vector(to_unsigned(1,8) ,
33575	 => std_logic_vector(to_unsigned(31,8) ,
33576	 => std_logic_vector(to_unsigned(92,8) ,
33577	 => std_logic_vector(to_unsigned(130,8) ,
33578	 => std_logic_vector(to_unsigned(156,8) ,
33579	 => std_logic_vector(to_unsigned(127,8) ,
33580	 => std_logic_vector(to_unsigned(88,8) ,
33581	 => std_logic_vector(to_unsigned(131,8) ,
33582	 => std_logic_vector(to_unsigned(166,8) ,
33583	 => std_logic_vector(to_unsigned(142,8) ,
33584	 => std_logic_vector(to_unsigned(138,8) ,
33585	 => std_logic_vector(to_unsigned(142,8) ,
33586	 => std_logic_vector(to_unsigned(28,8) ,
33587	 => std_logic_vector(to_unsigned(23,8) ,
33588	 => std_logic_vector(to_unsigned(125,8) ,
33589	 => std_logic_vector(to_unsigned(139,8) ,
33590	 => std_logic_vector(to_unsigned(130,8) ,
33591	 => std_logic_vector(to_unsigned(128,8) ,
33592	 => std_logic_vector(to_unsigned(133,8) ,
33593	 => std_logic_vector(to_unsigned(142,8) ,
33594	 => std_logic_vector(to_unsigned(149,8) ,
33595	 => std_logic_vector(to_unsigned(154,8) ,
33596	 => std_logic_vector(to_unsigned(152,8) ,
33597	 => std_logic_vector(to_unsigned(154,8) ,
33598	 => std_logic_vector(to_unsigned(149,8) ,
33599	 => std_logic_vector(to_unsigned(147,8) ,
33600	 => std_logic_vector(to_unsigned(151,8) ,
33601	 => std_logic_vector(to_unsigned(4,8) ,
33602	 => std_logic_vector(to_unsigned(4,8) ,
33603	 => std_logic_vector(to_unsigned(4,8) ,
33604	 => std_logic_vector(to_unsigned(4,8) ,
33605	 => std_logic_vector(to_unsigned(4,8) ,
33606	 => std_logic_vector(to_unsigned(5,8) ,
33607	 => std_logic_vector(to_unsigned(2,8) ,
33608	 => std_logic_vector(to_unsigned(2,8) ,
33609	 => std_logic_vector(to_unsigned(2,8) ,
33610	 => std_logic_vector(to_unsigned(2,8) ,
33611	 => std_logic_vector(to_unsigned(1,8) ,
33612	 => std_logic_vector(to_unsigned(2,8) ,
33613	 => std_logic_vector(to_unsigned(2,8) ,
33614	 => std_logic_vector(to_unsigned(1,8) ,
33615	 => std_logic_vector(to_unsigned(0,8) ,
33616	 => std_logic_vector(to_unsigned(1,8) ,
33617	 => std_logic_vector(to_unsigned(1,8) ,
33618	 => std_logic_vector(to_unsigned(0,8) ,
33619	 => std_logic_vector(to_unsigned(3,8) ,
33620	 => std_logic_vector(to_unsigned(3,8) ,
33621	 => std_logic_vector(to_unsigned(1,8) ,
33622	 => std_logic_vector(to_unsigned(1,8) ,
33623	 => std_logic_vector(to_unsigned(0,8) ,
33624	 => std_logic_vector(to_unsigned(0,8) ,
33625	 => std_logic_vector(to_unsigned(0,8) ,
33626	 => std_logic_vector(to_unsigned(0,8) ,
33627	 => std_logic_vector(to_unsigned(4,8) ,
33628	 => std_logic_vector(to_unsigned(16,8) ,
33629	 => std_logic_vector(to_unsigned(12,8) ,
33630	 => std_logic_vector(to_unsigned(9,8) ,
33631	 => std_logic_vector(to_unsigned(13,8) ,
33632	 => std_logic_vector(to_unsigned(8,8) ,
33633	 => std_logic_vector(to_unsigned(3,8) ,
33634	 => std_logic_vector(to_unsigned(15,8) ,
33635	 => std_logic_vector(to_unsigned(39,8) ,
33636	 => std_logic_vector(to_unsigned(28,8) ,
33637	 => std_logic_vector(to_unsigned(28,8) ,
33638	 => std_logic_vector(to_unsigned(30,8) ,
33639	 => std_logic_vector(to_unsigned(11,8) ,
33640	 => std_logic_vector(to_unsigned(4,8) ,
33641	 => std_logic_vector(to_unsigned(4,8) ,
33642	 => std_logic_vector(to_unsigned(5,8) ,
33643	 => std_logic_vector(to_unsigned(3,8) ,
33644	 => std_logic_vector(to_unsigned(7,8) ,
33645	 => std_logic_vector(to_unsigned(22,8) ,
33646	 => std_logic_vector(to_unsigned(9,8) ,
33647	 => std_logic_vector(to_unsigned(1,8) ,
33648	 => std_logic_vector(to_unsigned(0,8) ,
33649	 => std_logic_vector(to_unsigned(0,8) ,
33650	 => std_logic_vector(to_unsigned(1,8) ,
33651	 => std_logic_vector(to_unsigned(1,8) ,
33652	 => std_logic_vector(to_unsigned(2,8) ,
33653	 => std_logic_vector(to_unsigned(8,8) ,
33654	 => std_logic_vector(to_unsigned(9,8) ,
33655	 => std_logic_vector(to_unsigned(20,8) ,
33656	 => std_logic_vector(to_unsigned(13,8) ,
33657	 => std_logic_vector(to_unsigned(13,8) ,
33658	 => std_logic_vector(to_unsigned(10,8) ,
33659	 => std_logic_vector(to_unsigned(4,8) ,
33660	 => std_logic_vector(to_unsigned(1,8) ,
33661	 => std_logic_vector(to_unsigned(6,8) ,
33662	 => std_logic_vector(to_unsigned(12,8) ,
33663	 => std_logic_vector(to_unsigned(8,8) ,
33664	 => std_logic_vector(to_unsigned(10,8) ,
33665	 => std_logic_vector(to_unsigned(3,8) ,
33666	 => std_logic_vector(to_unsigned(1,8) ,
33667	 => std_logic_vector(to_unsigned(1,8) ,
33668	 => std_logic_vector(to_unsigned(0,8) ,
33669	 => std_logic_vector(to_unsigned(1,8) ,
33670	 => std_logic_vector(to_unsigned(1,8) ,
33671	 => std_logic_vector(to_unsigned(4,8) ,
33672	 => std_logic_vector(to_unsigned(3,8) ,
33673	 => std_logic_vector(to_unsigned(2,8) ,
33674	 => std_logic_vector(to_unsigned(6,8) ,
33675	 => std_logic_vector(to_unsigned(8,8) ,
33676	 => std_logic_vector(to_unsigned(7,8) ,
33677	 => std_logic_vector(to_unsigned(1,8) ,
33678	 => std_logic_vector(to_unsigned(7,8) ,
33679	 => std_logic_vector(to_unsigned(8,8) ,
33680	 => std_logic_vector(to_unsigned(6,8) ,
33681	 => std_logic_vector(to_unsigned(4,8) ,
33682	 => std_logic_vector(to_unsigned(2,8) ,
33683	 => std_logic_vector(to_unsigned(1,8) ,
33684	 => std_logic_vector(to_unsigned(1,8) ,
33685	 => std_logic_vector(to_unsigned(1,8) ,
33686	 => std_logic_vector(to_unsigned(0,8) ,
33687	 => std_logic_vector(to_unsigned(0,8) ,
33688	 => std_logic_vector(to_unsigned(0,8) ,
33689	 => std_logic_vector(to_unsigned(0,8) ,
33690	 => std_logic_vector(to_unsigned(0,8) ,
33691	 => std_logic_vector(to_unsigned(1,8) ,
33692	 => std_logic_vector(to_unsigned(4,8) ,
33693	 => std_logic_vector(to_unsigned(9,8) ,
33694	 => std_logic_vector(to_unsigned(8,8) ,
33695	 => std_logic_vector(to_unsigned(8,8) ,
33696	 => std_logic_vector(to_unsigned(8,8) ,
33697	 => std_logic_vector(to_unsigned(7,8) ,
33698	 => std_logic_vector(to_unsigned(1,8) ,
33699	 => std_logic_vector(to_unsigned(4,8) ,
33700	 => std_logic_vector(to_unsigned(18,8) ,
33701	 => std_logic_vector(to_unsigned(11,8) ,
33702	 => std_logic_vector(to_unsigned(10,8) ,
33703	 => std_logic_vector(to_unsigned(8,8) ,
33704	 => std_logic_vector(to_unsigned(4,8) ,
33705	 => std_logic_vector(to_unsigned(1,8) ,
33706	 => std_logic_vector(to_unsigned(7,8) ,
33707	 => std_logic_vector(to_unsigned(44,8) ,
33708	 => std_logic_vector(to_unsigned(19,8) ,
33709	 => std_logic_vector(to_unsigned(2,8) ,
33710	 => std_logic_vector(to_unsigned(6,8) ,
33711	 => std_logic_vector(to_unsigned(6,8) ,
33712	 => std_logic_vector(to_unsigned(9,8) ,
33713	 => std_logic_vector(to_unsigned(17,8) ,
33714	 => std_logic_vector(to_unsigned(15,8) ,
33715	 => std_logic_vector(to_unsigned(7,8) ,
33716	 => std_logic_vector(to_unsigned(2,8) ,
33717	 => std_logic_vector(to_unsigned(5,8) ,
33718	 => std_logic_vector(to_unsigned(9,8) ,
33719	 => std_logic_vector(to_unsigned(19,8) ,
33720	 => std_logic_vector(to_unsigned(15,8) ,
33721	 => std_logic_vector(to_unsigned(9,8) ,
33722	 => std_logic_vector(to_unsigned(5,8) ,
33723	 => std_logic_vector(to_unsigned(3,8) ,
33724	 => std_logic_vector(to_unsigned(6,8) ,
33725	 => std_logic_vector(to_unsigned(13,8) ,
33726	 => std_logic_vector(to_unsigned(14,8) ,
33727	 => std_logic_vector(to_unsigned(17,8) ,
33728	 => std_logic_vector(to_unsigned(8,8) ,
33729	 => std_logic_vector(to_unsigned(9,8) ,
33730	 => std_logic_vector(to_unsigned(37,8) ,
33731	 => std_logic_vector(to_unsigned(125,8) ,
33732	 => std_logic_vector(to_unsigned(152,8) ,
33733	 => std_logic_vector(to_unsigned(147,8) ,
33734	 => std_logic_vector(to_unsigned(152,8) ,
33735	 => std_logic_vector(to_unsigned(147,8) ,
33736	 => std_logic_vector(to_unsigned(149,8) ,
33737	 => std_logic_vector(to_unsigned(156,8) ,
33738	 => std_logic_vector(to_unsigned(157,8) ,
33739	 => std_logic_vector(to_unsigned(163,8) ,
33740	 => std_logic_vector(to_unsigned(164,8) ,
33741	 => std_logic_vector(to_unsigned(170,8) ,
33742	 => std_logic_vector(to_unsigned(170,8) ,
33743	 => std_logic_vector(to_unsigned(163,8) ,
33744	 => std_logic_vector(to_unsigned(154,8) ,
33745	 => std_logic_vector(to_unsigned(149,8) ,
33746	 => std_logic_vector(to_unsigned(27,8) ,
33747	 => std_logic_vector(to_unsigned(2,8) ,
33748	 => std_logic_vector(to_unsigned(6,8) ,
33749	 => std_logic_vector(to_unsigned(6,8) ,
33750	 => std_logic_vector(to_unsigned(4,8) ,
33751	 => std_logic_vector(to_unsigned(1,8) ,
33752	 => std_logic_vector(to_unsigned(1,8) ,
33753	 => std_logic_vector(to_unsigned(2,8) ,
33754	 => std_logic_vector(to_unsigned(4,8) ,
33755	 => std_logic_vector(to_unsigned(7,8) ,
33756	 => std_logic_vector(to_unsigned(7,8) ,
33757	 => std_logic_vector(to_unsigned(2,8) ,
33758	 => std_logic_vector(to_unsigned(4,8) ,
33759	 => std_logic_vector(to_unsigned(10,8) ,
33760	 => std_logic_vector(to_unsigned(12,8) ,
33761	 => std_logic_vector(to_unsigned(8,8) ,
33762	 => std_logic_vector(to_unsigned(4,8) ,
33763	 => std_logic_vector(to_unsigned(3,8) ,
33764	 => std_logic_vector(to_unsigned(3,8) ,
33765	 => std_logic_vector(to_unsigned(3,8) ,
33766	 => std_logic_vector(to_unsigned(1,8) ,
33767	 => std_logic_vector(to_unsigned(1,8) ,
33768	 => std_logic_vector(to_unsigned(1,8) ,
33769	 => std_logic_vector(to_unsigned(0,8) ,
33770	 => std_logic_vector(to_unsigned(0,8) ,
33771	 => std_logic_vector(to_unsigned(1,8) ,
33772	 => std_logic_vector(to_unsigned(1,8) ,
33773	 => std_logic_vector(to_unsigned(1,8) ,
33774	 => std_logic_vector(to_unsigned(3,8) ,
33775	 => std_logic_vector(to_unsigned(9,8) ,
33776	 => std_logic_vector(to_unsigned(12,8) ,
33777	 => std_logic_vector(to_unsigned(9,8) ,
33778	 => std_logic_vector(to_unsigned(7,8) ,
33779	 => std_logic_vector(to_unsigned(8,8) ,
33780	 => std_logic_vector(to_unsigned(4,8) ,
33781	 => std_logic_vector(to_unsigned(3,8) ,
33782	 => std_logic_vector(to_unsigned(8,8) ,
33783	 => std_logic_vector(to_unsigned(7,8) ,
33784	 => std_logic_vector(to_unsigned(6,8) ,
33785	 => std_logic_vector(to_unsigned(5,8) ,
33786	 => std_logic_vector(to_unsigned(10,8) ,
33787	 => std_logic_vector(to_unsigned(23,8) ,
33788	 => std_logic_vector(to_unsigned(17,8) ,
33789	 => std_logic_vector(to_unsigned(9,8) ,
33790	 => std_logic_vector(to_unsigned(5,8) ,
33791	 => std_logic_vector(to_unsigned(2,8) ,
33792	 => std_logic_vector(to_unsigned(4,8) ,
33793	 => std_logic_vector(to_unsigned(3,8) ,
33794	 => std_logic_vector(to_unsigned(2,8) ,
33795	 => std_logic_vector(to_unsigned(2,8) ,
33796	 => std_logic_vector(to_unsigned(5,8) ,
33797	 => std_logic_vector(to_unsigned(7,8) ,
33798	 => std_logic_vector(to_unsigned(6,8) ,
33799	 => std_logic_vector(to_unsigned(7,8) ,
33800	 => std_logic_vector(to_unsigned(5,8) ,
33801	 => std_logic_vector(to_unsigned(3,8) ,
33802	 => std_logic_vector(to_unsigned(2,8) ,
33803	 => std_logic_vector(to_unsigned(5,8) ,
33804	 => std_logic_vector(to_unsigned(17,8) ,
33805	 => std_logic_vector(to_unsigned(12,8) ,
33806	 => std_logic_vector(to_unsigned(4,8) ,
33807	 => std_logic_vector(to_unsigned(6,8) ,
33808	 => std_logic_vector(to_unsigned(2,8) ,
33809	 => std_logic_vector(to_unsigned(13,8) ,
33810	 => std_logic_vector(to_unsigned(144,8) ,
33811	 => std_logic_vector(to_unsigned(166,8) ,
33812	 => std_logic_vector(to_unsigned(151,8) ,
33813	 => std_logic_vector(to_unsigned(157,8) ,
33814	 => std_logic_vector(to_unsigned(159,8) ,
33815	 => std_logic_vector(to_unsigned(156,8) ,
33816	 => std_logic_vector(to_unsigned(152,8) ,
33817	 => std_logic_vector(to_unsigned(152,8) ,
33818	 => std_logic_vector(to_unsigned(154,8) ,
33819	 => std_logic_vector(to_unsigned(159,8) ,
33820	 => std_logic_vector(to_unsigned(146,8) ,
33821	 => std_logic_vector(to_unsigned(146,8) ,
33822	 => std_logic_vector(to_unsigned(154,8) ,
33823	 => std_logic_vector(to_unsigned(147,8) ,
33824	 => std_logic_vector(to_unsigned(144,8) ,
33825	 => std_logic_vector(to_unsigned(35,8) ,
33826	 => std_logic_vector(to_unsigned(1,8) ,
33827	 => std_logic_vector(to_unsigned(2,8) ,
33828	 => std_logic_vector(to_unsigned(2,8) ,
33829	 => std_logic_vector(to_unsigned(3,8) ,
33830	 => std_logic_vector(to_unsigned(3,8) ,
33831	 => std_logic_vector(to_unsigned(1,8) ,
33832	 => std_logic_vector(to_unsigned(3,8) ,
33833	 => std_logic_vector(to_unsigned(10,8) ,
33834	 => std_logic_vector(to_unsigned(18,8) ,
33835	 => std_logic_vector(to_unsigned(17,8) ,
33836	 => std_logic_vector(to_unsigned(12,8) ,
33837	 => std_logic_vector(to_unsigned(14,8) ,
33838	 => std_logic_vector(to_unsigned(8,8) ,
33839	 => std_logic_vector(to_unsigned(30,8) ,
33840	 => std_logic_vector(to_unsigned(142,8) ,
33841	 => std_logic_vector(to_unsigned(157,8) ,
33842	 => std_logic_vector(to_unsigned(142,8) ,
33843	 => std_logic_vector(to_unsigned(149,8) ,
33844	 => std_logic_vector(to_unsigned(26,8) ,
33845	 => std_logic_vector(to_unsigned(2,8) ,
33846	 => std_logic_vector(to_unsigned(21,8) ,
33847	 => std_logic_vector(to_unsigned(142,8) ,
33848	 => std_logic_vector(to_unsigned(163,8) ,
33849	 => std_logic_vector(to_unsigned(149,8) ,
33850	 => std_logic_vector(to_unsigned(157,8) ,
33851	 => std_logic_vector(to_unsigned(159,8) ,
33852	 => std_logic_vector(to_unsigned(157,8) ,
33853	 => std_logic_vector(to_unsigned(157,8) ,
33854	 => std_logic_vector(to_unsigned(149,8) ,
33855	 => std_logic_vector(to_unsigned(175,8) ,
33856	 => std_logic_vector(to_unsigned(36,8) ,
33857	 => std_logic_vector(to_unsigned(1,8) ,
33858	 => std_logic_vector(to_unsigned(8,8) ,
33859	 => std_logic_vector(to_unsigned(8,8) ,
33860	 => std_logic_vector(to_unsigned(5,8) ,
33861	 => std_logic_vector(to_unsigned(13,8) ,
33862	 => std_logic_vector(to_unsigned(14,8) ,
33863	 => std_logic_vector(to_unsigned(7,8) ,
33864	 => std_logic_vector(to_unsigned(12,8) ,
33865	 => std_logic_vector(to_unsigned(21,8) ,
33866	 => std_logic_vector(to_unsigned(95,8) ,
33867	 => std_logic_vector(to_unsigned(74,8) ,
33868	 => std_logic_vector(to_unsigned(49,8) ,
33869	 => std_logic_vector(to_unsigned(139,8) ,
33870	 => std_logic_vector(to_unsigned(151,8) ,
33871	 => std_logic_vector(to_unsigned(128,8) ,
33872	 => std_logic_vector(to_unsigned(70,8) ,
33873	 => std_logic_vector(to_unsigned(12,8) ,
33874	 => std_logic_vector(to_unsigned(3,8) ,
33875	 => std_logic_vector(to_unsigned(9,8) ,
33876	 => std_logic_vector(to_unsigned(7,8) ,
33877	 => std_logic_vector(to_unsigned(3,8) ,
33878	 => std_logic_vector(to_unsigned(2,8) ,
33879	 => std_logic_vector(to_unsigned(3,8) ,
33880	 => std_logic_vector(to_unsigned(4,8) ,
33881	 => std_logic_vector(to_unsigned(4,8) ,
33882	 => std_logic_vector(to_unsigned(4,8) ,
33883	 => std_logic_vector(to_unsigned(5,8) ,
33884	 => std_logic_vector(to_unsigned(6,8) ,
33885	 => std_logic_vector(to_unsigned(9,8) ,
33886	 => std_logic_vector(to_unsigned(7,8) ,
33887	 => std_logic_vector(to_unsigned(4,8) ,
33888	 => std_logic_vector(to_unsigned(2,8) ,
33889	 => std_logic_vector(to_unsigned(2,8) ,
33890	 => std_logic_vector(to_unsigned(1,8) ,
33891	 => std_logic_vector(to_unsigned(29,8) ,
33892	 => std_logic_vector(to_unsigned(118,8) ,
33893	 => std_logic_vector(to_unsigned(19,8) ,
33894	 => std_logic_vector(to_unsigned(2,8) ,
33895	 => std_logic_vector(to_unsigned(65,8) ,
33896	 => std_logic_vector(to_unsigned(138,8) ,
33897	 => std_logic_vector(to_unsigned(152,8) ,
33898	 => std_logic_vector(to_unsigned(141,8) ,
33899	 => std_logic_vector(to_unsigned(116,8) ,
33900	 => std_logic_vector(to_unsigned(90,8) ,
33901	 => std_logic_vector(to_unsigned(115,8) ,
33902	 => std_logic_vector(to_unsigned(147,8) ,
33903	 => std_logic_vector(to_unsigned(128,8) ,
33904	 => std_logic_vector(to_unsigned(130,8) ,
33905	 => std_logic_vector(to_unsigned(101,8) ,
33906	 => std_logic_vector(to_unsigned(3,8) ,
33907	 => std_logic_vector(to_unsigned(7,8) ,
33908	 => std_logic_vector(to_unsigned(109,8) ,
33909	 => std_logic_vector(to_unsigned(138,8) ,
33910	 => std_logic_vector(to_unsigned(124,8) ,
33911	 => std_logic_vector(to_unsigned(128,8) ,
33912	 => std_logic_vector(to_unsigned(127,8) ,
33913	 => std_logic_vector(to_unsigned(133,8) ,
33914	 => std_logic_vector(to_unsigned(146,8) ,
33915	 => std_logic_vector(to_unsigned(146,8) ,
33916	 => std_logic_vector(to_unsigned(124,8) ,
33917	 => std_logic_vector(to_unsigned(125,8) ,
33918	 => std_logic_vector(to_unsigned(122,8) ,
33919	 => std_logic_vector(to_unsigned(130,8) ,
33920	 => std_logic_vector(to_unsigned(136,8) ,
33921	 => std_logic_vector(to_unsigned(6,8) ,
33922	 => std_logic_vector(to_unsigned(4,8) ,
33923	 => std_logic_vector(to_unsigned(4,8) ,
33924	 => std_logic_vector(to_unsigned(5,8) ,
33925	 => std_logic_vector(to_unsigned(4,8) ,
33926	 => std_logic_vector(to_unsigned(5,8) ,
33927	 => std_logic_vector(to_unsigned(4,8) ,
33928	 => std_logic_vector(to_unsigned(2,8) ,
33929	 => std_logic_vector(to_unsigned(2,8) ,
33930	 => std_logic_vector(to_unsigned(2,8) ,
33931	 => std_logic_vector(to_unsigned(1,8) ,
33932	 => std_logic_vector(to_unsigned(1,8) ,
33933	 => std_logic_vector(to_unsigned(2,8) ,
33934	 => std_logic_vector(to_unsigned(1,8) ,
33935	 => std_logic_vector(to_unsigned(0,8) ,
33936	 => std_logic_vector(to_unsigned(1,8) ,
33937	 => std_logic_vector(to_unsigned(3,8) ,
33938	 => std_logic_vector(to_unsigned(2,8) ,
33939	 => std_logic_vector(to_unsigned(3,8) ,
33940	 => std_logic_vector(to_unsigned(1,8) ,
33941	 => std_logic_vector(to_unsigned(0,8) ,
33942	 => std_logic_vector(to_unsigned(0,8) ,
33943	 => std_logic_vector(to_unsigned(0,8) ,
33944	 => std_logic_vector(to_unsigned(0,8) ,
33945	 => std_logic_vector(to_unsigned(0,8) ,
33946	 => std_logic_vector(to_unsigned(0,8) ,
33947	 => std_logic_vector(to_unsigned(1,8) ,
33948	 => std_logic_vector(to_unsigned(11,8) ,
33949	 => std_logic_vector(to_unsigned(15,8) ,
33950	 => std_logic_vector(to_unsigned(12,8) ,
33951	 => std_logic_vector(to_unsigned(12,8) ,
33952	 => std_logic_vector(to_unsigned(6,8) ,
33953	 => std_logic_vector(to_unsigned(5,8) ,
33954	 => std_logic_vector(to_unsigned(17,8) ,
33955	 => std_logic_vector(to_unsigned(31,8) ,
33956	 => std_logic_vector(to_unsigned(35,8) ,
33957	 => std_logic_vector(to_unsigned(37,8) ,
33958	 => std_logic_vector(to_unsigned(31,8) ,
33959	 => std_logic_vector(to_unsigned(8,8) ,
33960	 => std_logic_vector(to_unsigned(6,8) ,
33961	 => std_logic_vector(to_unsigned(5,8) ,
33962	 => std_logic_vector(to_unsigned(3,8) ,
33963	 => std_logic_vector(to_unsigned(6,8) ,
33964	 => std_logic_vector(to_unsigned(17,8) ,
33965	 => std_logic_vector(to_unsigned(14,8) ,
33966	 => std_logic_vector(to_unsigned(4,8) ,
33967	 => std_logic_vector(to_unsigned(0,8) ,
33968	 => std_logic_vector(to_unsigned(0,8) ,
33969	 => std_logic_vector(to_unsigned(0,8) ,
33970	 => std_logic_vector(to_unsigned(0,8) ,
33971	 => std_logic_vector(to_unsigned(0,8) ,
33972	 => std_logic_vector(to_unsigned(12,8) ,
33973	 => std_logic_vector(to_unsigned(16,8) ,
33974	 => std_logic_vector(to_unsigned(6,8) ,
33975	 => std_logic_vector(to_unsigned(20,8) ,
33976	 => std_logic_vector(to_unsigned(10,8) ,
33977	 => std_logic_vector(to_unsigned(7,8) ,
33978	 => std_logic_vector(to_unsigned(8,8) ,
33979	 => std_logic_vector(to_unsigned(7,8) ,
33980	 => std_logic_vector(to_unsigned(5,8) ,
33981	 => std_logic_vector(to_unsigned(2,8) ,
33982	 => std_logic_vector(to_unsigned(3,8) ,
33983	 => std_logic_vector(to_unsigned(8,8) ,
33984	 => std_logic_vector(to_unsigned(9,8) ,
33985	 => std_logic_vector(to_unsigned(1,8) ,
33986	 => std_logic_vector(to_unsigned(1,8) ,
33987	 => std_logic_vector(to_unsigned(1,8) ,
33988	 => std_logic_vector(to_unsigned(0,8) ,
33989	 => std_logic_vector(to_unsigned(1,8) ,
33990	 => std_logic_vector(to_unsigned(3,8) ,
33991	 => std_logic_vector(to_unsigned(3,8) ,
33992	 => std_logic_vector(to_unsigned(2,8) ,
33993	 => std_logic_vector(to_unsigned(3,8) ,
33994	 => std_logic_vector(to_unsigned(6,8) ,
33995	 => std_logic_vector(to_unsigned(12,8) ,
33996	 => std_logic_vector(to_unsigned(5,8) ,
33997	 => std_logic_vector(to_unsigned(1,8) ,
33998	 => std_logic_vector(to_unsigned(7,8) ,
33999	 => std_logic_vector(to_unsigned(8,8) ,
34000	 => std_logic_vector(to_unsigned(7,8) ,
34001	 => std_logic_vector(to_unsigned(4,8) ,
34002	 => std_logic_vector(to_unsigned(1,8) ,
34003	 => std_logic_vector(to_unsigned(1,8) ,
34004	 => std_logic_vector(to_unsigned(1,8) ,
34005	 => std_logic_vector(to_unsigned(0,8) ,
34006	 => std_logic_vector(to_unsigned(0,8) ,
34007	 => std_logic_vector(to_unsigned(0,8) ,
34008	 => std_logic_vector(to_unsigned(0,8) ,
34009	 => std_logic_vector(to_unsigned(0,8) ,
34010	 => std_logic_vector(to_unsigned(0,8) ,
34011	 => std_logic_vector(to_unsigned(3,8) ,
34012	 => std_logic_vector(to_unsigned(8,8) ,
34013	 => std_logic_vector(to_unsigned(9,8) ,
34014	 => std_logic_vector(to_unsigned(8,8) ,
34015	 => std_logic_vector(to_unsigned(8,8) ,
34016	 => std_logic_vector(to_unsigned(6,8) ,
34017	 => std_logic_vector(to_unsigned(5,8) ,
34018	 => std_logic_vector(to_unsigned(3,8) ,
34019	 => std_logic_vector(to_unsigned(6,8) ,
34020	 => std_logic_vector(to_unsigned(15,8) ,
34021	 => std_logic_vector(to_unsigned(13,8) ,
34022	 => std_logic_vector(to_unsigned(10,8) ,
34023	 => std_logic_vector(to_unsigned(7,8) ,
34024	 => std_logic_vector(to_unsigned(6,8) ,
34025	 => std_logic_vector(to_unsigned(2,8) ,
34026	 => std_logic_vector(to_unsigned(7,8) ,
34027	 => std_logic_vector(to_unsigned(71,8) ,
34028	 => std_logic_vector(to_unsigned(28,8) ,
34029	 => std_logic_vector(to_unsigned(3,8) ,
34030	 => std_logic_vector(to_unsigned(4,8) ,
34031	 => std_logic_vector(to_unsigned(6,8) ,
34032	 => std_logic_vector(to_unsigned(5,8) ,
34033	 => std_logic_vector(to_unsigned(6,8) ,
34034	 => std_logic_vector(to_unsigned(7,8) ,
34035	 => std_logic_vector(to_unsigned(2,8) ,
34036	 => std_logic_vector(to_unsigned(1,8) ,
34037	 => std_logic_vector(to_unsigned(1,8) ,
34038	 => std_logic_vector(to_unsigned(1,8) ,
34039	 => std_logic_vector(to_unsigned(3,8) ,
34040	 => std_logic_vector(to_unsigned(3,8) ,
34041	 => std_logic_vector(to_unsigned(2,8) ,
34042	 => std_logic_vector(to_unsigned(1,8) ,
34043	 => std_logic_vector(to_unsigned(1,8) ,
34044	 => std_logic_vector(to_unsigned(7,8) ,
34045	 => std_logic_vector(to_unsigned(13,8) ,
34046	 => std_logic_vector(to_unsigned(12,8) ,
34047	 => std_logic_vector(to_unsigned(15,8) ,
34048	 => std_logic_vector(to_unsigned(11,8) ,
34049	 => std_logic_vector(to_unsigned(3,8) ,
34050	 => std_logic_vector(to_unsigned(15,8) ,
34051	 => std_logic_vector(to_unsigned(134,8) ,
34052	 => std_logic_vector(to_unsigned(181,8) ,
34053	 => std_logic_vector(to_unsigned(163,8) ,
34054	 => std_logic_vector(to_unsigned(161,8) ,
34055	 => std_logic_vector(to_unsigned(149,8) ,
34056	 => std_logic_vector(to_unsigned(141,8) ,
34057	 => std_logic_vector(to_unsigned(141,8) ,
34058	 => std_logic_vector(to_unsigned(112,8) ,
34059	 => std_logic_vector(to_unsigned(96,8) ,
34060	 => std_logic_vector(to_unsigned(78,8) ,
34061	 => std_logic_vector(to_unsigned(61,8) ,
34062	 => std_logic_vector(to_unsigned(46,8) ,
34063	 => std_logic_vector(to_unsigned(36,8) ,
34064	 => std_logic_vector(to_unsigned(27,8) ,
34065	 => std_logic_vector(to_unsigned(19,8) ,
34066	 => std_logic_vector(to_unsigned(6,8) ,
34067	 => std_logic_vector(to_unsigned(5,8) ,
34068	 => std_logic_vector(to_unsigned(7,8) ,
34069	 => std_logic_vector(to_unsigned(4,8) ,
34070	 => std_logic_vector(to_unsigned(2,8) ,
34071	 => std_logic_vector(to_unsigned(1,8) ,
34072	 => std_logic_vector(to_unsigned(2,8) ,
34073	 => std_logic_vector(to_unsigned(2,8) ,
34074	 => std_logic_vector(to_unsigned(4,8) ,
34075	 => std_logic_vector(to_unsigned(9,8) ,
34076	 => std_logic_vector(to_unsigned(8,8) ,
34077	 => std_logic_vector(to_unsigned(2,8) ,
34078	 => std_logic_vector(to_unsigned(5,8) ,
34079	 => std_logic_vector(to_unsigned(10,8) ,
34080	 => std_logic_vector(to_unsigned(10,8) ,
34081	 => std_logic_vector(to_unsigned(6,8) ,
34082	 => std_logic_vector(to_unsigned(5,8) ,
34083	 => std_logic_vector(to_unsigned(3,8) ,
34084	 => std_logic_vector(to_unsigned(2,8) ,
34085	 => std_logic_vector(to_unsigned(5,8) ,
34086	 => std_logic_vector(to_unsigned(2,8) ,
34087	 => std_logic_vector(to_unsigned(0,8) ,
34088	 => std_logic_vector(to_unsigned(1,8) ,
34089	 => std_logic_vector(to_unsigned(1,8) ,
34090	 => std_logic_vector(to_unsigned(0,8) ,
34091	 => std_logic_vector(to_unsigned(0,8) ,
34092	 => std_logic_vector(to_unsigned(0,8) ,
34093	 => std_logic_vector(to_unsigned(0,8) ,
34094	 => std_logic_vector(to_unsigned(3,8) ,
34095	 => std_logic_vector(to_unsigned(7,8) ,
34096	 => std_logic_vector(to_unsigned(8,8) ,
34097	 => std_logic_vector(to_unsigned(9,8) ,
34098	 => std_logic_vector(to_unsigned(7,8) ,
34099	 => std_logic_vector(to_unsigned(7,8) ,
34100	 => std_logic_vector(to_unsigned(5,8) ,
34101	 => std_logic_vector(to_unsigned(2,8) ,
34102	 => std_logic_vector(to_unsigned(5,8) ,
34103	 => std_logic_vector(to_unsigned(4,8) ,
34104	 => std_logic_vector(to_unsigned(5,8) ,
34105	 => std_logic_vector(to_unsigned(2,8) ,
34106	 => std_logic_vector(to_unsigned(6,8) ,
34107	 => std_logic_vector(to_unsigned(15,8) ,
34108	 => std_logic_vector(to_unsigned(12,8) ,
34109	 => std_logic_vector(to_unsigned(9,8) ,
34110	 => std_logic_vector(to_unsigned(8,8) ,
34111	 => std_logic_vector(to_unsigned(3,8) ,
34112	 => std_logic_vector(to_unsigned(2,8) ,
34113	 => std_logic_vector(to_unsigned(2,8) ,
34114	 => std_logic_vector(to_unsigned(2,8) ,
34115	 => std_logic_vector(to_unsigned(6,8) ,
34116	 => std_logic_vector(to_unsigned(7,8) ,
34117	 => std_logic_vector(to_unsigned(3,8) ,
34118	 => std_logic_vector(to_unsigned(2,8) ,
34119	 => std_logic_vector(to_unsigned(2,8) ,
34120	 => std_logic_vector(to_unsigned(1,8) ,
34121	 => std_logic_vector(to_unsigned(1,8) ,
34122	 => std_logic_vector(to_unsigned(2,8) ,
34123	 => std_logic_vector(to_unsigned(3,8) ,
34124	 => std_logic_vector(to_unsigned(2,8) ,
34125	 => std_logic_vector(to_unsigned(1,8) ,
34126	 => std_logic_vector(to_unsigned(1,8) ,
34127	 => std_logic_vector(to_unsigned(2,8) ,
34128	 => std_logic_vector(to_unsigned(1,8) ,
34129	 => std_logic_vector(to_unsigned(49,8) ,
34130	 => std_logic_vector(to_unsigned(186,8) ,
34131	 => std_logic_vector(to_unsigned(152,8) ,
34132	 => std_logic_vector(to_unsigned(147,8) ,
34133	 => std_logic_vector(to_unsigned(156,8) ,
34134	 => std_logic_vector(to_unsigned(157,8) ,
34135	 => std_logic_vector(to_unsigned(154,8) ,
34136	 => std_logic_vector(to_unsigned(151,8) ,
34137	 => std_logic_vector(to_unsigned(149,8) ,
34138	 => std_logic_vector(to_unsigned(152,8) ,
34139	 => std_logic_vector(to_unsigned(154,8) ,
34140	 => std_logic_vector(to_unsigned(151,8) ,
34141	 => std_logic_vector(to_unsigned(149,8) ,
34142	 => std_logic_vector(to_unsigned(151,8) ,
34143	 => std_logic_vector(to_unsigned(149,8) ,
34144	 => std_logic_vector(to_unsigned(144,8) ,
34145	 => std_logic_vector(to_unsigned(131,8) ,
34146	 => std_logic_vector(to_unsigned(38,8) ,
34147	 => std_logic_vector(to_unsigned(2,8) ,
34148	 => std_logic_vector(to_unsigned(1,8) ,
34149	 => std_logic_vector(to_unsigned(1,8) ,
34150	 => std_logic_vector(to_unsigned(1,8) ,
34151	 => std_logic_vector(to_unsigned(1,8) ,
34152	 => std_logic_vector(to_unsigned(2,8) ,
34153	 => std_logic_vector(to_unsigned(3,8) ,
34154	 => std_logic_vector(to_unsigned(4,8) ,
34155	 => std_logic_vector(to_unsigned(6,8) ,
34156	 => std_logic_vector(to_unsigned(6,8) ,
34157	 => std_logic_vector(to_unsigned(9,8) ,
34158	 => std_logic_vector(to_unsigned(9,8) ,
34159	 => std_logic_vector(to_unsigned(8,8) ,
34160	 => std_logic_vector(to_unsigned(66,8) ,
34161	 => std_logic_vector(to_unsigned(157,8) ,
34162	 => std_logic_vector(to_unsigned(149,8) ,
34163	 => std_logic_vector(to_unsigned(151,8) ,
34164	 => std_logic_vector(to_unsigned(30,8) ,
34165	 => std_logic_vector(to_unsigned(2,8) ,
34166	 => std_logic_vector(to_unsigned(19,8) ,
34167	 => std_logic_vector(to_unsigned(136,8) ,
34168	 => std_logic_vector(to_unsigned(159,8) ,
34169	 => std_logic_vector(to_unsigned(152,8) ,
34170	 => std_logic_vector(to_unsigned(157,8) ,
34171	 => std_logic_vector(to_unsigned(156,8) ,
34172	 => std_logic_vector(to_unsigned(156,8) ,
34173	 => std_logic_vector(to_unsigned(164,8) ,
34174	 => std_logic_vector(to_unsigned(170,8) ,
34175	 => std_logic_vector(to_unsigned(154,8) ,
34176	 => std_logic_vector(to_unsigned(53,8) ,
34177	 => std_logic_vector(to_unsigned(4,8) ,
34178	 => std_logic_vector(to_unsigned(6,8) ,
34179	 => std_logic_vector(to_unsigned(17,8) ,
34180	 => std_logic_vector(to_unsigned(25,8) ,
34181	 => std_logic_vector(to_unsigned(23,8) ,
34182	 => std_logic_vector(to_unsigned(10,8) ,
34183	 => std_logic_vector(to_unsigned(6,8) ,
34184	 => std_logic_vector(to_unsigned(8,8) ,
34185	 => std_logic_vector(to_unsigned(18,8) ,
34186	 => std_logic_vector(to_unsigned(54,8) ,
34187	 => std_logic_vector(to_unsigned(20,8) ,
34188	 => std_logic_vector(to_unsigned(32,8) ,
34189	 => std_logic_vector(to_unsigned(124,8) ,
34190	 => std_logic_vector(to_unsigned(127,8) ,
34191	 => std_logic_vector(to_unsigned(130,8) ,
34192	 => std_logic_vector(to_unsigned(42,8) ,
34193	 => std_logic_vector(to_unsigned(5,8) ,
34194	 => std_logic_vector(to_unsigned(7,8) ,
34195	 => std_logic_vector(to_unsigned(13,8) ,
34196	 => std_logic_vector(to_unsigned(13,8) ,
34197	 => std_logic_vector(to_unsigned(7,8) ,
34198	 => std_logic_vector(to_unsigned(2,8) ,
34199	 => std_logic_vector(to_unsigned(1,8) ,
34200	 => std_logic_vector(to_unsigned(1,8) ,
34201	 => std_logic_vector(to_unsigned(1,8) ,
34202	 => std_logic_vector(to_unsigned(1,8) ,
34203	 => std_logic_vector(to_unsigned(1,8) ,
34204	 => std_logic_vector(to_unsigned(1,8) ,
34205	 => std_logic_vector(to_unsigned(5,8) ,
34206	 => std_logic_vector(to_unsigned(6,8) ,
34207	 => std_logic_vector(to_unsigned(3,8) ,
34208	 => std_logic_vector(to_unsigned(2,8) ,
34209	 => std_logic_vector(to_unsigned(1,8) ,
34210	 => std_logic_vector(to_unsigned(1,8) ,
34211	 => std_logic_vector(to_unsigned(35,8) ,
34212	 => std_logic_vector(to_unsigned(124,8) ,
34213	 => std_logic_vector(to_unsigned(13,8) ,
34214	 => std_logic_vector(to_unsigned(1,8) ,
34215	 => std_logic_vector(to_unsigned(80,8) ,
34216	 => std_logic_vector(to_unsigned(157,8) ,
34217	 => std_logic_vector(to_unsigned(152,8) ,
34218	 => std_logic_vector(to_unsigned(144,8) ,
34219	 => std_logic_vector(to_unsigned(128,8) ,
34220	 => std_logic_vector(to_unsigned(121,8) ,
34221	 => std_logic_vector(to_unsigned(90,8) ,
34222	 => std_logic_vector(to_unsigned(127,8) ,
34223	 => std_logic_vector(to_unsigned(141,8) ,
34224	 => std_logic_vector(to_unsigned(125,8) ,
34225	 => std_logic_vector(to_unsigned(95,8) ,
34226	 => std_logic_vector(to_unsigned(50,8) ,
34227	 => std_logic_vector(to_unsigned(51,8) ,
34228	 => std_logic_vector(to_unsigned(107,8) ,
34229	 => std_logic_vector(to_unsigned(127,8) ,
34230	 => std_logic_vector(to_unsigned(124,8) ,
34231	 => std_logic_vector(to_unsigned(138,8) ,
34232	 => std_logic_vector(to_unsigned(138,8) ,
34233	 => std_logic_vector(to_unsigned(95,8) ,
34234	 => std_logic_vector(to_unsigned(99,8) ,
34235	 => std_logic_vector(to_unsigned(128,8) ,
34236	 => std_logic_vector(to_unsigned(108,8) ,
34237	 => std_logic_vector(to_unsigned(103,8) ,
34238	 => std_logic_vector(to_unsigned(119,8) ,
34239	 => std_logic_vector(to_unsigned(122,8) ,
34240	 => std_logic_vector(to_unsigned(115,8) ,
34241	 => std_logic_vector(to_unsigned(10,8) ,
34242	 => std_logic_vector(to_unsigned(6,8) ,
34243	 => std_logic_vector(to_unsigned(5,8) ,
34244	 => std_logic_vector(to_unsigned(6,8) ,
34245	 => std_logic_vector(to_unsigned(5,8) ,
34246	 => std_logic_vector(to_unsigned(6,8) ,
34247	 => std_logic_vector(to_unsigned(5,8) ,
34248	 => std_logic_vector(to_unsigned(3,8) ,
34249	 => std_logic_vector(to_unsigned(2,8) ,
34250	 => std_logic_vector(to_unsigned(2,8) ,
34251	 => std_logic_vector(to_unsigned(2,8) ,
34252	 => std_logic_vector(to_unsigned(1,8) ,
34253	 => std_logic_vector(to_unsigned(1,8) ,
34254	 => std_logic_vector(to_unsigned(1,8) ,
34255	 => std_logic_vector(to_unsigned(0,8) ,
34256	 => std_logic_vector(to_unsigned(0,8) ,
34257	 => std_logic_vector(to_unsigned(2,8) ,
34258	 => std_logic_vector(to_unsigned(3,8) ,
34259	 => std_logic_vector(to_unsigned(3,8) ,
34260	 => std_logic_vector(to_unsigned(1,8) ,
34261	 => std_logic_vector(to_unsigned(0,8) ,
34262	 => std_logic_vector(to_unsigned(0,8) ,
34263	 => std_logic_vector(to_unsigned(0,8) ,
34264	 => std_logic_vector(to_unsigned(0,8) ,
34265	 => std_logic_vector(to_unsigned(0,8) ,
34266	 => std_logic_vector(to_unsigned(0,8) ,
34267	 => std_logic_vector(to_unsigned(0,8) ,
34268	 => std_logic_vector(to_unsigned(6,8) ,
34269	 => std_logic_vector(to_unsigned(16,8) ,
34270	 => std_logic_vector(to_unsigned(10,8) ,
34271	 => std_logic_vector(to_unsigned(13,8) ,
34272	 => std_logic_vector(to_unsigned(10,8) ,
34273	 => std_logic_vector(to_unsigned(13,8) ,
34274	 => std_logic_vector(to_unsigned(31,8) ,
34275	 => std_logic_vector(to_unsigned(39,8) ,
34276	 => std_logic_vector(to_unsigned(40,8) ,
34277	 => std_logic_vector(to_unsigned(33,8) ,
34278	 => std_logic_vector(to_unsigned(22,8) ,
34279	 => std_logic_vector(to_unsigned(6,8) ,
34280	 => std_logic_vector(to_unsigned(12,8) ,
34281	 => std_logic_vector(to_unsigned(23,8) ,
34282	 => std_logic_vector(to_unsigned(12,8) ,
34283	 => std_logic_vector(to_unsigned(23,8) ,
34284	 => std_logic_vector(to_unsigned(19,8) ,
34285	 => std_logic_vector(to_unsigned(6,8) ,
34286	 => std_logic_vector(to_unsigned(2,8) ,
34287	 => std_logic_vector(to_unsigned(0,8) ,
34288	 => std_logic_vector(to_unsigned(0,8) ,
34289	 => std_logic_vector(to_unsigned(0,8) ,
34290	 => std_logic_vector(to_unsigned(1,8) ,
34291	 => std_logic_vector(to_unsigned(0,8) ,
34292	 => std_logic_vector(to_unsigned(10,8) ,
34293	 => std_logic_vector(to_unsigned(8,8) ,
34294	 => std_logic_vector(to_unsigned(3,8) ,
34295	 => std_logic_vector(to_unsigned(16,8) ,
34296	 => std_logic_vector(to_unsigned(9,8) ,
34297	 => std_logic_vector(to_unsigned(6,8) ,
34298	 => std_logic_vector(to_unsigned(6,8) ,
34299	 => std_logic_vector(to_unsigned(5,8) ,
34300	 => std_logic_vector(to_unsigned(5,8) ,
34301	 => std_logic_vector(to_unsigned(5,8) ,
34302	 => std_logic_vector(to_unsigned(2,8) ,
34303	 => std_logic_vector(to_unsigned(2,8) ,
34304	 => std_logic_vector(to_unsigned(2,8) ,
34305	 => std_logic_vector(to_unsigned(1,8) ,
34306	 => std_logic_vector(to_unsigned(1,8) ,
34307	 => std_logic_vector(to_unsigned(1,8) ,
34308	 => std_logic_vector(to_unsigned(1,8) ,
34309	 => std_logic_vector(to_unsigned(1,8) ,
34310	 => std_logic_vector(to_unsigned(2,8) ,
34311	 => std_logic_vector(to_unsigned(2,8) ,
34312	 => std_logic_vector(to_unsigned(4,8) ,
34313	 => std_logic_vector(to_unsigned(8,8) ,
34314	 => std_logic_vector(to_unsigned(11,8) ,
34315	 => std_logic_vector(to_unsigned(12,8) ,
34316	 => std_logic_vector(to_unsigned(3,8) ,
34317	 => std_logic_vector(to_unsigned(1,8) ,
34318	 => std_logic_vector(to_unsigned(7,8) ,
34319	 => std_logic_vector(to_unsigned(7,8) ,
34320	 => std_logic_vector(to_unsigned(7,8) ,
34321	 => std_logic_vector(to_unsigned(4,8) ,
34322	 => std_logic_vector(to_unsigned(2,8) ,
34323	 => std_logic_vector(to_unsigned(1,8) ,
34324	 => std_logic_vector(to_unsigned(1,8) ,
34325	 => std_logic_vector(to_unsigned(0,8) ,
34326	 => std_logic_vector(to_unsigned(0,8) ,
34327	 => std_logic_vector(to_unsigned(0,8) ,
34328	 => std_logic_vector(to_unsigned(0,8) ,
34329	 => std_logic_vector(to_unsigned(0,8) ,
34330	 => std_logic_vector(to_unsigned(1,8) ,
34331	 => std_logic_vector(to_unsigned(5,8) ,
34332	 => std_logic_vector(to_unsigned(8,8) ,
34333	 => std_logic_vector(to_unsigned(10,8) ,
34334	 => std_logic_vector(to_unsigned(11,8) ,
34335	 => std_logic_vector(to_unsigned(8,8) ,
34336	 => std_logic_vector(to_unsigned(10,8) ,
34337	 => std_logic_vector(to_unsigned(7,8) ,
34338	 => std_logic_vector(to_unsigned(4,8) ,
34339	 => std_logic_vector(to_unsigned(7,8) ,
34340	 => std_logic_vector(to_unsigned(10,8) ,
34341	 => std_logic_vector(to_unsigned(10,8) ,
34342	 => std_logic_vector(to_unsigned(4,8) ,
34343	 => std_logic_vector(to_unsigned(3,8) ,
34344	 => std_logic_vector(to_unsigned(2,8) ,
34345	 => std_logic_vector(to_unsigned(1,8) ,
34346	 => std_logic_vector(to_unsigned(5,8) ,
34347	 => std_logic_vector(to_unsigned(51,8) ,
34348	 => std_logic_vector(to_unsigned(25,8) ,
34349	 => std_logic_vector(to_unsigned(5,8) ,
34350	 => std_logic_vector(to_unsigned(2,8) ,
34351	 => std_logic_vector(to_unsigned(4,8) ,
34352	 => std_logic_vector(to_unsigned(7,8) ,
34353	 => std_logic_vector(to_unsigned(5,8) ,
34354	 => std_logic_vector(to_unsigned(2,8) ,
34355	 => std_logic_vector(to_unsigned(1,8) ,
34356	 => std_logic_vector(to_unsigned(0,8) ,
34357	 => std_logic_vector(to_unsigned(0,8) ,
34358	 => std_logic_vector(to_unsigned(0,8) ,
34359	 => std_logic_vector(to_unsigned(0,8) ,
34360	 => std_logic_vector(to_unsigned(0,8) ,
34361	 => std_logic_vector(to_unsigned(1,8) ,
34362	 => std_logic_vector(to_unsigned(2,8) ,
34363	 => std_logic_vector(to_unsigned(2,8) ,
34364	 => std_logic_vector(to_unsigned(5,8) ,
34365	 => std_logic_vector(to_unsigned(10,8) ,
34366	 => std_logic_vector(to_unsigned(17,8) ,
34367	 => std_logic_vector(to_unsigned(16,8) ,
34368	 => std_logic_vector(to_unsigned(6,8) ,
34369	 => std_logic_vector(to_unsigned(2,8) ,
34370	 => std_logic_vector(to_unsigned(7,8) ,
34371	 => std_logic_vector(to_unsigned(68,8) ,
34372	 => std_logic_vector(to_unsigned(64,8) ,
34373	 => std_logic_vector(to_unsigned(44,8) ,
34374	 => std_logic_vector(to_unsigned(35,8) ,
34375	 => std_logic_vector(to_unsigned(25,8) ,
34376	 => std_logic_vector(to_unsigned(17,8) ,
34377	 => std_logic_vector(to_unsigned(11,8) ,
34378	 => std_logic_vector(to_unsigned(5,8) ,
34379	 => std_logic_vector(to_unsigned(4,8) ,
34380	 => std_logic_vector(to_unsigned(2,8) ,
34381	 => std_logic_vector(to_unsigned(1,8) ,
34382	 => std_logic_vector(to_unsigned(0,8) ,
34383	 => std_logic_vector(to_unsigned(1,8) ,
34384	 => std_logic_vector(to_unsigned(0,8) ,
34385	 => std_logic_vector(to_unsigned(1,8) ,
34386	 => std_logic_vector(to_unsigned(4,8) ,
34387	 => std_logic_vector(to_unsigned(6,8) ,
34388	 => std_logic_vector(to_unsigned(2,8) ,
34389	 => std_logic_vector(to_unsigned(1,8) ,
34390	 => std_logic_vector(to_unsigned(0,8) ,
34391	 => std_logic_vector(to_unsigned(0,8) ,
34392	 => std_logic_vector(to_unsigned(2,8) ,
34393	 => std_logic_vector(to_unsigned(2,8) ,
34394	 => std_logic_vector(to_unsigned(4,8) ,
34395	 => std_logic_vector(to_unsigned(8,8) ,
34396	 => std_logic_vector(to_unsigned(7,8) ,
34397	 => std_logic_vector(to_unsigned(2,8) ,
34398	 => std_logic_vector(to_unsigned(6,8) ,
34399	 => std_logic_vector(to_unsigned(10,8) ,
34400	 => std_logic_vector(to_unsigned(9,8) ,
34401	 => std_logic_vector(to_unsigned(6,8) ,
34402	 => std_logic_vector(to_unsigned(6,8) ,
34403	 => std_logic_vector(to_unsigned(5,8) ,
34404	 => std_logic_vector(to_unsigned(3,8) ,
34405	 => std_logic_vector(to_unsigned(3,8) ,
34406	 => std_logic_vector(to_unsigned(2,8) ,
34407	 => std_logic_vector(to_unsigned(1,8) ,
34408	 => std_logic_vector(to_unsigned(0,8) ,
34409	 => std_logic_vector(to_unsigned(0,8) ,
34410	 => std_logic_vector(to_unsigned(1,8) ,
34411	 => std_logic_vector(to_unsigned(1,8) ,
34412	 => std_logic_vector(to_unsigned(0,8) ,
34413	 => std_logic_vector(to_unsigned(0,8) ,
34414	 => std_logic_vector(to_unsigned(3,8) ,
34415	 => std_logic_vector(to_unsigned(6,8) ,
34416	 => std_logic_vector(to_unsigned(7,8) ,
34417	 => std_logic_vector(to_unsigned(8,8) ,
34418	 => std_logic_vector(to_unsigned(7,8) ,
34419	 => std_logic_vector(to_unsigned(3,8) ,
34420	 => std_logic_vector(to_unsigned(4,8) ,
34421	 => std_logic_vector(to_unsigned(2,8) ,
34422	 => std_logic_vector(to_unsigned(5,8) ,
34423	 => std_logic_vector(to_unsigned(4,8) ,
34424	 => std_logic_vector(to_unsigned(4,8) ,
34425	 => std_logic_vector(to_unsigned(2,8) ,
34426	 => std_logic_vector(to_unsigned(4,8) ,
34427	 => std_logic_vector(to_unsigned(16,8) ,
34428	 => std_logic_vector(to_unsigned(8,8) ,
34429	 => std_logic_vector(to_unsigned(7,8) ,
34430	 => std_logic_vector(to_unsigned(8,8) ,
34431	 => std_logic_vector(to_unsigned(3,8) ,
34432	 => std_logic_vector(to_unsigned(1,8) ,
34433	 => std_logic_vector(to_unsigned(2,8) ,
34434	 => std_logic_vector(to_unsigned(2,8) ,
34435	 => std_logic_vector(to_unsigned(1,8) ,
34436	 => std_logic_vector(to_unsigned(3,8) ,
34437	 => std_logic_vector(to_unsigned(3,8) ,
34438	 => std_logic_vector(to_unsigned(2,8) ,
34439	 => std_logic_vector(to_unsigned(2,8) ,
34440	 => std_logic_vector(to_unsigned(1,8) ,
34441	 => std_logic_vector(to_unsigned(1,8) ,
34442	 => std_logic_vector(to_unsigned(1,8) ,
34443	 => std_logic_vector(to_unsigned(1,8) ,
34444	 => std_logic_vector(to_unsigned(0,8) ,
34445	 => std_logic_vector(to_unsigned(0,8) ,
34446	 => std_logic_vector(to_unsigned(1,8) ,
34447	 => std_logic_vector(to_unsigned(0,8) ,
34448	 => std_logic_vector(to_unsigned(0,8) ,
34449	 => std_logic_vector(to_unsigned(30,8) ,
34450	 => std_logic_vector(to_unsigned(122,8) ,
34451	 => std_logic_vector(to_unsigned(168,8) ,
34452	 => std_logic_vector(to_unsigned(173,8) ,
34453	 => std_logic_vector(to_unsigned(161,8) ,
34454	 => std_logic_vector(to_unsigned(154,8) ,
34455	 => std_logic_vector(to_unsigned(152,8) ,
34456	 => std_logic_vector(to_unsigned(157,8) ,
34457	 => std_logic_vector(to_unsigned(156,8) ,
34458	 => std_logic_vector(to_unsigned(154,8) ,
34459	 => std_logic_vector(to_unsigned(152,8) ,
34460	 => std_logic_vector(to_unsigned(154,8) ,
34461	 => std_logic_vector(to_unsigned(159,8) ,
34462	 => std_logic_vector(to_unsigned(149,8) ,
34463	 => std_logic_vector(to_unsigned(149,8) ,
34464	 => std_logic_vector(to_unsigned(146,8) ,
34465	 => std_logic_vector(to_unsigned(151,8) ,
34466	 => std_logic_vector(to_unsigned(128,8) ,
34467	 => std_logic_vector(to_unsigned(10,8) ,
34468	 => std_logic_vector(to_unsigned(0,8) ,
34469	 => std_logic_vector(to_unsigned(1,8) ,
34470	 => std_logic_vector(to_unsigned(0,8) ,
34471	 => std_logic_vector(to_unsigned(0,8) ,
34472	 => std_logic_vector(to_unsigned(0,8) ,
34473	 => std_logic_vector(to_unsigned(1,8) ,
34474	 => std_logic_vector(to_unsigned(2,8) ,
34475	 => std_logic_vector(to_unsigned(2,8) ,
34476	 => std_logic_vector(to_unsigned(4,8) ,
34477	 => std_logic_vector(to_unsigned(8,8) ,
34478	 => std_logic_vector(to_unsigned(12,8) ,
34479	 => std_logic_vector(to_unsigned(8,8) ,
34480	 => std_logic_vector(to_unsigned(51,8) ,
34481	 => std_logic_vector(to_unsigned(156,8) ,
34482	 => std_logic_vector(to_unsigned(154,8) ,
34483	 => std_logic_vector(to_unsigned(152,8) ,
34484	 => std_logic_vector(to_unsigned(30,8) ,
34485	 => std_logic_vector(to_unsigned(2,8) ,
34486	 => std_logic_vector(to_unsigned(23,8) ,
34487	 => std_logic_vector(to_unsigned(139,8) ,
34488	 => std_logic_vector(to_unsigned(152,8) ,
34489	 => std_logic_vector(to_unsigned(156,8) ,
34490	 => std_logic_vector(to_unsigned(157,8) ,
34491	 => std_logic_vector(to_unsigned(154,8) ,
34492	 => std_logic_vector(to_unsigned(166,8) ,
34493	 => std_logic_vector(to_unsigned(108,8) ,
34494	 => std_logic_vector(to_unsigned(45,8) ,
34495	 => std_logic_vector(to_unsigned(35,8) ,
34496	 => std_logic_vector(to_unsigned(17,8) ,
34497	 => std_logic_vector(to_unsigned(18,8) ,
34498	 => std_logic_vector(to_unsigned(27,8) ,
34499	 => std_logic_vector(to_unsigned(18,8) ,
34500	 => std_logic_vector(to_unsigned(9,8) ,
34501	 => std_logic_vector(to_unsigned(30,8) ,
34502	 => std_logic_vector(to_unsigned(16,8) ,
34503	 => std_logic_vector(to_unsigned(7,8) ,
34504	 => std_logic_vector(to_unsigned(5,8) ,
34505	 => std_logic_vector(to_unsigned(14,8) ,
34506	 => std_logic_vector(to_unsigned(38,8) ,
34507	 => std_logic_vector(to_unsigned(8,8) ,
34508	 => std_logic_vector(to_unsigned(13,8) ,
34509	 => std_logic_vector(to_unsigned(112,8) ,
34510	 => std_logic_vector(to_unsigned(118,8) ,
34511	 => std_logic_vector(to_unsigned(146,8) ,
34512	 => std_logic_vector(to_unsigned(35,8) ,
34513	 => std_logic_vector(to_unsigned(1,8) ,
34514	 => std_logic_vector(to_unsigned(5,8) ,
34515	 => std_logic_vector(to_unsigned(10,8) ,
34516	 => std_logic_vector(to_unsigned(11,8) ,
34517	 => std_logic_vector(to_unsigned(10,8) ,
34518	 => std_logic_vector(to_unsigned(8,8) ,
34519	 => std_logic_vector(to_unsigned(4,8) ,
34520	 => std_logic_vector(to_unsigned(2,8) ,
34521	 => std_logic_vector(to_unsigned(5,8) ,
34522	 => std_logic_vector(to_unsigned(5,8) ,
34523	 => std_logic_vector(to_unsigned(4,8) ,
34524	 => std_logic_vector(to_unsigned(2,8) ,
34525	 => std_logic_vector(to_unsigned(1,8) ,
34526	 => std_logic_vector(to_unsigned(2,8) ,
34527	 => std_logic_vector(to_unsigned(6,8) ,
34528	 => std_logic_vector(to_unsigned(4,8) ,
34529	 => std_logic_vector(to_unsigned(7,8) ,
34530	 => std_logic_vector(to_unsigned(32,8) ,
34531	 => std_logic_vector(to_unsigned(29,8) ,
34532	 => std_logic_vector(to_unsigned(90,8) ,
34533	 => std_logic_vector(to_unsigned(99,8) ,
34534	 => std_logic_vector(to_unsigned(29,8) ,
34535	 => std_logic_vector(to_unsigned(81,8) ,
34536	 => std_logic_vector(to_unsigned(154,8) ,
34537	 => std_logic_vector(to_unsigned(152,8) ,
34538	 => std_logic_vector(to_unsigned(128,8) ,
34539	 => std_logic_vector(to_unsigned(79,8) ,
34540	 => std_logic_vector(to_unsigned(55,8) ,
34541	 => std_logic_vector(to_unsigned(81,8) ,
34542	 => std_logic_vector(to_unsigned(139,8) ,
34543	 => std_logic_vector(to_unsigned(121,8) ,
34544	 => std_logic_vector(to_unsigned(37,8) ,
34545	 => std_logic_vector(to_unsigned(13,8) ,
34546	 => std_logic_vector(to_unsigned(71,8) ,
34547	 => std_logic_vector(to_unsigned(139,8) ,
34548	 => std_logic_vector(to_unsigned(119,8) ,
34549	 => std_logic_vector(to_unsigned(118,8) ,
34550	 => std_logic_vector(to_unsigned(114,8) ,
34551	 => std_logic_vector(to_unsigned(119,8) ,
34552	 => std_logic_vector(to_unsigned(128,8) ,
34553	 => std_logic_vector(to_unsigned(114,8) ,
34554	 => std_logic_vector(to_unsigned(116,8) ,
34555	 => std_logic_vector(to_unsigned(136,8) ,
34556	 => std_logic_vector(to_unsigned(112,8) ,
34557	 => std_logic_vector(to_unsigned(97,8) ,
34558	 => std_logic_vector(to_unsigned(105,8) ,
34559	 => std_logic_vector(to_unsigned(107,8) ,
34560	 => std_logic_vector(to_unsigned(108,8) ,
34561	 => std_logic_vector(to_unsigned(9,8) ,
34562	 => std_logic_vector(to_unsigned(8,8) ,
34563	 => std_logic_vector(to_unsigned(7,8) ,
34564	 => std_logic_vector(to_unsigned(7,8) ,
34565	 => std_logic_vector(to_unsigned(6,8) ,
34566	 => std_logic_vector(to_unsigned(7,8) ,
34567	 => std_logic_vector(to_unsigned(7,8) ,
34568	 => std_logic_vector(to_unsigned(7,8) ,
34569	 => std_logic_vector(to_unsigned(3,8) ,
34570	 => std_logic_vector(to_unsigned(2,8) ,
34571	 => std_logic_vector(to_unsigned(2,8) ,
34572	 => std_logic_vector(to_unsigned(1,8) ,
34573	 => std_logic_vector(to_unsigned(1,8) ,
34574	 => std_logic_vector(to_unsigned(1,8) ,
34575	 => std_logic_vector(to_unsigned(1,8) ,
34576	 => std_logic_vector(to_unsigned(0,8) ,
34577	 => std_logic_vector(to_unsigned(0,8) ,
34578	 => std_logic_vector(to_unsigned(1,8) ,
34579	 => std_logic_vector(to_unsigned(2,8) ,
34580	 => std_logic_vector(to_unsigned(1,8) ,
34581	 => std_logic_vector(to_unsigned(0,8) ,
34582	 => std_logic_vector(to_unsigned(0,8) ,
34583	 => std_logic_vector(to_unsigned(0,8) ,
34584	 => std_logic_vector(to_unsigned(0,8) ,
34585	 => std_logic_vector(to_unsigned(0,8) ,
34586	 => std_logic_vector(to_unsigned(0,8) ,
34587	 => std_logic_vector(to_unsigned(0,8) ,
34588	 => std_logic_vector(to_unsigned(2,8) ,
34589	 => std_logic_vector(to_unsigned(13,8) ,
34590	 => std_logic_vector(to_unsigned(9,8) ,
34591	 => std_logic_vector(to_unsigned(8,8) ,
34592	 => std_logic_vector(to_unsigned(7,8) ,
34593	 => std_logic_vector(to_unsigned(18,8) ,
34594	 => std_logic_vector(to_unsigned(35,8) ,
34595	 => std_logic_vector(to_unsigned(35,8) ,
34596	 => std_logic_vector(to_unsigned(32,8) ,
34597	 => std_logic_vector(to_unsigned(22,8) ,
34598	 => std_logic_vector(to_unsigned(14,8) ,
34599	 => std_logic_vector(to_unsigned(6,8) ,
34600	 => std_logic_vector(to_unsigned(17,8) ,
34601	 => std_logic_vector(to_unsigned(24,8) ,
34602	 => std_logic_vector(to_unsigned(17,8) ,
34603	 => std_logic_vector(to_unsigned(14,8) ,
34604	 => std_logic_vector(to_unsigned(4,8) ,
34605	 => std_logic_vector(to_unsigned(3,8) ,
34606	 => std_logic_vector(to_unsigned(2,8) ,
34607	 => std_logic_vector(to_unsigned(0,8) ,
34608	 => std_logic_vector(to_unsigned(0,8) ,
34609	 => std_logic_vector(to_unsigned(0,8) ,
34610	 => std_logic_vector(to_unsigned(0,8) ,
34611	 => std_logic_vector(to_unsigned(0,8) ,
34612	 => std_logic_vector(to_unsigned(3,8) ,
34613	 => std_logic_vector(to_unsigned(7,8) ,
34614	 => std_logic_vector(to_unsigned(3,8) ,
34615	 => std_logic_vector(to_unsigned(11,8) ,
34616	 => std_logic_vector(to_unsigned(10,8) ,
34617	 => std_logic_vector(to_unsigned(6,8) ,
34618	 => std_logic_vector(to_unsigned(6,8) ,
34619	 => std_logic_vector(to_unsigned(9,8) ,
34620	 => std_logic_vector(to_unsigned(7,8) ,
34621	 => std_logic_vector(to_unsigned(5,8) ,
34622	 => std_logic_vector(to_unsigned(3,8) ,
34623	 => std_logic_vector(to_unsigned(2,8) ,
34624	 => std_logic_vector(to_unsigned(1,8) ,
34625	 => std_logic_vector(to_unsigned(1,8) ,
34626	 => std_logic_vector(to_unsigned(1,8) ,
34627	 => std_logic_vector(to_unsigned(1,8) ,
34628	 => std_logic_vector(to_unsigned(1,8) ,
34629	 => std_logic_vector(to_unsigned(2,8) ,
34630	 => std_logic_vector(to_unsigned(3,8) ,
34631	 => std_logic_vector(to_unsigned(5,8) ,
34632	 => std_logic_vector(to_unsigned(9,8) ,
34633	 => std_logic_vector(to_unsigned(10,8) ,
34634	 => std_logic_vector(to_unsigned(11,8) ,
34635	 => std_logic_vector(to_unsigned(12,8) ,
34636	 => std_logic_vector(to_unsigned(2,8) ,
34637	 => std_logic_vector(to_unsigned(2,8) ,
34638	 => std_logic_vector(to_unsigned(9,8) ,
34639	 => std_logic_vector(to_unsigned(7,8) ,
34640	 => std_logic_vector(to_unsigned(7,8) ,
34641	 => std_logic_vector(to_unsigned(5,8) ,
34642	 => std_logic_vector(to_unsigned(3,8) ,
34643	 => std_logic_vector(to_unsigned(2,8) ,
34644	 => std_logic_vector(to_unsigned(1,8) ,
34645	 => std_logic_vector(to_unsigned(2,8) ,
34646	 => std_logic_vector(to_unsigned(1,8) ,
34647	 => std_logic_vector(to_unsigned(0,8) ,
34648	 => std_logic_vector(to_unsigned(0,8) ,
34649	 => std_logic_vector(to_unsigned(0,8) ,
34650	 => std_logic_vector(to_unsigned(1,8) ,
34651	 => std_logic_vector(to_unsigned(6,8) ,
34652	 => std_logic_vector(to_unsigned(8,8) ,
34653	 => std_logic_vector(to_unsigned(14,8) ,
34654	 => std_logic_vector(to_unsigned(11,8) ,
34655	 => std_logic_vector(to_unsigned(10,8) ,
34656	 => std_logic_vector(to_unsigned(9,8) ,
34657	 => std_logic_vector(to_unsigned(6,8) ,
34658	 => std_logic_vector(to_unsigned(3,8) ,
34659	 => std_logic_vector(to_unsigned(7,8) ,
34660	 => std_logic_vector(to_unsigned(10,8) ,
34661	 => std_logic_vector(to_unsigned(17,8) ,
34662	 => std_logic_vector(to_unsigned(10,8) ,
34663	 => std_logic_vector(to_unsigned(5,8) ,
34664	 => std_logic_vector(to_unsigned(4,8) ,
34665	 => std_logic_vector(to_unsigned(3,8) ,
34666	 => std_logic_vector(to_unsigned(1,8) ,
34667	 => std_logic_vector(to_unsigned(4,8) ,
34668	 => std_logic_vector(to_unsigned(17,8) ,
34669	 => std_logic_vector(to_unsigned(9,8) ,
34670	 => std_logic_vector(to_unsigned(4,8) ,
34671	 => std_logic_vector(to_unsigned(4,8) ,
34672	 => std_logic_vector(to_unsigned(4,8) ,
34673	 => std_logic_vector(to_unsigned(1,8) ,
34674	 => std_logic_vector(to_unsigned(0,8) ,
34675	 => std_logic_vector(to_unsigned(0,8) ,
34676	 => std_logic_vector(to_unsigned(0,8) ,
34677	 => std_logic_vector(to_unsigned(0,8) ,
34678	 => std_logic_vector(to_unsigned(0,8) ,
34679	 => std_logic_vector(to_unsigned(0,8) ,
34680	 => std_logic_vector(to_unsigned(0,8) ,
34681	 => std_logic_vector(to_unsigned(2,8) ,
34682	 => std_logic_vector(to_unsigned(4,8) ,
34683	 => std_logic_vector(to_unsigned(5,8) ,
34684	 => std_logic_vector(to_unsigned(5,8) ,
34685	 => std_logic_vector(to_unsigned(8,8) ,
34686	 => std_logic_vector(to_unsigned(27,8) ,
34687	 => std_logic_vector(to_unsigned(17,8) ,
34688	 => std_logic_vector(to_unsigned(4,8) ,
34689	 => std_logic_vector(to_unsigned(1,8) ,
34690	 => std_logic_vector(to_unsigned(1,8) ,
34691	 => std_logic_vector(to_unsigned(3,8) ,
34692	 => std_logic_vector(to_unsigned(1,8) ,
34693	 => std_logic_vector(to_unsigned(1,8) ,
34694	 => std_logic_vector(to_unsigned(1,8) ,
34695	 => std_logic_vector(to_unsigned(1,8) ,
34696	 => std_logic_vector(to_unsigned(2,8) ,
34697	 => std_logic_vector(to_unsigned(1,8) ,
34698	 => std_logic_vector(to_unsigned(0,8) ,
34699	 => std_logic_vector(to_unsigned(2,8) ,
34700	 => std_logic_vector(to_unsigned(2,8) ,
34701	 => std_logic_vector(to_unsigned(1,8) ,
34702	 => std_logic_vector(to_unsigned(1,8) ,
34703	 => std_logic_vector(to_unsigned(2,8) ,
34704	 => std_logic_vector(to_unsigned(6,8) ,
34705	 => std_logic_vector(to_unsigned(7,8) ,
34706	 => std_logic_vector(to_unsigned(5,8) ,
34707	 => std_logic_vector(to_unsigned(3,8) ,
34708	 => std_logic_vector(to_unsigned(4,8) ,
34709	 => std_logic_vector(to_unsigned(3,8) ,
34710	 => std_logic_vector(to_unsigned(3,8) ,
34711	 => std_logic_vector(to_unsigned(1,8) ,
34712	 => std_logic_vector(to_unsigned(2,8) ,
34713	 => std_logic_vector(to_unsigned(2,8) ,
34714	 => std_logic_vector(to_unsigned(5,8) ,
34715	 => std_logic_vector(to_unsigned(11,8) ,
34716	 => std_logic_vector(to_unsigned(5,8) ,
34717	 => std_logic_vector(to_unsigned(3,8) ,
34718	 => std_logic_vector(to_unsigned(5,8) ,
34719	 => std_logic_vector(to_unsigned(8,8) ,
34720	 => std_logic_vector(to_unsigned(10,8) ,
34721	 => std_logic_vector(to_unsigned(5,8) ,
34722	 => std_logic_vector(to_unsigned(5,8) ,
34723	 => std_logic_vector(to_unsigned(7,8) ,
34724	 => std_logic_vector(to_unsigned(6,8) ,
34725	 => std_logic_vector(to_unsigned(3,8) ,
34726	 => std_logic_vector(to_unsigned(1,8) ,
34727	 => std_logic_vector(to_unsigned(0,8) ,
34728	 => std_logic_vector(to_unsigned(1,8) ,
34729	 => std_logic_vector(to_unsigned(0,8) ,
34730	 => std_logic_vector(to_unsigned(0,8) ,
34731	 => std_logic_vector(to_unsigned(0,8) ,
34732	 => std_logic_vector(to_unsigned(0,8) ,
34733	 => std_logic_vector(to_unsigned(0,8) ,
34734	 => std_logic_vector(to_unsigned(3,8) ,
34735	 => std_logic_vector(to_unsigned(5,8) ,
34736	 => std_logic_vector(to_unsigned(6,8) ,
34737	 => std_logic_vector(to_unsigned(8,8) ,
34738	 => std_logic_vector(to_unsigned(8,8) ,
34739	 => std_logic_vector(to_unsigned(3,8) ,
34740	 => std_logic_vector(to_unsigned(1,8) ,
34741	 => std_logic_vector(to_unsigned(1,8) ,
34742	 => std_logic_vector(to_unsigned(4,8) ,
34743	 => std_logic_vector(to_unsigned(5,8) ,
34744	 => std_logic_vector(to_unsigned(3,8) ,
34745	 => std_logic_vector(to_unsigned(2,8) ,
34746	 => std_logic_vector(to_unsigned(2,8) ,
34747	 => std_logic_vector(to_unsigned(10,8) ,
34748	 => std_logic_vector(to_unsigned(9,8) ,
34749	 => std_logic_vector(to_unsigned(4,8) ,
34750	 => std_logic_vector(to_unsigned(2,8) ,
34751	 => std_logic_vector(to_unsigned(1,8) ,
34752	 => std_logic_vector(to_unsigned(0,8) ,
34753	 => std_logic_vector(to_unsigned(1,8) ,
34754	 => std_logic_vector(to_unsigned(1,8) ,
34755	 => std_logic_vector(to_unsigned(1,8) ,
34756	 => std_logic_vector(to_unsigned(1,8) ,
34757	 => std_logic_vector(to_unsigned(1,8) ,
34758	 => std_logic_vector(to_unsigned(1,8) ,
34759	 => std_logic_vector(to_unsigned(1,8) ,
34760	 => std_logic_vector(to_unsigned(1,8) ,
34761	 => std_logic_vector(to_unsigned(1,8) ,
34762	 => std_logic_vector(to_unsigned(0,8) ,
34763	 => std_logic_vector(to_unsigned(0,8) ,
34764	 => std_logic_vector(to_unsigned(0,8) ,
34765	 => std_logic_vector(to_unsigned(0,8) ,
34766	 => std_logic_vector(to_unsigned(0,8) ,
34767	 => std_logic_vector(to_unsigned(1,8) ,
34768	 => std_logic_vector(to_unsigned(1,8) ,
34769	 => std_logic_vector(to_unsigned(1,8) ,
34770	 => std_logic_vector(to_unsigned(6,8) ,
34771	 => std_logic_vector(to_unsigned(27,8) ,
34772	 => std_logic_vector(to_unsigned(90,8) ,
34773	 => std_logic_vector(to_unsigned(157,8) ,
34774	 => std_logic_vector(to_unsigned(179,8) ,
34775	 => std_logic_vector(to_unsigned(168,8) ,
34776	 => std_logic_vector(to_unsigned(154,8) ,
34777	 => std_logic_vector(to_unsigned(151,8) ,
34778	 => std_logic_vector(to_unsigned(152,8) ,
34779	 => std_logic_vector(to_unsigned(154,8) ,
34780	 => std_logic_vector(to_unsigned(154,8) ,
34781	 => std_logic_vector(to_unsigned(159,8) ,
34782	 => std_logic_vector(to_unsigned(156,8) ,
34783	 => std_logic_vector(to_unsigned(152,8) ,
34784	 => std_logic_vector(to_unsigned(149,8) ,
34785	 => std_logic_vector(to_unsigned(154,8) ,
34786	 => std_logic_vector(to_unsigned(101,8) ,
34787	 => std_logic_vector(to_unsigned(9,8) ,
34788	 => std_logic_vector(to_unsigned(0,8) ,
34789	 => std_logic_vector(to_unsigned(1,8) ,
34790	 => std_logic_vector(to_unsigned(1,8) ,
34791	 => std_logic_vector(to_unsigned(1,8) ,
34792	 => std_logic_vector(to_unsigned(2,8) ,
34793	 => std_logic_vector(to_unsigned(2,8) ,
34794	 => std_logic_vector(to_unsigned(2,8) ,
34795	 => std_logic_vector(to_unsigned(1,8) ,
34796	 => std_logic_vector(to_unsigned(2,8) ,
34797	 => std_logic_vector(to_unsigned(5,8) ,
34798	 => std_logic_vector(to_unsigned(9,8) ,
34799	 => std_logic_vector(to_unsigned(18,8) ,
34800	 => std_logic_vector(to_unsigned(111,8) ,
34801	 => std_logic_vector(to_unsigned(164,8) ,
34802	 => std_logic_vector(to_unsigned(147,8) ,
34803	 => std_logic_vector(to_unsigned(161,8) ,
34804	 => std_logic_vector(to_unsigned(38,8) ,
34805	 => std_logic_vector(to_unsigned(2,8) ,
34806	 => std_logic_vector(to_unsigned(27,8) ,
34807	 => std_logic_vector(to_unsigned(144,8) ,
34808	 => std_logic_vector(to_unsigned(159,8) ,
34809	 => std_logic_vector(to_unsigned(149,8) ,
34810	 => std_logic_vector(to_unsigned(152,8) ,
34811	 => std_logic_vector(to_unsigned(151,8) ,
34812	 => std_logic_vector(to_unsigned(177,8) ,
34813	 => std_logic_vector(to_unsigned(60,8) ,
34814	 => std_logic_vector(to_unsigned(1,8) ,
34815	 => std_logic_vector(to_unsigned(4,8) ,
34816	 => std_logic_vector(to_unsigned(5,8) ,
34817	 => std_logic_vector(to_unsigned(4,8) ,
34818	 => std_logic_vector(to_unsigned(6,8) ,
34819	 => std_logic_vector(to_unsigned(8,8) ,
34820	 => std_logic_vector(to_unsigned(6,8) ,
34821	 => std_logic_vector(to_unsigned(36,8) ,
34822	 => std_logic_vector(to_unsigned(51,8) ,
34823	 => std_logic_vector(to_unsigned(10,8) ,
34824	 => std_logic_vector(to_unsigned(5,8) ,
34825	 => std_logic_vector(to_unsigned(11,8) ,
34826	 => std_logic_vector(to_unsigned(36,8) ,
34827	 => std_logic_vector(to_unsigned(20,8) ,
34828	 => std_logic_vector(to_unsigned(5,8) ,
34829	 => std_logic_vector(to_unsigned(93,8) ,
34830	 => std_logic_vector(to_unsigned(119,8) ,
34831	 => std_logic_vector(to_unsigned(133,8) ,
34832	 => std_logic_vector(to_unsigned(65,8) ,
34833	 => std_logic_vector(to_unsigned(4,8) ,
34834	 => std_logic_vector(to_unsigned(6,8) ,
34835	 => std_logic_vector(to_unsigned(12,8) ,
34836	 => std_logic_vector(to_unsigned(8,8) ,
34837	 => std_logic_vector(to_unsigned(7,8) ,
34838	 => std_logic_vector(to_unsigned(11,8) ,
34839	 => std_logic_vector(to_unsigned(16,8) ,
34840	 => std_logic_vector(to_unsigned(11,8) ,
34841	 => std_logic_vector(to_unsigned(19,8) ,
34842	 => std_logic_vector(to_unsigned(25,8) ,
34843	 => std_logic_vector(to_unsigned(15,8) ,
34844	 => std_logic_vector(to_unsigned(12,8) ,
34845	 => std_logic_vector(to_unsigned(4,8) ,
34846	 => std_logic_vector(to_unsigned(1,8) ,
34847	 => std_logic_vector(to_unsigned(1,8) ,
34848	 => std_logic_vector(to_unsigned(17,8) ,
34849	 => std_logic_vector(to_unsigned(104,8) ,
34850	 => std_logic_vector(to_unsigned(181,8) ,
34851	 => std_logic_vector(to_unsigned(121,8) ,
34852	 => std_logic_vector(to_unsigned(77,8) ,
34853	 => std_logic_vector(to_unsigned(127,8) ,
34854	 => std_logic_vector(to_unsigned(112,8) ,
34855	 => std_logic_vector(to_unsigned(91,8) ,
34856	 => std_logic_vector(to_unsigned(130,8) ,
34857	 => std_logic_vector(to_unsigned(130,8) ,
34858	 => std_logic_vector(to_unsigned(116,8) ,
34859	 => std_logic_vector(to_unsigned(60,8) ,
34860	 => std_logic_vector(to_unsigned(47,8) ,
34861	 => std_logic_vector(to_unsigned(100,8) ,
34862	 => std_logic_vector(to_unsigned(136,8) ,
34863	 => std_logic_vector(to_unsigned(87,8) ,
34864	 => std_logic_vector(to_unsigned(4,8) ,
34865	 => std_logic_vector(to_unsigned(0,8) ,
34866	 => std_logic_vector(to_unsigned(21,8) ,
34867	 => std_logic_vector(to_unsigned(133,8) ,
34868	 => std_logic_vector(to_unsigned(134,8) ,
34869	 => std_logic_vector(to_unsigned(122,8) ,
34870	 => std_logic_vector(to_unsigned(131,8) ,
34871	 => std_logic_vector(to_unsigned(138,8) ,
34872	 => std_logic_vector(to_unsigned(119,8) ,
34873	 => std_logic_vector(to_unsigned(133,8) ,
34874	 => std_logic_vector(to_unsigned(142,8) ,
34875	 => std_logic_vector(to_unsigned(128,8) ,
34876	 => std_logic_vector(to_unsigned(121,8) ,
34877	 => std_logic_vector(to_unsigned(114,8) ,
34878	 => std_logic_vector(to_unsigned(107,8) ,
34879	 => std_logic_vector(to_unsigned(107,8) ,
34880	 => std_logic_vector(to_unsigned(105,8) ,
34881	 => std_logic_vector(to_unsigned(9,8) ,
34882	 => std_logic_vector(to_unsigned(8,8) ,
34883	 => std_logic_vector(to_unsigned(6,8) ,
34884	 => std_logic_vector(to_unsigned(6,8) ,
34885	 => std_logic_vector(to_unsigned(6,8) ,
34886	 => std_logic_vector(to_unsigned(6,8) ,
34887	 => std_logic_vector(to_unsigned(7,8) ,
34888	 => std_logic_vector(to_unsigned(7,8) ,
34889	 => std_logic_vector(to_unsigned(4,8) ,
34890	 => std_logic_vector(to_unsigned(2,8) ,
34891	 => std_logic_vector(to_unsigned(2,8) ,
34892	 => std_logic_vector(to_unsigned(1,8) ,
34893	 => std_logic_vector(to_unsigned(1,8) ,
34894	 => std_logic_vector(to_unsigned(1,8) ,
34895	 => std_logic_vector(to_unsigned(1,8) ,
34896	 => std_logic_vector(to_unsigned(0,8) ,
34897	 => std_logic_vector(to_unsigned(0,8) ,
34898	 => std_logic_vector(to_unsigned(1,8) ,
34899	 => std_logic_vector(to_unsigned(1,8) ,
34900	 => std_logic_vector(to_unsigned(0,8) ,
34901	 => std_logic_vector(to_unsigned(0,8) ,
34902	 => std_logic_vector(to_unsigned(0,8) ,
34903	 => std_logic_vector(to_unsigned(0,8) ,
34904	 => std_logic_vector(to_unsigned(0,8) ,
34905	 => std_logic_vector(to_unsigned(0,8) ,
34906	 => std_logic_vector(to_unsigned(0,8) ,
34907	 => std_logic_vector(to_unsigned(0,8) ,
34908	 => std_logic_vector(to_unsigned(0,8) ,
34909	 => std_logic_vector(to_unsigned(6,8) ,
34910	 => std_logic_vector(to_unsigned(15,8) ,
34911	 => std_logic_vector(to_unsigned(8,8) ,
34912	 => std_logic_vector(to_unsigned(4,8) ,
34913	 => std_logic_vector(to_unsigned(26,8) ,
34914	 => std_logic_vector(to_unsigned(33,8) ,
34915	 => std_logic_vector(to_unsigned(29,8) ,
34916	 => std_logic_vector(to_unsigned(30,8) ,
34917	 => std_logic_vector(to_unsigned(22,8) ,
34918	 => std_logic_vector(to_unsigned(12,8) ,
34919	 => std_logic_vector(to_unsigned(12,8) ,
34920	 => std_logic_vector(to_unsigned(20,8) ,
34921	 => std_logic_vector(to_unsigned(8,8) ,
34922	 => std_logic_vector(to_unsigned(5,8) ,
34923	 => std_logic_vector(to_unsigned(3,8) ,
34924	 => std_logic_vector(to_unsigned(3,8) ,
34925	 => std_logic_vector(to_unsigned(5,8) ,
34926	 => std_logic_vector(to_unsigned(2,8) ,
34927	 => std_logic_vector(to_unsigned(0,8) ,
34928	 => std_logic_vector(to_unsigned(0,8) ,
34929	 => std_logic_vector(to_unsigned(0,8) ,
34930	 => std_logic_vector(to_unsigned(0,8) ,
34931	 => std_logic_vector(to_unsigned(1,8) ,
34932	 => std_logic_vector(to_unsigned(2,8) ,
34933	 => std_logic_vector(to_unsigned(3,8) ,
34934	 => std_logic_vector(to_unsigned(3,8) ,
34935	 => std_logic_vector(to_unsigned(10,8) ,
34936	 => std_logic_vector(to_unsigned(10,8) ,
34937	 => std_logic_vector(to_unsigned(7,8) ,
34938	 => std_logic_vector(to_unsigned(6,8) ,
34939	 => std_logic_vector(to_unsigned(4,8) ,
34940	 => std_logic_vector(to_unsigned(8,8) ,
34941	 => std_logic_vector(to_unsigned(11,8) ,
34942	 => std_logic_vector(to_unsigned(6,8) ,
34943	 => std_logic_vector(to_unsigned(3,8) ,
34944	 => std_logic_vector(to_unsigned(3,8) ,
34945	 => std_logic_vector(to_unsigned(1,8) ,
34946	 => std_logic_vector(to_unsigned(1,8) ,
34947	 => std_logic_vector(to_unsigned(1,8) ,
34948	 => std_logic_vector(to_unsigned(0,8) ,
34949	 => std_logic_vector(to_unsigned(2,8) ,
34950	 => std_logic_vector(to_unsigned(7,8) ,
34951	 => std_logic_vector(to_unsigned(9,8) ,
34952	 => std_logic_vector(to_unsigned(10,8) ,
34953	 => std_logic_vector(to_unsigned(7,8) ,
34954	 => std_logic_vector(to_unsigned(9,8) ,
34955	 => std_logic_vector(to_unsigned(11,8) ,
34956	 => std_logic_vector(to_unsigned(1,8) ,
34957	 => std_logic_vector(to_unsigned(2,8) ,
34958	 => std_logic_vector(to_unsigned(8,8) ,
34959	 => std_logic_vector(to_unsigned(4,8) ,
34960	 => std_logic_vector(to_unsigned(5,8) ,
34961	 => std_logic_vector(to_unsigned(5,8) ,
34962	 => std_logic_vector(to_unsigned(5,8) ,
34963	 => std_logic_vector(to_unsigned(2,8) ,
34964	 => std_logic_vector(to_unsigned(1,8) ,
34965	 => std_logic_vector(to_unsigned(3,8) ,
34966	 => std_logic_vector(to_unsigned(2,8) ,
34967	 => std_logic_vector(to_unsigned(0,8) ,
34968	 => std_logic_vector(to_unsigned(0,8) ,
34969	 => std_logic_vector(to_unsigned(0,8) ,
34970	 => std_logic_vector(to_unsigned(0,8) ,
34971	 => std_logic_vector(to_unsigned(4,8) ,
34972	 => std_logic_vector(to_unsigned(9,8) ,
34973	 => std_logic_vector(to_unsigned(17,8) ,
34974	 => std_logic_vector(to_unsigned(10,8) ,
34975	 => std_logic_vector(to_unsigned(9,8) ,
34976	 => std_logic_vector(to_unsigned(9,8) ,
34977	 => std_logic_vector(to_unsigned(7,8) ,
34978	 => std_logic_vector(to_unsigned(5,8) ,
34979	 => std_logic_vector(to_unsigned(8,8) ,
34980	 => std_logic_vector(to_unsigned(10,8) ,
34981	 => std_logic_vector(to_unsigned(10,8) ,
34982	 => std_logic_vector(to_unsigned(21,8) ,
34983	 => std_logic_vector(to_unsigned(22,8) ,
34984	 => std_logic_vector(to_unsigned(17,8) ,
34985	 => std_logic_vector(to_unsigned(13,8) ,
34986	 => std_logic_vector(to_unsigned(5,8) ,
34987	 => std_logic_vector(to_unsigned(17,8) ,
34988	 => std_logic_vector(to_unsigned(61,8) ,
34989	 => std_logic_vector(to_unsigned(15,8) ,
34990	 => std_logic_vector(to_unsigned(3,8) ,
34991	 => std_logic_vector(to_unsigned(3,8) ,
34992	 => std_logic_vector(to_unsigned(1,8) ,
34993	 => std_logic_vector(to_unsigned(1,8) ,
34994	 => std_logic_vector(to_unsigned(0,8) ,
34995	 => std_logic_vector(to_unsigned(0,8) ,
34996	 => std_logic_vector(to_unsigned(0,8) ,
34997	 => std_logic_vector(to_unsigned(0,8) ,
34998	 => std_logic_vector(to_unsigned(0,8) ,
34999	 => std_logic_vector(to_unsigned(0,8) ,
35000	 => std_logic_vector(to_unsigned(0,8) ,
35001	 => std_logic_vector(to_unsigned(2,8) ,
35002	 => std_logic_vector(to_unsigned(6,8) ,
35003	 => std_logic_vector(to_unsigned(6,8) ,
35004	 => std_logic_vector(to_unsigned(5,8) ,
35005	 => std_logic_vector(to_unsigned(11,8) ,
35006	 => std_logic_vector(to_unsigned(15,8) ,
35007	 => std_logic_vector(to_unsigned(6,8) ,
35008	 => std_logic_vector(to_unsigned(3,8) ,
35009	 => std_logic_vector(to_unsigned(2,8) ,
35010	 => std_logic_vector(to_unsigned(0,8) ,
35011	 => std_logic_vector(to_unsigned(3,8) ,
35012	 => std_logic_vector(to_unsigned(4,8) ,
35013	 => std_logic_vector(to_unsigned(3,8) ,
35014	 => std_logic_vector(to_unsigned(3,8) ,
35015	 => std_logic_vector(to_unsigned(2,8) ,
35016	 => std_logic_vector(to_unsigned(3,8) ,
35017	 => std_logic_vector(to_unsigned(2,8) ,
35018	 => std_logic_vector(to_unsigned(1,8) ,
35019	 => std_logic_vector(to_unsigned(3,8) ,
35020	 => std_logic_vector(to_unsigned(3,8) ,
35021	 => std_logic_vector(to_unsigned(1,8) ,
35022	 => std_logic_vector(to_unsigned(1,8) ,
35023	 => std_logic_vector(to_unsigned(1,8) ,
35024	 => std_logic_vector(to_unsigned(1,8) ,
35025	 => std_logic_vector(to_unsigned(2,8) ,
35026	 => std_logic_vector(to_unsigned(1,8) ,
35027	 => std_logic_vector(to_unsigned(2,8) ,
35028	 => std_logic_vector(to_unsigned(4,8) ,
35029	 => std_logic_vector(to_unsigned(4,8) ,
35030	 => std_logic_vector(to_unsigned(5,8) ,
35031	 => std_logic_vector(to_unsigned(4,8) ,
35032	 => std_logic_vector(to_unsigned(3,8) ,
35033	 => std_logic_vector(to_unsigned(3,8) ,
35034	 => std_logic_vector(to_unsigned(5,8) ,
35035	 => std_logic_vector(to_unsigned(12,8) ,
35036	 => std_logic_vector(to_unsigned(6,8) ,
35037	 => std_logic_vector(to_unsigned(3,8) ,
35038	 => std_logic_vector(to_unsigned(4,8) ,
35039	 => std_logic_vector(to_unsigned(6,8) ,
35040	 => std_logic_vector(to_unsigned(11,8) ,
35041	 => std_logic_vector(to_unsigned(5,8) ,
35042	 => std_logic_vector(to_unsigned(5,8) ,
35043	 => std_logic_vector(to_unsigned(8,8) ,
35044	 => std_logic_vector(to_unsigned(8,8) ,
35045	 => std_logic_vector(to_unsigned(6,8) ,
35046	 => std_logic_vector(to_unsigned(3,8) ,
35047	 => std_logic_vector(to_unsigned(1,8) ,
35048	 => std_logic_vector(to_unsigned(1,8) ,
35049	 => std_logic_vector(to_unsigned(0,8) ,
35050	 => std_logic_vector(to_unsigned(1,8) ,
35051	 => std_logic_vector(to_unsigned(1,8) ,
35052	 => std_logic_vector(to_unsigned(1,8) ,
35053	 => std_logic_vector(to_unsigned(1,8) ,
35054	 => std_logic_vector(to_unsigned(2,8) ,
35055	 => std_logic_vector(to_unsigned(3,8) ,
35056	 => std_logic_vector(to_unsigned(4,8) ,
35057	 => std_logic_vector(to_unsigned(8,8) ,
35058	 => std_logic_vector(to_unsigned(6,8) ,
35059	 => std_logic_vector(to_unsigned(4,8) ,
35060	 => std_logic_vector(to_unsigned(1,8) ,
35061	 => std_logic_vector(to_unsigned(1,8) ,
35062	 => std_logic_vector(to_unsigned(4,8) ,
35063	 => std_logic_vector(to_unsigned(4,8) ,
35064	 => std_logic_vector(to_unsigned(2,8) ,
35065	 => std_logic_vector(to_unsigned(2,8) ,
35066	 => std_logic_vector(to_unsigned(1,8) ,
35067	 => std_logic_vector(to_unsigned(4,8) ,
35068	 => std_logic_vector(to_unsigned(8,8) ,
35069	 => std_logic_vector(to_unsigned(2,8) ,
35070	 => std_logic_vector(to_unsigned(0,8) ,
35071	 => std_logic_vector(to_unsigned(0,8) ,
35072	 => std_logic_vector(to_unsigned(0,8) ,
35073	 => std_logic_vector(to_unsigned(0,8) ,
35074	 => std_logic_vector(to_unsigned(1,8) ,
35075	 => std_logic_vector(to_unsigned(1,8) ,
35076	 => std_logic_vector(to_unsigned(0,8) ,
35077	 => std_logic_vector(to_unsigned(0,8) ,
35078	 => std_logic_vector(to_unsigned(1,8) ,
35079	 => std_logic_vector(to_unsigned(0,8) ,
35080	 => std_logic_vector(to_unsigned(0,8) ,
35081	 => std_logic_vector(to_unsigned(0,8) ,
35082	 => std_logic_vector(to_unsigned(0,8) ,
35083	 => std_logic_vector(to_unsigned(0,8) ,
35084	 => std_logic_vector(to_unsigned(0,8) ,
35085	 => std_logic_vector(to_unsigned(0,8) ,
35086	 => std_logic_vector(to_unsigned(0,8) ,
35087	 => std_logic_vector(to_unsigned(1,8) ,
35088	 => std_logic_vector(to_unsigned(1,8) ,
35089	 => std_logic_vector(to_unsigned(2,8) ,
35090	 => std_logic_vector(to_unsigned(1,8) ,
35091	 => std_logic_vector(to_unsigned(1,8) ,
35092	 => std_logic_vector(to_unsigned(2,8) ,
35093	 => std_logic_vector(to_unsigned(14,8) ,
35094	 => std_logic_vector(to_unsigned(62,8) ,
35095	 => std_logic_vector(to_unsigned(133,8) ,
35096	 => std_logic_vector(to_unsigned(183,8) ,
35097	 => std_logic_vector(to_unsigned(173,8) ,
35098	 => std_logic_vector(to_unsigned(161,8) ,
35099	 => std_logic_vector(to_unsigned(151,8) ,
35100	 => std_logic_vector(to_unsigned(151,8) ,
35101	 => std_logic_vector(to_unsigned(156,8) ,
35102	 => std_logic_vector(to_unsigned(157,8) ,
35103	 => std_logic_vector(to_unsigned(157,8) ,
35104	 => std_logic_vector(to_unsigned(152,8) ,
35105	 => std_logic_vector(to_unsigned(161,8) ,
35106	 => std_logic_vector(to_unsigned(77,8) ,
35107	 => std_logic_vector(to_unsigned(9,8) ,
35108	 => std_logic_vector(to_unsigned(0,8) ,
35109	 => std_logic_vector(to_unsigned(1,8) ,
35110	 => std_logic_vector(to_unsigned(8,8) ,
35111	 => std_logic_vector(to_unsigned(12,8) ,
35112	 => std_logic_vector(to_unsigned(12,8) ,
35113	 => std_logic_vector(to_unsigned(14,8) ,
35114	 => std_logic_vector(to_unsigned(17,8) ,
35115	 => std_logic_vector(to_unsigned(4,8) ,
35116	 => std_logic_vector(to_unsigned(2,8) ,
35117	 => std_logic_vector(to_unsigned(4,8) ,
35118	 => std_logic_vector(to_unsigned(3,8) ,
35119	 => std_logic_vector(to_unsigned(7,8) ,
35120	 => std_logic_vector(to_unsigned(107,8) ,
35121	 => std_logic_vector(to_unsigned(163,8) ,
35122	 => std_logic_vector(to_unsigned(144,8) ,
35123	 => std_logic_vector(to_unsigned(159,8) ,
35124	 => std_logic_vector(to_unsigned(34,8) ,
35125	 => std_logic_vector(to_unsigned(2,8) ,
35126	 => std_logic_vector(to_unsigned(24,8) ,
35127	 => std_logic_vector(to_unsigned(144,8) ,
35128	 => std_logic_vector(to_unsigned(156,8) ,
35129	 => std_logic_vector(to_unsigned(151,8) ,
35130	 => std_logic_vector(to_unsigned(156,8) ,
35131	 => std_logic_vector(to_unsigned(156,8) ,
35132	 => std_logic_vector(to_unsigned(161,8) ,
35133	 => std_logic_vector(to_unsigned(51,8) ,
35134	 => std_logic_vector(to_unsigned(5,8) ,
35135	 => std_logic_vector(to_unsigned(3,8) ,
35136	 => std_logic_vector(to_unsigned(4,8) ,
35137	 => std_logic_vector(to_unsigned(4,8) ,
35138	 => std_logic_vector(to_unsigned(4,8) ,
35139	 => std_logic_vector(to_unsigned(7,8) ,
35140	 => std_logic_vector(to_unsigned(5,8) ,
35141	 => std_logic_vector(to_unsigned(47,8) ,
35142	 => std_logic_vector(to_unsigned(62,8) ,
35143	 => std_logic_vector(to_unsigned(8,8) ,
35144	 => std_logic_vector(to_unsigned(6,8) ,
35145	 => std_logic_vector(to_unsigned(6,8) ,
35146	 => std_logic_vector(to_unsigned(23,8) ,
35147	 => std_logic_vector(to_unsigned(31,8) ,
35148	 => std_logic_vector(to_unsigned(4,8) ,
35149	 => std_logic_vector(to_unsigned(46,8) ,
35150	 => std_logic_vector(to_unsigned(85,8) ,
35151	 => std_logic_vector(to_unsigned(77,8) ,
35152	 => std_logic_vector(to_unsigned(95,8) ,
35153	 => std_logic_vector(to_unsigned(27,8) ,
35154	 => std_logic_vector(to_unsigned(5,8) ,
35155	 => std_logic_vector(to_unsigned(9,8) ,
35156	 => std_logic_vector(to_unsigned(11,8) ,
35157	 => std_logic_vector(to_unsigned(6,8) ,
35158	 => std_logic_vector(to_unsigned(2,8) ,
35159	 => std_logic_vector(to_unsigned(3,8) ,
35160	 => std_logic_vector(to_unsigned(8,8) ,
35161	 => std_logic_vector(to_unsigned(23,8) ,
35162	 => std_logic_vector(to_unsigned(34,8) ,
35163	 => std_logic_vector(to_unsigned(32,8) ,
35164	 => std_logic_vector(to_unsigned(12,8) ,
35165	 => std_logic_vector(to_unsigned(2,8) ,
35166	 => std_logic_vector(to_unsigned(4,8) ,
35167	 => std_logic_vector(to_unsigned(2,8) ,
35168	 => std_logic_vector(to_unsigned(33,8) ,
35169	 => std_logic_vector(to_unsigned(139,8) ,
35170	 => std_logic_vector(to_unsigned(121,8) ,
35171	 => std_logic_vector(to_unsigned(78,8) ,
35172	 => std_logic_vector(to_unsigned(28,8) ,
35173	 => std_logic_vector(to_unsigned(23,8) ,
35174	 => std_logic_vector(to_unsigned(92,8) ,
35175	 => std_logic_vector(to_unsigned(141,8) ,
35176	 => std_logic_vector(to_unsigned(122,8) ,
35177	 => std_logic_vector(to_unsigned(80,8) ,
35178	 => std_logic_vector(to_unsigned(103,8) ,
35179	 => std_logic_vector(to_unsigned(34,8) ,
35180	 => std_logic_vector(to_unsigned(11,8) ,
35181	 => std_logic_vector(to_unsigned(97,8) ,
35182	 => std_logic_vector(to_unsigned(124,8) ,
35183	 => std_logic_vector(to_unsigned(111,8) ,
35184	 => std_logic_vector(to_unsigned(34,8) ,
35185	 => std_logic_vector(to_unsigned(13,8) ,
35186	 => std_logic_vector(to_unsigned(59,8) ,
35187	 => std_logic_vector(to_unsigned(125,8) ,
35188	 => std_logic_vector(to_unsigned(131,8) ,
35189	 => std_logic_vector(to_unsigned(136,8) ,
35190	 => std_logic_vector(to_unsigned(146,8) ,
35191	 => std_logic_vector(to_unsigned(138,8) ,
35192	 => std_logic_vector(to_unsigned(134,8) ,
35193	 => std_logic_vector(to_unsigned(133,8) ,
35194	 => std_logic_vector(to_unsigned(127,8) ,
35195	 => std_logic_vector(to_unsigned(128,8) ,
35196	 => std_logic_vector(to_unsigned(138,8) ,
35197	 => std_logic_vector(to_unsigned(138,8) ,
35198	 => std_logic_vector(to_unsigned(122,8) ,
35199	 => std_logic_vector(to_unsigned(115,8) ,
35200	 => std_logic_vector(to_unsigned(107,8) ,
35201	 => std_logic_vector(to_unsigned(9,8) ,
35202	 => std_logic_vector(to_unsigned(8,8) ,
35203	 => std_logic_vector(to_unsigned(7,8) ,
35204	 => std_logic_vector(to_unsigned(6,8) ,
35205	 => std_logic_vector(to_unsigned(6,8) ,
35206	 => std_logic_vector(to_unsigned(6,8) ,
35207	 => std_logic_vector(to_unsigned(5,8) ,
35208	 => std_logic_vector(to_unsigned(6,8) ,
35209	 => std_logic_vector(to_unsigned(6,8) ,
35210	 => std_logic_vector(to_unsigned(3,8) ,
35211	 => std_logic_vector(to_unsigned(2,8) ,
35212	 => std_logic_vector(to_unsigned(1,8) ,
35213	 => std_logic_vector(to_unsigned(1,8) ,
35214	 => std_logic_vector(to_unsigned(1,8) ,
35215	 => std_logic_vector(to_unsigned(1,8) ,
35216	 => std_logic_vector(to_unsigned(1,8) ,
35217	 => std_logic_vector(to_unsigned(0,8) ,
35218	 => std_logic_vector(to_unsigned(1,8) ,
35219	 => std_logic_vector(to_unsigned(1,8) ,
35220	 => std_logic_vector(to_unsigned(0,8) ,
35221	 => std_logic_vector(to_unsigned(0,8) ,
35222	 => std_logic_vector(to_unsigned(0,8) ,
35223	 => std_logic_vector(to_unsigned(0,8) ,
35224	 => std_logic_vector(to_unsigned(0,8) ,
35225	 => std_logic_vector(to_unsigned(0,8) ,
35226	 => std_logic_vector(to_unsigned(0,8) ,
35227	 => std_logic_vector(to_unsigned(0,8) ,
35228	 => std_logic_vector(to_unsigned(0,8) ,
35229	 => std_logic_vector(to_unsigned(1,8) ,
35230	 => std_logic_vector(to_unsigned(13,8) ,
35231	 => std_logic_vector(to_unsigned(12,8) ,
35232	 => std_logic_vector(to_unsigned(7,8) ,
35233	 => std_logic_vector(to_unsigned(25,8) ,
35234	 => std_logic_vector(to_unsigned(30,8) ,
35235	 => std_logic_vector(to_unsigned(21,8) ,
35236	 => std_logic_vector(to_unsigned(29,8) ,
35237	 => std_logic_vector(to_unsigned(23,8) ,
35238	 => std_logic_vector(to_unsigned(10,8) ,
35239	 => std_logic_vector(to_unsigned(14,8) ,
35240	 => std_logic_vector(to_unsigned(8,8) ,
35241	 => std_logic_vector(to_unsigned(3,8) ,
35242	 => std_logic_vector(to_unsigned(3,8) ,
35243	 => std_logic_vector(to_unsigned(3,8) ,
35244	 => std_logic_vector(to_unsigned(4,8) ,
35245	 => std_logic_vector(to_unsigned(4,8) ,
35246	 => std_logic_vector(to_unsigned(1,8) ,
35247	 => std_logic_vector(to_unsigned(0,8) ,
35248	 => std_logic_vector(to_unsigned(1,8) ,
35249	 => std_logic_vector(to_unsigned(1,8) ,
35250	 => std_logic_vector(to_unsigned(1,8) ,
35251	 => std_logic_vector(to_unsigned(1,8) ,
35252	 => std_logic_vector(to_unsigned(1,8) ,
35253	 => std_logic_vector(to_unsigned(2,8) ,
35254	 => std_logic_vector(to_unsigned(3,8) ,
35255	 => std_logic_vector(to_unsigned(10,8) ,
35256	 => std_logic_vector(to_unsigned(10,8) ,
35257	 => std_logic_vector(to_unsigned(10,8) ,
35258	 => std_logic_vector(to_unsigned(8,8) ,
35259	 => std_logic_vector(to_unsigned(4,8) ,
35260	 => std_logic_vector(to_unsigned(5,8) ,
35261	 => std_logic_vector(to_unsigned(9,8) ,
35262	 => std_logic_vector(to_unsigned(9,8) ,
35263	 => std_logic_vector(to_unsigned(8,8) ,
35264	 => std_logic_vector(to_unsigned(5,8) ,
35265	 => std_logic_vector(to_unsigned(3,8) ,
35266	 => std_logic_vector(to_unsigned(2,8) ,
35267	 => std_logic_vector(to_unsigned(1,8) ,
35268	 => std_logic_vector(to_unsigned(1,8) ,
35269	 => std_logic_vector(to_unsigned(2,8) ,
35270	 => std_logic_vector(to_unsigned(5,8) ,
35271	 => std_logic_vector(to_unsigned(6,8) ,
35272	 => std_logic_vector(to_unsigned(7,8) ,
35273	 => std_logic_vector(to_unsigned(8,8) ,
35274	 => std_logic_vector(to_unsigned(12,8) ,
35275	 => std_logic_vector(to_unsigned(7,8) ,
35276	 => std_logic_vector(to_unsigned(0,8) ,
35277	 => std_logic_vector(to_unsigned(4,8) ,
35278	 => std_logic_vector(to_unsigned(9,8) ,
35279	 => std_logic_vector(to_unsigned(4,8) ,
35280	 => std_logic_vector(to_unsigned(6,8) ,
35281	 => std_logic_vector(to_unsigned(6,8) ,
35282	 => std_logic_vector(to_unsigned(5,8) ,
35283	 => std_logic_vector(to_unsigned(3,8) ,
35284	 => std_logic_vector(to_unsigned(2,8) ,
35285	 => std_logic_vector(to_unsigned(3,8) ,
35286	 => std_logic_vector(to_unsigned(3,8) ,
35287	 => std_logic_vector(to_unsigned(0,8) ,
35288	 => std_logic_vector(to_unsigned(0,8) ,
35289	 => std_logic_vector(to_unsigned(0,8) ,
35290	 => std_logic_vector(to_unsigned(0,8) ,
35291	 => std_logic_vector(to_unsigned(3,8) ,
35292	 => std_logic_vector(to_unsigned(9,8) ,
35293	 => std_logic_vector(to_unsigned(16,8) ,
35294	 => std_logic_vector(to_unsigned(10,8) ,
35295	 => std_logic_vector(to_unsigned(9,8) ,
35296	 => std_logic_vector(to_unsigned(11,8) ,
35297	 => std_logic_vector(to_unsigned(7,8) ,
35298	 => std_logic_vector(to_unsigned(5,8) ,
35299	 => std_logic_vector(to_unsigned(8,8) ,
35300	 => std_logic_vector(to_unsigned(11,8) ,
35301	 => std_logic_vector(to_unsigned(9,8) ,
35302	 => std_logic_vector(to_unsigned(8,8) ,
35303	 => std_logic_vector(to_unsigned(12,8) ,
35304	 => std_logic_vector(to_unsigned(17,8) ,
35305	 => std_logic_vector(to_unsigned(12,8) ,
35306	 => std_logic_vector(to_unsigned(10,8) ,
35307	 => std_logic_vector(to_unsigned(46,8) ,
35308	 => std_logic_vector(to_unsigned(62,8) ,
35309	 => std_logic_vector(to_unsigned(15,8) ,
35310	 => std_logic_vector(to_unsigned(3,8) ,
35311	 => std_logic_vector(to_unsigned(1,8) ,
35312	 => std_logic_vector(to_unsigned(0,8) ,
35313	 => std_logic_vector(to_unsigned(1,8) ,
35314	 => std_logic_vector(to_unsigned(1,8) ,
35315	 => std_logic_vector(to_unsigned(0,8) ,
35316	 => std_logic_vector(to_unsigned(0,8) ,
35317	 => std_logic_vector(to_unsigned(1,8) ,
35318	 => std_logic_vector(to_unsigned(1,8) ,
35319	 => std_logic_vector(to_unsigned(0,8) ,
35320	 => std_logic_vector(to_unsigned(0,8) ,
35321	 => std_logic_vector(to_unsigned(1,8) ,
35322	 => std_logic_vector(to_unsigned(5,8) ,
35323	 => std_logic_vector(to_unsigned(8,8) ,
35324	 => std_logic_vector(to_unsigned(6,8) ,
35325	 => std_logic_vector(to_unsigned(13,8) ,
35326	 => std_logic_vector(to_unsigned(12,8) ,
35327	 => std_logic_vector(to_unsigned(5,8) ,
35328	 => std_logic_vector(to_unsigned(4,8) ,
35329	 => std_logic_vector(to_unsigned(2,8) ,
35330	 => std_logic_vector(to_unsigned(1,8) ,
35331	 => std_logic_vector(to_unsigned(3,8) ,
35332	 => std_logic_vector(to_unsigned(6,8) ,
35333	 => std_logic_vector(to_unsigned(4,8) ,
35334	 => std_logic_vector(to_unsigned(3,8) ,
35335	 => std_logic_vector(to_unsigned(2,8) ,
35336	 => std_logic_vector(to_unsigned(2,8) ,
35337	 => std_logic_vector(to_unsigned(2,8) ,
35338	 => std_logic_vector(to_unsigned(2,8) ,
35339	 => std_logic_vector(to_unsigned(3,8) ,
35340	 => std_logic_vector(to_unsigned(2,8) ,
35341	 => std_logic_vector(to_unsigned(0,8) ,
35342	 => std_logic_vector(to_unsigned(0,8) ,
35343	 => std_logic_vector(to_unsigned(0,8) ,
35344	 => std_logic_vector(to_unsigned(0,8) ,
35345	 => std_logic_vector(to_unsigned(0,8) ,
35346	 => std_logic_vector(to_unsigned(0,8) ,
35347	 => std_logic_vector(to_unsigned(1,8) ,
35348	 => std_logic_vector(to_unsigned(1,8) ,
35349	 => std_logic_vector(to_unsigned(2,8) ,
35350	 => std_logic_vector(to_unsigned(2,8) ,
35351	 => std_logic_vector(to_unsigned(1,8) ,
35352	 => std_logic_vector(to_unsigned(2,8) ,
35353	 => std_logic_vector(to_unsigned(4,8) ,
35354	 => std_logic_vector(to_unsigned(6,8) ,
35355	 => std_logic_vector(to_unsigned(10,8) ,
35356	 => std_logic_vector(to_unsigned(7,8) ,
35357	 => std_logic_vector(to_unsigned(3,8) ,
35358	 => std_logic_vector(to_unsigned(3,8) ,
35359	 => std_logic_vector(to_unsigned(7,8) ,
35360	 => std_logic_vector(to_unsigned(12,8) ,
35361	 => std_logic_vector(to_unsigned(7,8) ,
35362	 => std_logic_vector(to_unsigned(5,8) ,
35363	 => std_logic_vector(to_unsigned(8,8) ,
35364	 => std_logic_vector(to_unsigned(6,8) ,
35365	 => std_logic_vector(to_unsigned(6,8) ,
35366	 => std_logic_vector(to_unsigned(5,8) ,
35367	 => std_logic_vector(to_unsigned(1,8) ,
35368	 => std_logic_vector(to_unsigned(1,8) ,
35369	 => std_logic_vector(to_unsigned(3,8) ,
35370	 => std_logic_vector(to_unsigned(6,8) ,
35371	 => std_logic_vector(to_unsigned(8,8) ,
35372	 => std_logic_vector(to_unsigned(5,8) ,
35373	 => std_logic_vector(to_unsigned(4,8) ,
35374	 => std_logic_vector(to_unsigned(3,8) ,
35375	 => std_logic_vector(to_unsigned(2,8) ,
35376	 => std_logic_vector(to_unsigned(2,8) ,
35377	 => std_logic_vector(to_unsigned(6,8) ,
35378	 => std_logic_vector(to_unsigned(5,8) ,
35379	 => std_logic_vector(to_unsigned(4,8) ,
35380	 => std_logic_vector(to_unsigned(3,8) ,
35381	 => std_logic_vector(to_unsigned(1,8) ,
35382	 => std_logic_vector(to_unsigned(3,8) ,
35383	 => std_logic_vector(to_unsigned(4,8) ,
35384	 => std_logic_vector(to_unsigned(3,8) ,
35385	 => std_logic_vector(to_unsigned(2,8) ,
35386	 => std_logic_vector(to_unsigned(1,8) ,
35387	 => std_logic_vector(to_unsigned(1,8) ,
35388	 => std_logic_vector(to_unsigned(1,8) ,
35389	 => std_logic_vector(to_unsigned(0,8) ,
35390	 => std_logic_vector(to_unsigned(0,8) ,
35391	 => std_logic_vector(to_unsigned(1,8) ,
35392	 => std_logic_vector(to_unsigned(1,8) ,
35393	 => std_logic_vector(to_unsigned(0,8) ,
35394	 => std_logic_vector(to_unsigned(0,8) ,
35395	 => std_logic_vector(to_unsigned(0,8) ,
35396	 => std_logic_vector(to_unsigned(0,8) ,
35397	 => std_logic_vector(to_unsigned(0,8) ,
35398	 => std_logic_vector(to_unsigned(0,8) ,
35399	 => std_logic_vector(to_unsigned(0,8) ,
35400	 => std_logic_vector(to_unsigned(0,8) ,
35401	 => std_logic_vector(to_unsigned(0,8) ,
35402	 => std_logic_vector(to_unsigned(0,8) ,
35403	 => std_logic_vector(to_unsigned(0,8) ,
35404	 => std_logic_vector(to_unsigned(0,8) ,
35405	 => std_logic_vector(to_unsigned(0,8) ,
35406	 => std_logic_vector(to_unsigned(0,8) ,
35407	 => std_logic_vector(to_unsigned(1,8) ,
35408	 => std_logic_vector(to_unsigned(1,8) ,
35409	 => std_logic_vector(to_unsigned(2,8) ,
35410	 => std_logic_vector(to_unsigned(3,8) ,
35411	 => std_logic_vector(to_unsigned(2,8) ,
35412	 => std_logic_vector(to_unsigned(1,8) ,
35413	 => std_logic_vector(to_unsigned(0,8) ,
35414	 => std_logic_vector(to_unsigned(2,8) ,
35415	 => std_logic_vector(to_unsigned(8,8) ,
35416	 => std_logic_vector(to_unsigned(45,8) ,
35417	 => std_logic_vector(to_unsigned(112,8) ,
35418	 => std_logic_vector(to_unsigned(163,8) ,
35419	 => std_logic_vector(to_unsigned(175,8) ,
35420	 => std_logic_vector(to_unsigned(170,8) ,
35421	 => std_logic_vector(to_unsigned(157,8) ,
35422	 => std_logic_vector(to_unsigned(149,8) ,
35423	 => std_logic_vector(to_unsigned(152,8) ,
35424	 => std_logic_vector(to_unsigned(159,8) ,
35425	 => std_logic_vector(to_unsigned(138,8) ,
35426	 => std_logic_vector(to_unsigned(72,8) ,
35427	 => std_logic_vector(to_unsigned(18,8) ,
35428	 => std_logic_vector(to_unsigned(0,8) ,
35429	 => std_logic_vector(to_unsigned(4,8) ,
35430	 => std_logic_vector(to_unsigned(31,8) ,
35431	 => std_logic_vector(to_unsigned(31,8) ,
35432	 => std_logic_vector(to_unsigned(20,8) ,
35433	 => std_logic_vector(to_unsigned(28,8) ,
35434	 => std_logic_vector(to_unsigned(29,8) ,
35435	 => std_logic_vector(to_unsigned(9,8) ,
35436	 => std_logic_vector(to_unsigned(2,8) ,
35437	 => std_logic_vector(to_unsigned(1,8) ,
35438	 => std_logic_vector(to_unsigned(8,8) ,
35439	 => std_logic_vector(to_unsigned(87,8) ,
35440	 => std_logic_vector(to_unsigned(151,8) ,
35441	 => std_logic_vector(to_unsigned(142,8) ,
35442	 => std_logic_vector(to_unsigned(144,8) ,
35443	 => std_logic_vector(to_unsigned(149,8) ,
35444	 => std_logic_vector(to_unsigned(29,8) ,
35445	 => std_logic_vector(to_unsigned(2,8) ,
35446	 => std_logic_vector(to_unsigned(30,8) ,
35447	 => std_logic_vector(to_unsigned(146,8) ,
35448	 => std_logic_vector(to_unsigned(147,8) ,
35449	 => std_logic_vector(to_unsigned(149,8) ,
35450	 => std_logic_vector(to_unsigned(149,8) ,
35451	 => std_logic_vector(to_unsigned(159,8) ,
35452	 => std_logic_vector(to_unsigned(156,8) ,
35453	 => std_logic_vector(to_unsigned(25,8) ,
35454	 => std_logic_vector(to_unsigned(3,8) ,
35455	 => std_logic_vector(to_unsigned(9,8) ,
35456	 => std_logic_vector(to_unsigned(5,8) ,
35457	 => std_logic_vector(to_unsigned(4,8) ,
35458	 => std_logic_vector(to_unsigned(5,8) ,
35459	 => std_logic_vector(to_unsigned(2,8) ,
35460	 => std_logic_vector(to_unsigned(4,8) ,
35461	 => std_logic_vector(to_unsigned(34,8) ,
35462	 => std_logic_vector(to_unsigned(49,8) ,
35463	 => std_logic_vector(to_unsigned(23,8) ,
35464	 => std_logic_vector(to_unsigned(7,8) ,
35465	 => std_logic_vector(to_unsigned(5,8) ,
35466	 => std_logic_vector(to_unsigned(19,8) ,
35467	 => std_logic_vector(to_unsigned(54,8) ,
35468	 => std_logic_vector(to_unsigned(20,8) ,
35469	 => std_logic_vector(to_unsigned(31,8) ,
35470	 => std_logic_vector(to_unsigned(69,8) ,
35471	 => std_logic_vector(to_unsigned(78,8) ,
35472	 => std_logic_vector(to_unsigned(96,8) ,
35473	 => std_logic_vector(to_unsigned(76,8) ,
35474	 => std_logic_vector(to_unsigned(51,8) ,
35475	 => std_logic_vector(to_unsigned(9,8) ,
35476	 => std_logic_vector(to_unsigned(7,8) ,
35477	 => std_logic_vector(to_unsigned(14,8) ,
35478	 => std_logic_vector(to_unsigned(6,8) ,
35479	 => std_logic_vector(to_unsigned(1,8) ,
35480	 => std_logic_vector(to_unsigned(1,8) ,
35481	 => std_logic_vector(to_unsigned(11,8) ,
35482	 => std_logic_vector(to_unsigned(20,8) ,
35483	 => std_logic_vector(to_unsigned(17,8) ,
35484	 => std_logic_vector(to_unsigned(9,8) ,
35485	 => std_logic_vector(to_unsigned(4,8) ,
35486	 => std_logic_vector(to_unsigned(5,8) ,
35487	 => std_logic_vector(to_unsigned(7,8) ,
35488	 => std_logic_vector(to_unsigned(29,8) ,
35489	 => std_logic_vector(to_unsigned(41,8) ,
35490	 => std_logic_vector(to_unsigned(23,8) ,
35491	 => std_logic_vector(to_unsigned(29,8) ,
35492	 => std_logic_vector(to_unsigned(33,8) ,
35493	 => std_logic_vector(to_unsigned(33,8) ,
35494	 => std_logic_vector(to_unsigned(93,8) ,
35495	 => std_logic_vector(to_unsigned(119,8) ,
35496	 => std_logic_vector(to_unsigned(108,8) ,
35497	 => std_logic_vector(to_unsigned(58,8) ,
35498	 => std_logic_vector(to_unsigned(30,8) ,
35499	 => std_logic_vector(to_unsigned(2,8) ,
35500	 => std_logic_vector(to_unsigned(1,8) ,
35501	 => std_logic_vector(to_unsigned(87,8) ,
35502	 => std_logic_vector(to_unsigned(151,8) ,
35503	 => std_logic_vector(to_unsigned(115,8) ,
35504	 => std_logic_vector(to_unsigned(124,8) ,
35505	 => std_logic_vector(to_unsigned(118,8) ,
35506	 => std_logic_vector(to_unsigned(142,8) ,
35507	 => std_logic_vector(to_unsigned(146,8) ,
35508	 => std_logic_vector(to_unsigned(149,8) ,
35509	 => std_logic_vector(to_unsigned(147,8) ,
35510	 => std_logic_vector(to_unsigned(134,8) ,
35511	 => std_logic_vector(to_unsigned(124,8) ,
35512	 => std_logic_vector(to_unsigned(134,8) ,
35513	 => std_logic_vector(to_unsigned(128,8) ,
35514	 => std_logic_vector(to_unsigned(124,8) ,
35515	 => std_logic_vector(to_unsigned(127,8) ,
35516	 => std_logic_vector(to_unsigned(124,8) ,
35517	 => std_logic_vector(to_unsigned(121,8) ,
35518	 => std_logic_vector(to_unsigned(112,8) ,
35519	 => std_logic_vector(to_unsigned(116,8) ,
35520	 => std_logic_vector(to_unsigned(115,8) ,
35521	 => std_logic_vector(to_unsigned(12,8) ,
35522	 => std_logic_vector(to_unsigned(10,8) ,
35523	 => std_logic_vector(to_unsigned(10,8) ,
35524	 => std_logic_vector(to_unsigned(8,8) ,
35525	 => std_logic_vector(to_unsigned(5,8) ,
35526	 => std_logic_vector(to_unsigned(6,8) ,
35527	 => std_logic_vector(to_unsigned(6,8) ,
35528	 => std_logic_vector(to_unsigned(7,8) ,
35529	 => std_logic_vector(to_unsigned(11,8) ,
35530	 => std_logic_vector(to_unsigned(3,8) ,
35531	 => std_logic_vector(to_unsigned(2,8) ,
35532	 => std_logic_vector(to_unsigned(2,8) ,
35533	 => std_logic_vector(to_unsigned(1,8) ,
35534	 => std_logic_vector(to_unsigned(1,8) ,
35535	 => std_logic_vector(to_unsigned(1,8) ,
35536	 => std_logic_vector(to_unsigned(1,8) ,
35537	 => std_logic_vector(to_unsigned(1,8) ,
35538	 => std_logic_vector(to_unsigned(1,8) ,
35539	 => std_logic_vector(to_unsigned(1,8) ,
35540	 => std_logic_vector(to_unsigned(0,8) ,
35541	 => std_logic_vector(to_unsigned(0,8) ,
35542	 => std_logic_vector(to_unsigned(0,8) ,
35543	 => std_logic_vector(to_unsigned(0,8) ,
35544	 => std_logic_vector(to_unsigned(0,8) ,
35545	 => std_logic_vector(to_unsigned(0,8) ,
35546	 => std_logic_vector(to_unsigned(0,8) ,
35547	 => std_logic_vector(to_unsigned(0,8) ,
35548	 => std_logic_vector(to_unsigned(0,8) ,
35549	 => std_logic_vector(to_unsigned(0,8) ,
35550	 => std_logic_vector(to_unsigned(5,8) ,
35551	 => std_logic_vector(to_unsigned(8,8) ,
35552	 => std_logic_vector(to_unsigned(12,8) ,
35553	 => std_logic_vector(to_unsigned(27,8) ,
35554	 => std_logic_vector(to_unsigned(26,8) ,
35555	 => std_logic_vector(to_unsigned(19,8) ,
35556	 => std_logic_vector(to_unsigned(18,8) ,
35557	 => std_logic_vector(to_unsigned(10,8) ,
35558	 => std_logic_vector(to_unsigned(5,8) ,
35559	 => std_logic_vector(to_unsigned(8,8) ,
35560	 => std_logic_vector(to_unsigned(4,8) ,
35561	 => std_logic_vector(to_unsigned(2,8) ,
35562	 => std_logic_vector(to_unsigned(2,8) ,
35563	 => std_logic_vector(to_unsigned(2,8) ,
35564	 => std_logic_vector(to_unsigned(2,8) ,
35565	 => std_logic_vector(to_unsigned(2,8) ,
35566	 => std_logic_vector(to_unsigned(0,8) ,
35567	 => std_logic_vector(to_unsigned(0,8) ,
35568	 => std_logic_vector(to_unsigned(0,8) ,
35569	 => std_logic_vector(to_unsigned(1,8) ,
35570	 => std_logic_vector(to_unsigned(2,8) ,
35571	 => std_logic_vector(to_unsigned(2,8) ,
35572	 => std_logic_vector(to_unsigned(1,8) ,
35573	 => std_logic_vector(to_unsigned(2,8) ,
35574	 => std_logic_vector(to_unsigned(3,8) ,
35575	 => std_logic_vector(to_unsigned(12,8) ,
35576	 => std_logic_vector(to_unsigned(13,8) ,
35577	 => std_logic_vector(to_unsigned(10,8) ,
35578	 => std_logic_vector(to_unsigned(8,8) ,
35579	 => std_logic_vector(to_unsigned(7,8) ,
35580	 => std_logic_vector(to_unsigned(6,8) ,
35581	 => std_logic_vector(to_unsigned(4,8) ,
35582	 => std_logic_vector(to_unsigned(4,8) ,
35583	 => std_logic_vector(to_unsigned(7,8) ,
35584	 => std_logic_vector(to_unsigned(4,8) ,
35585	 => std_logic_vector(to_unsigned(3,8) ,
35586	 => std_logic_vector(to_unsigned(2,8) ,
35587	 => std_logic_vector(to_unsigned(1,8) ,
35588	 => std_logic_vector(to_unsigned(2,8) ,
35589	 => std_logic_vector(to_unsigned(5,8) ,
35590	 => std_logic_vector(to_unsigned(2,8) ,
35591	 => std_logic_vector(to_unsigned(5,8) ,
35592	 => std_logic_vector(to_unsigned(9,8) ,
35593	 => std_logic_vector(to_unsigned(8,8) ,
35594	 => std_logic_vector(to_unsigned(11,8) ,
35595	 => std_logic_vector(to_unsigned(3,8) ,
35596	 => std_logic_vector(to_unsigned(0,8) ,
35597	 => std_logic_vector(to_unsigned(5,8) ,
35598	 => std_logic_vector(to_unsigned(9,8) ,
35599	 => std_logic_vector(to_unsigned(5,8) ,
35600	 => std_logic_vector(to_unsigned(6,8) ,
35601	 => std_logic_vector(to_unsigned(6,8) ,
35602	 => std_logic_vector(to_unsigned(6,8) ,
35603	 => std_logic_vector(to_unsigned(5,8) ,
35604	 => std_logic_vector(to_unsigned(4,8) ,
35605	 => std_logic_vector(to_unsigned(3,8) ,
35606	 => std_logic_vector(to_unsigned(3,8) ,
35607	 => std_logic_vector(to_unsigned(1,8) ,
35608	 => std_logic_vector(to_unsigned(0,8) ,
35609	 => std_logic_vector(to_unsigned(0,8) ,
35610	 => std_logic_vector(to_unsigned(0,8) ,
35611	 => std_logic_vector(to_unsigned(3,8) ,
35612	 => std_logic_vector(to_unsigned(9,8) ,
35613	 => std_logic_vector(to_unsigned(12,8) ,
35614	 => std_logic_vector(to_unsigned(11,8) ,
35615	 => std_logic_vector(to_unsigned(13,8) ,
35616	 => std_logic_vector(to_unsigned(9,8) ,
35617	 => std_logic_vector(to_unsigned(7,8) ,
35618	 => std_logic_vector(to_unsigned(4,8) ,
35619	 => std_logic_vector(to_unsigned(6,8) ,
35620	 => std_logic_vector(to_unsigned(13,8) ,
35621	 => std_logic_vector(to_unsigned(10,8) ,
35622	 => std_logic_vector(to_unsigned(7,8) ,
35623	 => std_logic_vector(to_unsigned(4,8) ,
35624	 => std_logic_vector(to_unsigned(2,8) ,
35625	 => std_logic_vector(to_unsigned(1,8) ,
35626	 => std_logic_vector(to_unsigned(2,8) ,
35627	 => std_logic_vector(to_unsigned(28,8) ,
35628	 => std_logic_vector(to_unsigned(29,8) ,
35629	 => std_logic_vector(to_unsigned(12,8) ,
35630	 => std_logic_vector(to_unsigned(7,8) ,
35631	 => std_logic_vector(to_unsigned(4,8) ,
35632	 => std_logic_vector(to_unsigned(11,8) ,
35633	 => std_logic_vector(to_unsigned(3,8) ,
35634	 => std_logic_vector(to_unsigned(1,8) ,
35635	 => std_logic_vector(to_unsigned(0,8) ,
35636	 => std_logic_vector(to_unsigned(0,8) ,
35637	 => std_logic_vector(to_unsigned(1,8) ,
35638	 => std_logic_vector(to_unsigned(0,8) ,
35639	 => std_logic_vector(to_unsigned(0,8) ,
35640	 => std_logic_vector(to_unsigned(1,8) ,
35641	 => std_logic_vector(to_unsigned(1,8) ,
35642	 => std_logic_vector(to_unsigned(6,8) ,
35643	 => std_logic_vector(to_unsigned(8,8) ,
35644	 => std_logic_vector(to_unsigned(7,8) ,
35645	 => std_logic_vector(to_unsigned(14,8) ,
35646	 => std_logic_vector(to_unsigned(13,8) ,
35647	 => std_logic_vector(to_unsigned(5,8) ,
35648	 => std_logic_vector(to_unsigned(3,8) ,
35649	 => std_logic_vector(to_unsigned(2,8) ,
35650	 => std_logic_vector(to_unsigned(1,8) ,
35651	 => std_logic_vector(to_unsigned(2,8) ,
35652	 => std_logic_vector(to_unsigned(5,8) ,
35653	 => std_logic_vector(to_unsigned(4,8) ,
35654	 => std_logic_vector(to_unsigned(4,8) ,
35655	 => std_logic_vector(to_unsigned(3,8) ,
35656	 => std_logic_vector(to_unsigned(2,8) ,
35657	 => std_logic_vector(to_unsigned(2,8) ,
35658	 => std_logic_vector(to_unsigned(2,8) ,
35659	 => std_logic_vector(to_unsigned(2,8) ,
35660	 => std_logic_vector(to_unsigned(1,8) ,
35661	 => std_logic_vector(to_unsigned(0,8) ,
35662	 => std_logic_vector(to_unsigned(0,8) ,
35663	 => std_logic_vector(to_unsigned(0,8) ,
35664	 => std_logic_vector(to_unsigned(1,8) ,
35665	 => std_logic_vector(to_unsigned(0,8) ,
35666	 => std_logic_vector(to_unsigned(1,8) ,
35667	 => std_logic_vector(to_unsigned(2,8) ,
35668	 => std_logic_vector(to_unsigned(2,8) ,
35669	 => std_logic_vector(to_unsigned(3,8) ,
35670	 => std_logic_vector(to_unsigned(3,8) ,
35671	 => std_logic_vector(to_unsigned(2,8) ,
35672	 => std_logic_vector(to_unsigned(2,8) ,
35673	 => std_logic_vector(to_unsigned(4,8) ,
35674	 => std_logic_vector(to_unsigned(7,8) ,
35675	 => std_logic_vector(to_unsigned(10,8) ,
35676	 => std_logic_vector(to_unsigned(4,8) ,
35677	 => std_logic_vector(to_unsigned(2,8) ,
35678	 => std_logic_vector(to_unsigned(2,8) ,
35679	 => std_logic_vector(to_unsigned(6,8) ,
35680	 => std_logic_vector(to_unsigned(12,8) ,
35681	 => std_logic_vector(to_unsigned(8,8) ,
35682	 => std_logic_vector(to_unsigned(5,8) ,
35683	 => std_logic_vector(to_unsigned(8,8) ,
35684	 => std_logic_vector(to_unsigned(7,8) ,
35685	 => std_logic_vector(to_unsigned(5,8) ,
35686	 => std_logic_vector(to_unsigned(3,8) ,
35687	 => std_logic_vector(to_unsigned(0,8) ,
35688	 => std_logic_vector(to_unsigned(0,8) ,
35689	 => std_logic_vector(to_unsigned(1,8) ,
35690	 => std_logic_vector(to_unsigned(1,8) ,
35691	 => std_logic_vector(to_unsigned(2,8) ,
35692	 => std_logic_vector(to_unsigned(3,8) ,
35693	 => std_logic_vector(to_unsigned(3,8) ,
35694	 => std_logic_vector(to_unsigned(3,8) ,
35695	 => std_logic_vector(to_unsigned(4,8) ,
35696	 => std_logic_vector(to_unsigned(2,8) ,
35697	 => std_logic_vector(to_unsigned(3,8) ,
35698	 => std_logic_vector(to_unsigned(5,8) ,
35699	 => std_logic_vector(to_unsigned(4,8) ,
35700	 => std_logic_vector(to_unsigned(3,8) ,
35701	 => std_logic_vector(to_unsigned(2,8) ,
35702	 => std_logic_vector(to_unsigned(2,8) ,
35703	 => std_logic_vector(to_unsigned(3,8) ,
35704	 => std_logic_vector(to_unsigned(2,8) ,
35705	 => std_logic_vector(to_unsigned(2,8) ,
35706	 => std_logic_vector(to_unsigned(1,8) ,
35707	 => std_logic_vector(to_unsigned(1,8) ,
35708	 => std_logic_vector(to_unsigned(0,8) ,
35709	 => std_logic_vector(to_unsigned(0,8) ,
35710	 => std_logic_vector(to_unsigned(1,8) ,
35711	 => std_logic_vector(to_unsigned(1,8) ,
35712	 => std_logic_vector(to_unsigned(1,8) ,
35713	 => std_logic_vector(to_unsigned(1,8) ,
35714	 => std_logic_vector(to_unsigned(0,8) ,
35715	 => std_logic_vector(to_unsigned(0,8) ,
35716	 => std_logic_vector(to_unsigned(0,8) ,
35717	 => std_logic_vector(to_unsigned(0,8) ,
35718	 => std_logic_vector(to_unsigned(0,8) ,
35719	 => std_logic_vector(to_unsigned(0,8) ,
35720	 => std_logic_vector(to_unsigned(0,8) ,
35721	 => std_logic_vector(to_unsigned(0,8) ,
35722	 => std_logic_vector(to_unsigned(0,8) ,
35723	 => std_logic_vector(to_unsigned(0,8) ,
35724	 => std_logic_vector(to_unsigned(0,8) ,
35725	 => std_logic_vector(to_unsigned(0,8) ,
35726	 => std_logic_vector(to_unsigned(0,8) ,
35727	 => std_logic_vector(to_unsigned(1,8) ,
35728	 => std_logic_vector(to_unsigned(2,8) ,
35729	 => std_logic_vector(to_unsigned(2,8) ,
35730	 => std_logic_vector(to_unsigned(2,8) ,
35731	 => std_logic_vector(to_unsigned(2,8) ,
35732	 => std_logic_vector(to_unsigned(1,8) ,
35733	 => std_logic_vector(to_unsigned(2,8) ,
35734	 => std_logic_vector(to_unsigned(6,8) ,
35735	 => std_logic_vector(to_unsigned(3,8) ,
35736	 => std_logic_vector(to_unsigned(2,8) ,
35737	 => std_logic_vector(to_unsigned(4,8) ,
35738	 => std_logic_vector(to_unsigned(23,8) ,
35739	 => std_logic_vector(to_unsigned(70,8) ,
35740	 => std_logic_vector(to_unsigned(136,8) ,
35741	 => std_logic_vector(to_unsigned(173,8) ,
35742	 => std_logic_vector(to_unsigned(171,8) ,
35743	 => std_logic_vector(to_unsigned(156,8) ,
35744	 => std_logic_vector(to_unsigned(152,8) ,
35745	 => std_logic_vector(to_unsigned(142,8) ,
35746	 => std_logic_vector(to_unsigned(81,8) ,
35747	 => std_logic_vector(to_unsigned(8,8) ,
35748	 => std_logic_vector(to_unsigned(0,8) ,
35749	 => std_logic_vector(to_unsigned(17,8) ,
35750	 => std_logic_vector(to_unsigned(37,8) ,
35751	 => std_logic_vector(to_unsigned(36,8) ,
35752	 => std_logic_vector(to_unsigned(41,8) ,
35753	 => std_logic_vector(to_unsigned(34,8) ,
35754	 => std_logic_vector(to_unsigned(22,8) ,
35755	 => std_logic_vector(to_unsigned(7,8) ,
35756	 => std_logic_vector(to_unsigned(2,8) ,
35757	 => std_logic_vector(to_unsigned(1,8) ,
35758	 => std_logic_vector(to_unsigned(16,8) ,
35759	 => std_logic_vector(to_unsigned(128,8) ,
35760	 => std_logic_vector(to_unsigned(168,8) ,
35761	 => std_logic_vector(to_unsigned(163,8) ,
35762	 => std_logic_vector(to_unsigned(177,8) ,
35763	 => std_logic_vector(to_unsigned(144,8) ,
35764	 => std_logic_vector(to_unsigned(13,8) ,
35765	 => std_logic_vector(to_unsigned(1,8) ,
35766	 => std_logic_vector(to_unsigned(35,8) ,
35767	 => std_logic_vector(to_unsigned(161,8) ,
35768	 => std_logic_vector(to_unsigned(152,8) ,
35769	 => std_logic_vector(to_unsigned(149,8) ,
35770	 => std_logic_vector(to_unsigned(154,8) ,
35771	 => std_logic_vector(to_unsigned(152,8) ,
35772	 => std_logic_vector(to_unsigned(156,8) ,
35773	 => std_logic_vector(to_unsigned(130,8) ,
35774	 => std_logic_vector(to_unsigned(37,8) ,
35775	 => std_logic_vector(to_unsigned(5,8) ,
35776	 => std_logic_vector(to_unsigned(6,8) ,
35777	 => std_logic_vector(to_unsigned(6,8) ,
35778	 => std_logic_vector(to_unsigned(6,8) ,
35779	 => std_logic_vector(to_unsigned(2,8) ,
35780	 => std_logic_vector(to_unsigned(11,8) ,
35781	 => std_logic_vector(to_unsigned(16,8) ,
35782	 => std_logic_vector(to_unsigned(30,8) ,
35783	 => std_logic_vector(to_unsigned(44,8) ,
35784	 => std_logic_vector(to_unsigned(13,8) ,
35785	 => std_logic_vector(to_unsigned(7,8) ,
35786	 => std_logic_vector(to_unsigned(16,8) ,
35787	 => std_logic_vector(to_unsigned(38,8) ,
35788	 => std_logic_vector(to_unsigned(66,8) ,
35789	 => std_logic_vector(to_unsigned(86,8) ,
35790	 => std_logic_vector(to_unsigned(84,8) ,
35791	 => std_logic_vector(to_unsigned(73,8) ,
35792	 => std_logic_vector(to_unsigned(86,8) ,
35793	 => std_logic_vector(to_unsigned(42,8) ,
35794	 => std_logic_vector(to_unsigned(61,8) ,
35795	 => std_logic_vector(to_unsigned(72,8) ,
35796	 => std_logic_vector(to_unsigned(10,8) ,
35797	 => std_logic_vector(to_unsigned(7,8) ,
35798	 => std_logic_vector(to_unsigned(16,8) ,
35799	 => std_logic_vector(to_unsigned(7,8) ,
35800	 => std_logic_vector(to_unsigned(1,8) ,
35801	 => std_logic_vector(to_unsigned(1,8) ,
35802	 => std_logic_vector(to_unsigned(4,8) ,
35803	 => std_logic_vector(to_unsigned(6,8) ,
35804	 => std_logic_vector(to_unsigned(8,8) ,
35805	 => std_logic_vector(to_unsigned(7,8) ,
35806	 => std_logic_vector(to_unsigned(4,8) ,
35807	 => std_logic_vector(to_unsigned(14,8) ,
35808	 => std_logic_vector(to_unsigned(35,8) ,
35809	 => std_logic_vector(to_unsigned(27,8) ,
35810	 => std_logic_vector(to_unsigned(13,8) ,
35811	 => std_logic_vector(to_unsigned(23,8) ,
35812	 => std_logic_vector(to_unsigned(46,8) ,
35813	 => std_logic_vector(to_unsigned(38,8) ,
35814	 => std_logic_vector(to_unsigned(59,8) ,
35815	 => std_logic_vector(to_unsigned(93,8) ,
35816	 => std_logic_vector(to_unsigned(77,8) ,
35817	 => std_logic_vector(to_unsigned(11,8) ,
35818	 => std_logic_vector(to_unsigned(2,8) ,
35819	 => std_logic_vector(to_unsigned(1,8) ,
35820	 => std_logic_vector(to_unsigned(2,8) ,
35821	 => std_logic_vector(to_unsigned(85,8) ,
35822	 => std_logic_vector(to_unsigned(154,8) ,
35823	 => std_logic_vector(to_unsigned(116,8) ,
35824	 => std_logic_vector(to_unsigned(124,8) ,
35825	 => std_logic_vector(to_unsigned(154,8) ,
35826	 => std_logic_vector(to_unsigned(171,8) ,
35827	 => std_logic_vector(to_unsigned(168,8) ,
35828	 => std_logic_vector(to_unsigned(152,8) ,
35829	 => std_logic_vector(to_unsigned(138,8) ,
35830	 => std_logic_vector(to_unsigned(130,8) ,
35831	 => std_logic_vector(to_unsigned(128,8) ,
35832	 => std_logic_vector(to_unsigned(131,8) ,
35833	 => std_logic_vector(to_unsigned(128,8) ,
35834	 => std_logic_vector(to_unsigned(133,8) ,
35835	 => std_logic_vector(to_unsigned(131,8) ,
35836	 => std_logic_vector(to_unsigned(130,8) ,
35837	 => std_logic_vector(to_unsigned(116,8) ,
35838	 => std_logic_vector(to_unsigned(107,8) ,
35839	 => std_logic_vector(to_unsigned(121,8) ,
35840	 => std_logic_vector(to_unsigned(124,8) ,
35841	 => std_logic_vector(to_unsigned(29,8) ,
35842	 => std_logic_vector(to_unsigned(29,8) ,
35843	 => std_logic_vector(to_unsigned(30,8) ,
35844	 => std_logic_vector(to_unsigned(24,8) ,
35845	 => std_logic_vector(to_unsigned(15,8) ,
35846	 => std_logic_vector(to_unsigned(13,8) ,
35847	 => std_logic_vector(to_unsigned(8,8) ,
35848	 => std_logic_vector(to_unsigned(13,8) ,
35849	 => std_logic_vector(to_unsigned(31,8) ,
35850	 => std_logic_vector(to_unsigned(5,8) ,
35851	 => std_logic_vector(to_unsigned(2,8) ,
35852	 => std_logic_vector(to_unsigned(2,8) ,
35853	 => std_logic_vector(to_unsigned(1,8) ,
35854	 => std_logic_vector(to_unsigned(1,8) ,
35855	 => std_logic_vector(to_unsigned(1,8) ,
35856	 => std_logic_vector(to_unsigned(0,8) ,
35857	 => std_logic_vector(to_unsigned(1,8) ,
35858	 => std_logic_vector(to_unsigned(1,8) ,
35859	 => std_logic_vector(to_unsigned(0,8) ,
35860	 => std_logic_vector(to_unsigned(0,8) ,
35861	 => std_logic_vector(to_unsigned(0,8) ,
35862	 => std_logic_vector(to_unsigned(0,8) ,
35863	 => std_logic_vector(to_unsigned(0,8) ,
35864	 => std_logic_vector(to_unsigned(0,8) ,
35865	 => std_logic_vector(to_unsigned(0,8) ,
35866	 => std_logic_vector(to_unsigned(0,8) ,
35867	 => std_logic_vector(to_unsigned(0,8) ,
35868	 => std_logic_vector(to_unsigned(0,8) ,
35869	 => std_logic_vector(to_unsigned(0,8) ,
35870	 => std_logic_vector(to_unsigned(2,8) ,
35871	 => std_logic_vector(to_unsigned(5,8) ,
35872	 => std_logic_vector(to_unsigned(17,8) ,
35873	 => std_logic_vector(to_unsigned(23,8) ,
35874	 => std_logic_vector(to_unsigned(22,8) ,
35875	 => std_logic_vector(to_unsigned(17,8) ,
35876	 => std_logic_vector(to_unsigned(7,8) ,
35877	 => std_logic_vector(to_unsigned(4,8) ,
35878	 => std_logic_vector(to_unsigned(3,8) ,
35879	 => std_logic_vector(to_unsigned(3,8) ,
35880	 => std_logic_vector(to_unsigned(3,8) ,
35881	 => std_logic_vector(to_unsigned(2,8) ,
35882	 => std_logic_vector(to_unsigned(3,8) ,
35883	 => std_logic_vector(to_unsigned(3,8) ,
35884	 => std_logic_vector(to_unsigned(4,8) ,
35885	 => std_logic_vector(to_unsigned(2,8) ,
35886	 => std_logic_vector(to_unsigned(0,8) ,
35887	 => std_logic_vector(to_unsigned(0,8) ,
35888	 => std_logic_vector(to_unsigned(0,8) ,
35889	 => std_logic_vector(to_unsigned(0,8) ,
35890	 => std_logic_vector(to_unsigned(1,8) ,
35891	 => std_logic_vector(to_unsigned(2,8) ,
35892	 => std_logic_vector(to_unsigned(3,8) ,
35893	 => std_logic_vector(to_unsigned(2,8) ,
35894	 => std_logic_vector(to_unsigned(3,8) ,
35895	 => std_logic_vector(to_unsigned(14,8) ,
35896	 => std_logic_vector(to_unsigned(12,8) ,
35897	 => std_logic_vector(to_unsigned(10,8) ,
35898	 => std_logic_vector(to_unsigned(8,8) ,
35899	 => std_logic_vector(to_unsigned(8,8) ,
35900	 => std_logic_vector(to_unsigned(10,8) ,
35901	 => std_logic_vector(to_unsigned(6,8) ,
35902	 => std_logic_vector(to_unsigned(4,8) ,
35903	 => std_logic_vector(to_unsigned(4,8) ,
35904	 => std_logic_vector(to_unsigned(2,8) ,
35905	 => std_logic_vector(to_unsigned(3,8) ,
35906	 => std_logic_vector(to_unsigned(2,8) ,
35907	 => std_logic_vector(to_unsigned(0,8) ,
35908	 => std_logic_vector(to_unsigned(1,8) ,
35909	 => std_logic_vector(to_unsigned(8,8) ,
35910	 => std_logic_vector(to_unsigned(6,8) ,
35911	 => std_logic_vector(to_unsigned(5,8) ,
35912	 => std_logic_vector(to_unsigned(5,8) ,
35913	 => std_logic_vector(to_unsigned(8,8) ,
35914	 => std_logic_vector(to_unsigned(10,8) ,
35915	 => std_logic_vector(to_unsigned(1,8) ,
35916	 => std_logic_vector(to_unsigned(0,8) ,
35917	 => std_logic_vector(to_unsigned(7,8) ,
35918	 => std_logic_vector(to_unsigned(9,8) ,
35919	 => std_logic_vector(to_unsigned(4,8) ,
35920	 => std_logic_vector(to_unsigned(5,8) ,
35921	 => std_logic_vector(to_unsigned(5,8) ,
35922	 => std_logic_vector(to_unsigned(5,8) ,
35923	 => std_logic_vector(to_unsigned(3,8) ,
35924	 => std_logic_vector(to_unsigned(4,8) ,
35925	 => std_logic_vector(to_unsigned(3,8) ,
35926	 => std_logic_vector(to_unsigned(1,8) ,
35927	 => std_logic_vector(to_unsigned(1,8) ,
35928	 => std_logic_vector(to_unsigned(0,8) ,
35929	 => std_logic_vector(to_unsigned(0,8) ,
35930	 => std_logic_vector(to_unsigned(0,8) ,
35931	 => std_logic_vector(to_unsigned(1,8) ,
35932	 => std_logic_vector(to_unsigned(10,8) ,
35933	 => std_logic_vector(to_unsigned(12,8) ,
35934	 => std_logic_vector(to_unsigned(8,8) ,
35935	 => std_logic_vector(to_unsigned(10,8) ,
35936	 => std_logic_vector(to_unsigned(10,8) ,
35937	 => std_logic_vector(to_unsigned(8,8) ,
35938	 => std_logic_vector(to_unsigned(3,8) ,
35939	 => std_logic_vector(to_unsigned(4,8) ,
35940	 => std_logic_vector(to_unsigned(13,8) ,
35941	 => std_logic_vector(to_unsigned(10,8) ,
35942	 => std_logic_vector(to_unsigned(7,8) ,
35943	 => std_logic_vector(to_unsigned(3,8) ,
35944	 => std_logic_vector(to_unsigned(1,8) ,
35945	 => std_logic_vector(to_unsigned(0,8) ,
35946	 => std_logic_vector(to_unsigned(3,8) ,
35947	 => std_logic_vector(to_unsigned(29,8) ,
35948	 => std_logic_vector(to_unsigned(19,8) ,
35949	 => std_logic_vector(to_unsigned(10,8) ,
35950	 => std_logic_vector(to_unsigned(7,8) ,
35951	 => std_logic_vector(to_unsigned(45,8) ,
35952	 => std_logic_vector(to_unsigned(152,8) ,
35953	 => std_logic_vector(to_unsigned(48,8) ,
35954	 => std_logic_vector(to_unsigned(1,8) ,
35955	 => std_logic_vector(to_unsigned(0,8) ,
35956	 => std_logic_vector(to_unsigned(1,8) ,
35957	 => std_logic_vector(to_unsigned(0,8) ,
35958	 => std_logic_vector(to_unsigned(0,8) ,
35959	 => std_logic_vector(to_unsigned(0,8) ,
35960	 => std_logic_vector(to_unsigned(0,8) ,
35961	 => std_logic_vector(to_unsigned(1,8) ,
35962	 => std_logic_vector(to_unsigned(8,8) ,
35963	 => std_logic_vector(to_unsigned(7,8) ,
35964	 => std_logic_vector(to_unsigned(6,8) ,
35965	 => std_logic_vector(to_unsigned(13,8) ,
35966	 => std_logic_vector(to_unsigned(9,8) ,
35967	 => std_logic_vector(to_unsigned(4,8) ,
35968	 => std_logic_vector(to_unsigned(3,8) ,
35969	 => std_logic_vector(to_unsigned(2,8) ,
35970	 => std_logic_vector(to_unsigned(0,8) ,
35971	 => std_logic_vector(to_unsigned(3,8) ,
35972	 => std_logic_vector(to_unsigned(5,8) ,
35973	 => std_logic_vector(to_unsigned(4,8) ,
35974	 => std_logic_vector(to_unsigned(4,8) ,
35975	 => std_logic_vector(to_unsigned(3,8) ,
35976	 => std_logic_vector(to_unsigned(2,8) ,
35977	 => std_logic_vector(to_unsigned(2,8) ,
35978	 => std_logic_vector(to_unsigned(2,8) ,
35979	 => std_logic_vector(to_unsigned(1,8) ,
35980	 => std_logic_vector(to_unsigned(1,8) ,
35981	 => std_logic_vector(to_unsigned(0,8) ,
35982	 => std_logic_vector(to_unsigned(0,8) ,
35983	 => std_logic_vector(to_unsigned(0,8) ,
35984	 => std_logic_vector(to_unsigned(0,8) ,
35985	 => std_logic_vector(to_unsigned(0,8) ,
35986	 => std_logic_vector(to_unsigned(1,8) ,
35987	 => std_logic_vector(to_unsigned(2,8) ,
35988	 => std_logic_vector(to_unsigned(2,8) ,
35989	 => std_logic_vector(to_unsigned(2,8) ,
35990	 => std_logic_vector(to_unsigned(3,8) ,
35991	 => std_logic_vector(to_unsigned(2,8) ,
35992	 => std_logic_vector(to_unsigned(2,8) ,
35993	 => std_logic_vector(to_unsigned(4,8) ,
35994	 => std_logic_vector(to_unsigned(7,8) ,
35995	 => std_logic_vector(to_unsigned(10,8) ,
35996	 => std_logic_vector(to_unsigned(3,8) ,
35997	 => std_logic_vector(to_unsigned(1,8) ,
35998	 => std_logic_vector(to_unsigned(1,8) ,
35999	 => std_logic_vector(to_unsigned(3,8) ,
36000	 => std_logic_vector(to_unsigned(10,8) ,
36001	 => std_logic_vector(to_unsigned(8,8) ,
36002	 => std_logic_vector(to_unsigned(4,8) ,
36003	 => std_logic_vector(to_unsigned(5,8) ,
36004	 => std_logic_vector(to_unsigned(6,8) ,
36005	 => std_logic_vector(to_unsigned(5,8) ,
36006	 => std_logic_vector(to_unsigned(2,8) ,
36007	 => std_logic_vector(to_unsigned(0,8) ,
36008	 => std_logic_vector(to_unsigned(0,8) ,
36009	 => std_logic_vector(to_unsigned(0,8) ,
36010	 => std_logic_vector(to_unsigned(0,8) ,
36011	 => std_logic_vector(to_unsigned(0,8) ,
36012	 => std_logic_vector(to_unsigned(0,8) ,
36013	 => std_logic_vector(to_unsigned(0,8) ,
36014	 => std_logic_vector(to_unsigned(1,8) ,
36015	 => std_logic_vector(to_unsigned(3,8) ,
36016	 => std_logic_vector(to_unsigned(1,8) ,
36017	 => std_logic_vector(to_unsigned(4,8) ,
36018	 => std_logic_vector(to_unsigned(4,8) ,
36019	 => std_logic_vector(to_unsigned(3,8) ,
36020	 => std_logic_vector(to_unsigned(3,8) ,
36021	 => std_logic_vector(to_unsigned(1,8) ,
36022	 => std_logic_vector(to_unsigned(2,8) ,
36023	 => std_logic_vector(to_unsigned(3,8) ,
36024	 => std_logic_vector(to_unsigned(2,8) ,
36025	 => std_logic_vector(to_unsigned(3,8) ,
36026	 => std_logic_vector(to_unsigned(1,8) ,
36027	 => std_logic_vector(to_unsigned(2,8) ,
36028	 => std_logic_vector(to_unsigned(1,8) ,
36029	 => std_logic_vector(to_unsigned(0,8) ,
36030	 => std_logic_vector(to_unsigned(1,8) ,
36031	 => std_logic_vector(to_unsigned(0,8) ,
36032	 => std_logic_vector(to_unsigned(0,8) ,
36033	 => std_logic_vector(to_unsigned(1,8) ,
36034	 => std_logic_vector(to_unsigned(1,8) ,
36035	 => std_logic_vector(to_unsigned(1,8) ,
36036	 => std_logic_vector(to_unsigned(1,8) ,
36037	 => std_logic_vector(to_unsigned(1,8) ,
36038	 => std_logic_vector(to_unsigned(1,8) ,
36039	 => std_logic_vector(to_unsigned(1,8) ,
36040	 => std_logic_vector(to_unsigned(1,8) ,
36041	 => std_logic_vector(to_unsigned(1,8) ,
36042	 => std_logic_vector(to_unsigned(1,8) ,
36043	 => std_logic_vector(to_unsigned(0,8) ,
36044	 => std_logic_vector(to_unsigned(0,8) ,
36045	 => std_logic_vector(to_unsigned(0,8) ,
36046	 => std_logic_vector(to_unsigned(1,8) ,
36047	 => std_logic_vector(to_unsigned(2,8) ,
36048	 => std_logic_vector(to_unsigned(2,8) ,
36049	 => std_logic_vector(to_unsigned(2,8) ,
36050	 => std_logic_vector(to_unsigned(3,8) ,
36051	 => std_logic_vector(to_unsigned(2,8) ,
36052	 => std_logic_vector(to_unsigned(0,8) ,
36053	 => std_logic_vector(to_unsigned(3,8) ,
36054	 => std_logic_vector(to_unsigned(10,8) ,
36055	 => std_logic_vector(to_unsigned(9,8) ,
36056	 => std_logic_vector(to_unsigned(7,8) ,
36057	 => std_logic_vector(to_unsigned(5,8) ,
36058	 => std_logic_vector(to_unsigned(2,8) ,
36059	 => std_logic_vector(to_unsigned(2,8) ,
36060	 => std_logic_vector(to_unsigned(12,8) ,
36061	 => std_logic_vector(to_unsigned(52,8) ,
36062	 => std_logic_vector(to_unsigned(116,8) ,
36063	 => std_logic_vector(to_unsigned(166,8) ,
36064	 => std_logic_vector(to_unsigned(177,8) ,
36065	 => std_logic_vector(to_unsigned(119,8) ,
36066	 => std_logic_vector(to_unsigned(33,8) ,
36067	 => std_logic_vector(to_unsigned(1,8) ,
36068	 => std_logic_vector(to_unsigned(1,8) ,
36069	 => std_logic_vector(to_unsigned(11,8) ,
36070	 => std_logic_vector(to_unsigned(25,8) ,
36071	 => std_logic_vector(to_unsigned(39,8) ,
36072	 => std_logic_vector(to_unsigned(51,8) ,
36073	 => std_logic_vector(to_unsigned(33,8) ,
36074	 => std_logic_vector(to_unsigned(19,8) ,
36075	 => std_logic_vector(to_unsigned(10,8) ,
36076	 => std_logic_vector(to_unsigned(2,8) ,
36077	 => std_logic_vector(to_unsigned(2,8) ,
36078	 => std_logic_vector(to_unsigned(2,8) ,
36079	 => std_logic_vector(to_unsigned(9,8) ,
36080	 => std_logic_vector(to_unsigned(28,8) ,
36081	 => std_logic_vector(to_unsigned(45,8) ,
36082	 => std_logic_vector(to_unsigned(70,8) ,
36083	 => std_logic_vector(to_unsigned(84,8) ,
36084	 => std_logic_vector(to_unsigned(18,8) ,
36085	 => std_logic_vector(to_unsigned(4,8) ,
36086	 => std_logic_vector(to_unsigned(45,8) ,
36087	 => std_logic_vector(to_unsigned(157,8) ,
36088	 => std_logic_vector(to_unsigned(152,8) ,
36089	 => std_logic_vector(to_unsigned(154,8) ,
36090	 => std_logic_vector(to_unsigned(164,8) ,
36091	 => std_logic_vector(to_unsigned(161,8) ,
36092	 => std_logic_vector(to_unsigned(164,8) ,
36093	 => std_logic_vector(to_unsigned(149,8) ,
36094	 => std_logic_vector(to_unsigned(46,8) ,
36095	 => std_logic_vector(to_unsigned(10,8) ,
36096	 => std_logic_vector(to_unsigned(6,8) ,
36097	 => std_logic_vector(to_unsigned(5,8) ,
36098	 => std_logic_vector(to_unsigned(5,8) ,
36099	 => std_logic_vector(to_unsigned(7,8) ,
36100	 => std_logic_vector(to_unsigned(11,8) ,
36101	 => std_logic_vector(to_unsigned(12,8) ,
36102	 => std_logic_vector(to_unsigned(14,8) ,
36103	 => std_logic_vector(to_unsigned(23,8) ,
36104	 => std_logic_vector(to_unsigned(29,8) ,
36105	 => std_logic_vector(to_unsigned(9,8) ,
36106	 => std_logic_vector(to_unsigned(8,8) ,
36107	 => std_logic_vector(to_unsigned(22,8) ,
36108	 => std_logic_vector(to_unsigned(65,8) ,
36109	 => std_logic_vector(to_unsigned(71,8) ,
36110	 => std_logic_vector(to_unsigned(51,8) ,
36111	 => std_logic_vector(to_unsigned(46,8) ,
36112	 => std_logic_vector(to_unsigned(65,8) ,
36113	 => std_logic_vector(to_unsigned(35,8) ,
36114	 => std_logic_vector(to_unsigned(12,8) ,
36115	 => std_logic_vector(to_unsigned(74,8) ,
36116	 => std_logic_vector(to_unsigned(26,8) ,
36117	 => std_logic_vector(to_unsigned(9,8) ,
36118	 => std_logic_vector(to_unsigned(8,8) ,
36119	 => std_logic_vector(to_unsigned(10,8) ,
36120	 => std_logic_vector(to_unsigned(3,8) ,
36121	 => std_logic_vector(to_unsigned(1,8) ,
36122	 => std_logic_vector(to_unsigned(2,8) ,
36123	 => std_logic_vector(to_unsigned(6,8) ,
36124	 => std_logic_vector(to_unsigned(6,8) ,
36125	 => std_logic_vector(to_unsigned(6,8) ,
36126	 => std_logic_vector(to_unsigned(5,8) ,
36127	 => std_logic_vector(to_unsigned(19,8) ,
36128	 => std_logic_vector(to_unsigned(18,8) ,
36129	 => std_logic_vector(to_unsigned(7,8) ,
36130	 => std_logic_vector(to_unsigned(6,8) ,
36131	 => std_logic_vector(to_unsigned(10,8) ,
36132	 => std_logic_vector(to_unsigned(7,8) ,
36133	 => std_logic_vector(to_unsigned(19,8) ,
36134	 => std_logic_vector(to_unsigned(57,8) ,
36135	 => std_logic_vector(to_unsigned(51,8) ,
36136	 => std_logic_vector(to_unsigned(22,8) ,
36137	 => std_logic_vector(to_unsigned(2,8) ,
36138	 => std_logic_vector(to_unsigned(1,8) ,
36139	 => std_logic_vector(to_unsigned(0,8) ,
36140	 => std_logic_vector(to_unsigned(8,8) ,
36141	 => std_logic_vector(to_unsigned(130,8) ,
36142	 => std_logic_vector(to_unsigned(152,8) ,
36143	 => std_logic_vector(to_unsigned(138,8) ,
36144	 => std_logic_vector(to_unsigned(139,8) ,
36145	 => std_logic_vector(to_unsigned(146,8) ,
36146	 => std_logic_vector(to_unsigned(154,8) ,
36147	 => std_logic_vector(to_unsigned(154,8) ,
36148	 => std_logic_vector(to_unsigned(156,8) ,
36149	 => std_logic_vector(to_unsigned(151,8) ,
36150	 => std_logic_vector(to_unsigned(141,8) ,
36151	 => std_logic_vector(to_unsigned(142,8) ,
36152	 => std_logic_vector(to_unsigned(141,8) ,
36153	 => std_logic_vector(to_unsigned(131,8) ,
36154	 => std_logic_vector(to_unsigned(144,8) ,
36155	 => std_logic_vector(to_unsigned(139,8) ,
36156	 => std_logic_vector(to_unsigned(121,8) ,
36157	 => std_logic_vector(to_unsigned(109,8) ,
36158	 => std_logic_vector(to_unsigned(111,8) ,
36159	 => std_logic_vector(to_unsigned(119,8) ,
36160	 => std_logic_vector(to_unsigned(116,8) ,
36161	 => std_logic_vector(to_unsigned(10,8) ,
36162	 => std_logic_vector(to_unsigned(11,8) ,
36163	 => std_logic_vector(to_unsigned(14,8) ,
36164	 => std_logic_vector(to_unsigned(14,8) ,
36165	 => std_logic_vector(to_unsigned(13,8) ,
36166	 => std_logic_vector(to_unsigned(17,8) ,
36167	 => std_logic_vector(to_unsigned(23,8) ,
36168	 => std_logic_vector(to_unsigned(35,8) ,
36169	 => std_logic_vector(to_unsigned(24,8) ,
36170	 => std_logic_vector(to_unsigned(3,8) ,
36171	 => std_logic_vector(to_unsigned(2,8) ,
36172	 => std_logic_vector(to_unsigned(1,8) ,
36173	 => std_logic_vector(to_unsigned(1,8) ,
36174	 => std_logic_vector(to_unsigned(1,8) ,
36175	 => std_logic_vector(to_unsigned(1,8) ,
36176	 => std_logic_vector(to_unsigned(0,8) ,
36177	 => std_logic_vector(to_unsigned(0,8) ,
36178	 => std_logic_vector(to_unsigned(0,8) ,
36179	 => std_logic_vector(to_unsigned(0,8) ,
36180	 => std_logic_vector(to_unsigned(0,8) ,
36181	 => std_logic_vector(to_unsigned(0,8) ,
36182	 => std_logic_vector(to_unsigned(0,8) ,
36183	 => std_logic_vector(to_unsigned(0,8) ,
36184	 => std_logic_vector(to_unsigned(0,8) ,
36185	 => std_logic_vector(to_unsigned(0,8) ,
36186	 => std_logic_vector(to_unsigned(0,8) ,
36187	 => std_logic_vector(to_unsigned(0,8) ,
36188	 => std_logic_vector(to_unsigned(0,8) ,
36189	 => std_logic_vector(to_unsigned(0,8) ,
36190	 => std_logic_vector(to_unsigned(0,8) ,
36191	 => std_logic_vector(to_unsigned(2,8) ,
36192	 => std_logic_vector(to_unsigned(17,8) ,
36193	 => std_logic_vector(to_unsigned(20,8) ,
36194	 => std_logic_vector(to_unsigned(23,8) ,
36195	 => std_logic_vector(to_unsigned(9,8) ,
36196	 => std_logic_vector(to_unsigned(3,8) ,
36197	 => std_logic_vector(to_unsigned(4,8) ,
36198	 => std_logic_vector(to_unsigned(3,8) ,
36199	 => std_logic_vector(to_unsigned(2,8) ,
36200	 => std_logic_vector(to_unsigned(3,8) ,
36201	 => std_logic_vector(to_unsigned(6,8) ,
36202	 => std_logic_vector(to_unsigned(7,8) ,
36203	 => std_logic_vector(to_unsigned(5,8) ,
36204	 => std_logic_vector(to_unsigned(7,8) ,
36205	 => std_logic_vector(to_unsigned(2,8) ,
36206	 => std_logic_vector(to_unsigned(0,8) ,
36207	 => std_logic_vector(to_unsigned(0,8) ,
36208	 => std_logic_vector(to_unsigned(0,8) ,
36209	 => std_logic_vector(to_unsigned(0,8) ,
36210	 => std_logic_vector(to_unsigned(1,8) ,
36211	 => std_logic_vector(to_unsigned(1,8) ,
36212	 => std_logic_vector(to_unsigned(3,8) ,
36213	 => std_logic_vector(to_unsigned(2,8) ,
36214	 => std_logic_vector(to_unsigned(2,8) ,
36215	 => std_logic_vector(to_unsigned(9,8) ,
36216	 => std_logic_vector(to_unsigned(11,8) ,
36217	 => std_logic_vector(to_unsigned(8,8) ,
36218	 => std_logic_vector(to_unsigned(8,8) ,
36219	 => std_logic_vector(to_unsigned(8,8) ,
36220	 => std_logic_vector(to_unsigned(9,8) ,
36221	 => std_logic_vector(to_unsigned(7,8) ,
36222	 => std_logic_vector(to_unsigned(6,8) ,
36223	 => std_logic_vector(to_unsigned(5,8) ,
36224	 => std_logic_vector(to_unsigned(3,8) ,
36225	 => std_logic_vector(to_unsigned(2,8) ,
36226	 => std_logic_vector(to_unsigned(2,8) ,
36227	 => std_logic_vector(to_unsigned(0,8) ,
36228	 => std_logic_vector(to_unsigned(0,8) ,
36229	 => std_logic_vector(to_unsigned(6,8) ,
36230	 => std_logic_vector(to_unsigned(15,8) ,
36231	 => std_logic_vector(to_unsigned(8,8) ,
36232	 => std_logic_vector(to_unsigned(5,8) ,
36233	 => std_logic_vector(to_unsigned(12,8) ,
36234	 => std_logic_vector(to_unsigned(6,8) ,
36235	 => std_logic_vector(to_unsigned(0,8) ,
36236	 => std_logic_vector(to_unsigned(1,8) ,
36237	 => std_logic_vector(to_unsigned(10,8) ,
36238	 => std_logic_vector(to_unsigned(8,8) ,
36239	 => std_logic_vector(to_unsigned(3,8) ,
36240	 => std_logic_vector(to_unsigned(6,8) ,
36241	 => std_logic_vector(to_unsigned(5,8) ,
36242	 => std_logic_vector(to_unsigned(5,8) ,
36243	 => std_logic_vector(to_unsigned(3,8) ,
36244	 => std_logic_vector(to_unsigned(4,8) ,
36245	 => std_logic_vector(to_unsigned(1,8) ,
36246	 => std_logic_vector(to_unsigned(2,8) ,
36247	 => std_logic_vector(to_unsigned(1,8) ,
36248	 => std_logic_vector(to_unsigned(0,8) ,
36249	 => std_logic_vector(to_unsigned(0,8) ,
36250	 => std_logic_vector(to_unsigned(0,8) ,
36251	 => std_logic_vector(to_unsigned(1,8) ,
36252	 => std_logic_vector(to_unsigned(8,8) ,
36253	 => std_logic_vector(to_unsigned(12,8) ,
36254	 => std_logic_vector(to_unsigned(9,8) ,
36255	 => std_logic_vector(to_unsigned(10,8) ,
36256	 => std_logic_vector(to_unsigned(10,8) ,
36257	 => std_logic_vector(to_unsigned(10,8) ,
36258	 => std_logic_vector(to_unsigned(5,8) ,
36259	 => std_logic_vector(to_unsigned(3,8) ,
36260	 => std_logic_vector(to_unsigned(9,8) ,
36261	 => std_logic_vector(to_unsigned(10,8) ,
36262	 => std_logic_vector(to_unsigned(7,8) ,
36263	 => std_logic_vector(to_unsigned(3,8) ,
36264	 => std_logic_vector(to_unsigned(3,8) ,
36265	 => std_logic_vector(to_unsigned(3,8) ,
36266	 => std_logic_vector(to_unsigned(4,8) ,
36267	 => std_logic_vector(to_unsigned(10,8) ,
36268	 => std_logic_vector(to_unsigned(8,8) ,
36269	 => std_logic_vector(to_unsigned(8,8) ,
36270	 => std_logic_vector(to_unsigned(5,8) ,
36271	 => std_logic_vector(to_unsigned(53,8) ,
36272	 => std_logic_vector(to_unsigned(183,8) ,
36273	 => std_logic_vector(to_unsigned(152,8) ,
36274	 => std_logic_vector(to_unsigned(27,8) ,
36275	 => std_logic_vector(to_unsigned(0,8) ,
36276	 => std_logic_vector(to_unsigned(0,8) ,
36277	 => std_logic_vector(to_unsigned(1,8) ,
36278	 => std_logic_vector(to_unsigned(1,8) ,
36279	 => std_logic_vector(to_unsigned(0,8) ,
36280	 => std_logic_vector(to_unsigned(0,8) ,
36281	 => std_logic_vector(to_unsigned(1,8) ,
36282	 => std_logic_vector(to_unsigned(6,8) ,
36283	 => std_logic_vector(to_unsigned(6,8) ,
36284	 => std_logic_vector(to_unsigned(7,8) ,
36285	 => std_logic_vector(to_unsigned(12,8) ,
36286	 => std_logic_vector(to_unsigned(4,8) ,
36287	 => std_logic_vector(to_unsigned(2,8) ,
36288	 => std_logic_vector(to_unsigned(4,8) ,
36289	 => std_logic_vector(to_unsigned(1,8) ,
36290	 => std_logic_vector(to_unsigned(0,8) ,
36291	 => std_logic_vector(to_unsigned(3,8) ,
36292	 => std_logic_vector(to_unsigned(6,8) ,
36293	 => std_logic_vector(to_unsigned(3,8) ,
36294	 => std_logic_vector(to_unsigned(3,8) ,
36295	 => std_logic_vector(to_unsigned(4,8) ,
36296	 => std_logic_vector(to_unsigned(3,8) ,
36297	 => std_logic_vector(to_unsigned(2,8) ,
36298	 => std_logic_vector(to_unsigned(2,8) ,
36299	 => std_logic_vector(to_unsigned(1,8) ,
36300	 => std_logic_vector(to_unsigned(1,8) ,
36301	 => std_logic_vector(to_unsigned(0,8) ,
36302	 => std_logic_vector(to_unsigned(0,8) ,
36303	 => std_logic_vector(to_unsigned(0,8) ,
36304	 => std_logic_vector(to_unsigned(0,8) ,
36305	 => std_logic_vector(to_unsigned(1,8) ,
36306	 => std_logic_vector(to_unsigned(1,8) ,
36307	 => std_logic_vector(to_unsigned(2,8) ,
36308	 => std_logic_vector(to_unsigned(2,8) ,
36309	 => std_logic_vector(to_unsigned(2,8) ,
36310	 => std_logic_vector(to_unsigned(2,8) ,
36311	 => std_logic_vector(to_unsigned(2,8) ,
36312	 => std_logic_vector(to_unsigned(2,8) ,
36313	 => std_logic_vector(to_unsigned(5,8) ,
36314	 => std_logic_vector(to_unsigned(7,8) ,
36315	 => std_logic_vector(to_unsigned(10,8) ,
36316	 => std_logic_vector(to_unsigned(5,8) ,
36317	 => std_logic_vector(to_unsigned(1,8) ,
36318	 => std_logic_vector(to_unsigned(1,8) ,
36319	 => std_logic_vector(to_unsigned(3,8) ,
36320	 => std_logic_vector(to_unsigned(12,8) ,
36321	 => std_logic_vector(to_unsigned(9,8) ,
36322	 => std_logic_vector(to_unsigned(4,8) ,
36323	 => std_logic_vector(to_unsigned(4,8) ,
36324	 => std_logic_vector(to_unsigned(5,8) ,
36325	 => std_logic_vector(to_unsigned(5,8) ,
36326	 => std_logic_vector(to_unsigned(3,8) ,
36327	 => std_logic_vector(to_unsigned(0,8) ,
36328	 => std_logic_vector(to_unsigned(0,8) ,
36329	 => std_logic_vector(to_unsigned(0,8) ,
36330	 => std_logic_vector(to_unsigned(0,8) ,
36331	 => std_logic_vector(to_unsigned(1,8) ,
36332	 => std_logic_vector(to_unsigned(1,8) ,
36333	 => std_logic_vector(to_unsigned(0,8) ,
36334	 => std_logic_vector(to_unsigned(2,8) ,
36335	 => std_logic_vector(to_unsigned(2,8) ,
36336	 => std_logic_vector(to_unsigned(2,8) ,
36337	 => std_logic_vector(to_unsigned(4,8) ,
36338	 => std_logic_vector(to_unsigned(6,8) ,
36339	 => std_logic_vector(to_unsigned(6,8) ,
36340	 => std_logic_vector(to_unsigned(3,8) ,
36341	 => std_logic_vector(to_unsigned(1,8) ,
36342	 => std_logic_vector(to_unsigned(2,8) ,
36343	 => std_logic_vector(to_unsigned(4,8) ,
36344	 => std_logic_vector(to_unsigned(3,8) ,
36345	 => std_logic_vector(to_unsigned(3,8) ,
36346	 => std_logic_vector(to_unsigned(2,8) ,
36347	 => std_logic_vector(to_unsigned(2,8) ,
36348	 => std_logic_vector(to_unsigned(2,8) ,
36349	 => std_logic_vector(to_unsigned(1,8) ,
36350	 => std_logic_vector(to_unsigned(0,8) ,
36351	 => std_logic_vector(to_unsigned(0,8) ,
36352	 => std_logic_vector(to_unsigned(0,8) ,
36353	 => std_logic_vector(to_unsigned(0,8) ,
36354	 => std_logic_vector(to_unsigned(1,8) ,
36355	 => std_logic_vector(to_unsigned(2,8) ,
36356	 => std_logic_vector(to_unsigned(2,8) ,
36357	 => std_logic_vector(to_unsigned(3,8) ,
36358	 => std_logic_vector(to_unsigned(3,8) ,
36359	 => std_logic_vector(to_unsigned(3,8) ,
36360	 => std_logic_vector(to_unsigned(4,8) ,
36361	 => std_logic_vector(to_unsigned(4,8) ,
36362	 => std_logic_vector(to_unsigned(3,8) ,
36363	 => std_logic_vector(to_unsigned(4,8) ,
36364	 => std_logic_vector(to_unsigned(4,8) ,
36365	 => std_logic_vector(to_unsigned(2,8) ,
36366	 => std_logic_vector(to_unsigned(1,8) ,
36367	 => std_logic_vector(to_unsigned(2,8) ,
36368	 => std_logic_vector(to_unsigned(1,8) ,
36369	 => std_logic_vector(to_unsigned(2,8) ,
36370	 => std_logic_vector(to_unsigned(3,8) ,
36371	 => std_logic_vector(to_unsigned(3,8) ,
36372	 => std_logic_vector(to_unsigned(1,8) ,
36373	 => std_logic_vector(to_unsigned(6,8) ,
36374	 => std_logic_vector(to_unsigned(15,8) ,
36375	 => std_logic_vector(to_unsigned(11,8) ,
36376	 => std_logic_vector(to_unsigned(9,8) ,
36377	 => std_logic_vector(to_unsigned(10,8) ,
36378	 => std_logic_vector(to_unsigned(13,8) ,
36379	 => std_logic_vector(to_unsigned(7,8) ,
36380	 => std_logic_vector(to_unsigned(3,8) ,
36381	 => std_logic_vector(to_unsigned(2,8) ,
36382	 => std_logic_vector(to_unsigned(4,8) ,
36383	 => std_logic_vector(to_unsigned(25,8) ,
36384	 => std_logic_vector(to_unsigned(81,8) ,
36385	 => std_logic_vector(to_unsigned(25,8) ,
36386	 => std_logic_vector(to_unsigned(0,8) ,
36387	 => std_logic_vector(to_unsigned(1,8) ,
36388	 => std_logic_vector(to_unsigned(5,8) ,
36389	 => std_logic_vector(to_unsigned(11,8) ,
36390	 => std_logic_vector(to_unsigned(37,8) ,
36391	 => std_logic_vector(to_unsigned(50,8) ,
36392	 => std_logic_vector(to_unsigned(46,8) ,
36393	 => std_logic_vector(to_unsigned(36,8) ,
36394	 => std_logic_vector(to_unsigned(21,8) ,
36395	 => std_logic_vector(to_unsigned(10,8) ,
36396	 => std_logic_vector(to_unsigned(3,8) ,
36397	 => std_logic_vector(to_unsigned(3,8) ,
36398	 => std_logic_vector(to_unsigned(4,8) ,
36399	 => std_logic_vector(to_unsigned(1,8) ,
36400	 => std_logic_vector(to_unsigned(1,8) ,
36401	 => std_logic_vector(to_unsigned(1,8) ,
36402	 => std_logic_vector(to_unsigned(1,8) ,
36403	 => std_logic_vector(to_unsigned(4,8) ,
36404	 => std_logic_vector(to_unsigned(24,8) ,
36405	 => std_logic_vector(to_unsigned(28,8) ,
36406	 => std_logic_vector(to_unsigned(22,8) ,
36407	 => std_logic_vector(to_unsigned(22,8) ,
36408	 => std_logic_vector(to_unsigned(30,8) ,
36409	 => std_logic_vector(to_unsigned(36,8) ,
36410	 => std_logic_vector(to_unsigned(44,8) ,
36411	 => std_logic_vector(to_unsigned(50,8) ,
36412	 => std_logic_vector(to_unsigned(57,8) ,
36413	 => std_logic_vector(to_unsigned(40,8) ,
36414	 => std_logic_vector(to_unsigned(9,8) ,
36415	 => std_logic_vector(to_unsigned(8,8) ,
36416	 => std_logic_vector(to_unsigned(6,8) ,
36417	 => std_logic_vector(to_unsigned(5,8) ,
36418	 => std_logic_vector(to_unsigned(3,8) ,
36419	 => std_logic_vector(to_unsigned(4,8) ,
36420	 => std_logic_vector(to_unsigned(6,8) ,
36421	 => std_logic_vector(to_unsigned(5,8) ,
36422	 => std_logic_vector(to_unsigned(6,8) ,
36423	 => std_logic_vector(to_unsigned(15,8) ,
36424	 => std_logic_vector(to_unsigned(32,8) ,
36425	 => std_logic_vector(to_unsigned(13,8) ,
36426	 => std_logic_vector(to_unsigned(7,8) ,
36427	 => std_logic_vector(to_unsigned(21,8) ,
36428	 => std_logic_vector(to_unsigned(53,8) ,
36429	 => std_logic_vector(to_unsigned(63,8) ,
36430	 => std_logic_vector(to_unsigned(28,8) ,
36431	 => std_logic_vector(to_unsigned(48,8) ,
36432	 => std_logic_vector(to_unsigned(32,8) ,
36433	 => std_logic_vector(to_unsigned(37,8) ,
36434	 => std_logic_vector(to_unsigned(8,8) ,
36435	 => std_logic_vector(to_unsigned(73,8) ,
36436	 => std_logic_vector(to_unsigned(22,8) ,
36437	 => std_logic_vector(to_unsigned(14,8) ,
36438	 => std_logic_vector(to_unsigned(7,8) ,
36439	 => std_logic_vector(to_unsigned(6,8) ,
36440	 => std_logic_vector(to_unsigned(4,8) ,
36441	 => std_logic_vector(to_unsigned(2,8) ,
36442	 => std_logic_vector(to_unsigned(1,8) ,
36443	 => std_logic_vector(to_unsigned(1,8) ,
36444	 => std_logic_vector(to_unsigned(1,8) ,
36445	 => std_logic_vector(to_unsigned(3,8) ,
36446	 => std_logic_vector(to_unsigned(8,8) ,
36447	 => std_logic_vector(to_unsigned(14,8) ,
36448	 => std_logic_vector(to_unsigned(12,8) ,
36449	 => std_logic_vector(to_unsigned(9,8) ,
36450	 => std_logic_vector(to_unsigned(9,8) ,
36451	 => std_logic_vector(to_unsigned(6,8) ,
36452	 => std_logic_vector(to_unsigned(18,8) ,
36453	 => std_logic_vector(to_unsigned(49,8) ,
36454	 => std_logic_vector(to_unsigned(19,8) ,
36455	 => std_logic_vector(to_unsigned(35,8) ,
36456	 => std_logic_vector(to_unsigned(19,8) ,
36457	 => std_logic_vector(to_unsigned(4,8) ,
36458	 => std_logic_vector(to_unsigned(3,8) ,
36459	 => std_logic_vector(to_unsigned(0,8) ,
36460	 => std_logic_vector(to_unsigned(22,8) ,
36461	 => std_logic_vector(to_unsigned(164,8) ,
36462	 => std_logic_vector(to_unsigned(156,8) ,
36463	 => std_logic_vector(to_unsigned(144,8) ,
36464	 => std_logic_vector(to_unsigned(141,8) ,
36465	 => std_logic_vector(to_unsigned(134,8) ,
36466	 => std_logic_vector(to_unsigned(142,8) ,
36467	 => std_logic_vector(to_unsigned(147,8) ,
36468	 => std_logic_vector(to_unsigned(159,8) ,
36469	 => std_logic_vector(to_unsigned(168,8) ,
36470	 => std_logic_vector(to_unsigned(152,8) ,
36471	 => std_logic_vector(to_unsigned(139,8) ,
36472	 => std_logic_vector(to_unsigned(144,8) ,
36473	 => std_logic_vector(to_unsigned(151,8) ,
36474	 => std_logic_vector(to_unsigned(163,8) ,
36475	 => std_logic_vector(to_unsigned(144,8) ,
36476	 => std_logic_vector(to_unsigned(119,8) ,
36477	 => std_logic_vector(to_unsigned(115,8) ,
36478	 => std_logic_vector(to_unsigned(115,8) ,
36479	 => std_logic_vector(to_unsigned(107,8) ,
36480	 => std_logic_vector(to_unsigned(107,8) ,
36481	 => std_logic_vector(to_unsigned(27,8) ,
36482	 => std_logic_vector(to_unsigned(21,8) ,
36483	 => std_logic_vector(to_unsigned(17,8) ,
36484	 => std_logic_vector(to_unsigned(10,8) ,
36485	 => std_logic_vector(to_unsigned(6,8) ,
36486	 => std_logic_vector(to_unsigned(12,8) ,
36487	 => std_logic_vector(to_unsigned(35,8) ,
36488	 => std_logic_vector(to_unsigned(27,8) ,
36489	 => std_logic_vector(to_unsigned(7,8) ,
36490	 => std_logic_vector(to_unsigned(2,8) ,
36491	 => std_logic_vector(to_unsigned(2,8) ,
36492	 => std_logic_vector(to_unsigned(2,8) ,
36493	 => std_logic_vector(to_unsigned(3,8) ,
36494	 => std_logic_vector(to_unsigned(1,8) ,
36495	 => std_logic_vector(to_unsigned(1,8) ,
36496	 => std_logic_vector(to_unsigned(1,8) ,
36497	 => std_logic_vector(to_unsigned(1,8) ,
36498	 => std_logic_vector(to_unsigned(1,8) ,
36499	 => std_logic_vector(to_unsigned(0,8) ,
36500	 => std_logic_vector(to_unsigned(0,8) ,
36501	 => std_logic_vector(to_unsigned(1,8) ,
36502	 => std_logic_vector(to_unsigned(0,8) ,
36503	 => std_logic_vector(to_unsigned(0,8) ,
36504	 => std_logic_vector(to_unsigned(0,8) ,
36505	 => std_logic_vector(to_unsigned(0,8) ,
36506	 => std_logic_vector(to_unsigned(0,8) ,
36507	 => std_logic_vector(to_unsigned(1,8) ,
36508	 => std_logic_vector(to_unsigned(1,8) ,
36509	 => std_logic_vector(to_unsigned(1,8) ,
36510	 => std_logic_vector(to_unsigned(1,8) ,
36511	 => std_logic_vector(to_unsigned(3,8) ,
36512	 => std_logic_vector(to_unsigned(15,8) ,
36513	 => std_logic_vector(to_unsigned(14,8) ,
36514	 => std_logic_vector(to_unsigned(12,8) ,
36515	 => std_logic_vector(to_unsigned(4,8) ,
36516	 => std_logic_vector(to_unsigned(4,8) ,
36517	 => std_logic_vector(to_unsigned(5,8) ,
36518	 => std_logic_vector(to_unsigned(3,8) ,
36519	 => std_logic_vector(to_unsigned(3,8) ,
36520	 => std_logic_vector(to_unsigned(3,8) ,
36521	 => std_logic_vector(to_unsigned(4,8) ,
36522	 => std_logic_vector(to_unsigned(4,8) ,
36523	 => std_logic_vector(to_unsigned(3,8) ,
36524	 => std_logic_vector(to_unsigned(4,8) ,
36525	 => std_logic_vector(to_unsigned(1,8) ,
36526	 => std_logic_vector(to_unsigned(0,8) ,
36527	 => std_logic_vector(to_unsigned(1,8) ,
36528	 => std_logic_vector(to_unsigned(1,8) ,
36529	 => std_logic_vector(to_unsigned(1,8) ,
36530	 => std_logic_vector(to_unsigned(1,8) ,
36531	 => std_logic_vector(to_unsigned(1,8) ,
36532	 => std_logic_vector(to_unsigned(1,8) ,
36533	 => std_logic_vector(to_unsigned(2,8) ,
36534	 => std_logic_vector(to_unsigned(1,8) ,
36535	 => std_logic_vector(to_unsigned(5,8) ,
36536	 => std_logic_vector(to_unsigned(11,8) ,
36537	 => std_logic_vector(to_unsigned(8,8) ,
36538	 => std_logic_vector(to_unsigned(8,8) ,
36539	 => std_logic_vector(to_unsigned(7,8) ,
36540	 => std_logic_vector(to_unsigned(7,8) ,
36541	 => std_logic_vector(to_unsigned(7,8) ,
36542	 => std_logic_vector(to_unsigned(4,8) ,
36543	 => std_logic_vector(to_unsigned(3,8) ,
36544	 => std_logic_vector(to_unsigned(3,8) ,
36545	 => std_logic_vector(to_unsigned(2,8) ,
36546	 => std_logic_vector(to_unsigned(1,8) ,
36547	 => std_logic_vector(to_unsigned(0,8) ,
36548	 => std_logic_vector(to_unsigned(1,8) ,
36549	 => std_logic_vector(to_unsigned(4,8) ,
36550	 => std_logic_vector(to_unsigned(17,8) ,
36551	 => std_logic_vector(to_unsigned(20,8) ,
36552	 => std_logic_vector(to_unsigned(12,8) ,
36553	 => std_logic_vector(to_unsigned(8,8) ,
36554	 => std_logic_vector(to_unsigned(2,8) ,
36555	 => std_logic_vector(to_unsigned(0,8) ,
36556	 => std_logic_vector(to_unsigned(1,8) ,
36557	 => std_logic_vector(to_unsigned(9,8) ,
36558	 => std_logic_vector(to_unsigned(9,8) ,
36559	 => std_logic_vector(to_unsigned(4,8) ,
36560	 => std_logic_vector(to_unsigned(6,8) ,
36561	 => std_logic_vector(to_unsigned(7,8) ,
36562	 => std_logic_vector(to_unsigned(6,8) ,
36563	 => std_logic_vector(to_unsigned(6,8) ,
36564	 => std_logic_vector(to_unsigned(4,8) ,
36565	 => std_logic_vector(to_unsigned(1,8) ,
36566	 => std_logic_vector(to_unsigned(4,8) ,
36567	 => std_logic_vector(to_unsigned(1,8) ,
36568	 => std_logic_vector(to_unsigned(0,8) ,
36569	 => std_logic_vector(to_unsigned(0,8) ,
36570	 => std_logic_vector(to_unsigned(0,8) ,
36571	 => std_logic_vector(to_unsigned(0,8) ,
36572	 => std_logic_vector(to_unsigned(5,8) ,
36573	 => std_logic_vector(to_unsigned(13,8) ,
36574	 => std_logic_vector(to_unsigned(10,8) ,
36575	 => std_logic_vector(to_unsigned(10,8) ,
36576	 => std_logic_vector(to_unsigned(9,8) ,
36577	 => std_logic_vector(to_unsigned(7,8) ,
36578	 => std_logic_vector(to_unsigned(6,8) ,
36579	 => std_logic_vector(to_unsigned(3,8) ,
36580	 => std_logic_vector(to_unsigned(8,8) ,
36581	 => std_logic_vector(to_unsigned(14,8) ,
36582	 => std_logic_vector(to_unsigned(8,8) ,
36583	 => std_logic_vector(to_unsigned(5,8) ,
36584	 => std_logic_vector(to_unsigned(4,8) ,
36585	 => std_logic_vector(to_unsigned(3,8) ,
36586	 => std_logic_vector(to_unsigned(3,8) ,
36587	 => std_logic_vector(to_unsigned(2,8) ,
36588	 => std_logic_vector(to_unsigned(4,8) ,
36589	 => std_logic_vector(to_unsigned(6,8) ,
36590	 => std_logic_vector(to_unsigned(6,8) ,
36591	 => std_logic_vector(to_unsigned(84,8) ,
36592	 => std_logic_vector(to_unsigned(161,8) ,
36593	 => std_logic_vector(to_unsigned(166,8) ,
36594	 => std_logic_vector(to_unsigned(116,8) ,
36595	 => std_logic_vector(to_unsigned(5,8) ,
36596	 => std_logic_vector(to_unsigned(0,8) ,
36597	 => std_logic_vector(to_unsigned(1,8) ,
36598	 => std_logic_vector(to_unsigned(1,8) ,
36599	 => std_logic_vector(to_unsigned(1,8) ,
36600	 => std_logic_vector(to_unsigned(0,8) ,
36601	 => std_logic_vector(to_unsigned(0,8) ,
36602	 => std_logic_vector(to_unsigned(4,8) ,
36603	 => std_logic_vector(to_unsigned(5,8) ,
36604	 => std_logic_vector(to_unsigned(7,8) ,
36605	 => std_logic_vector(to_unsigned(10,8) ,
36606	 => std_logic_vector(to_unsigned(3,8) ,
36607	 => std_logic_vector(to_unsigned(5,8) ,
36608	 => std_logic_vector(to_unsigned(4,8) ,
36609	 => std_logic_vector(to_unsigned(2,8) ,
36610	 => std_logic_vector(to_unsigned(0,8) ,
36611	 => std_logic_vector(to_unsigned(3,8) ,
36612	 => std_logic_vector(to_unsigned(6,8) ,
36613	 => std_logic_vector(to_unsigned(3,8) ,
36614	 => std_logic_vector(to_unsigned(3,8) ,
36615	 => std_logic_vector(to_unsigned(5,8) ,
36616	 => std_logic_vector(to_unsigned(3,8) ,
36617	 => std_logic_vector(to_unsigned(2,8) ,
36618	 => std_logic_vector(to_unsigned(2,8) ,
36619	 => std_logic_vector(to_unsigned(3,8) ,
36620	 => std_logic_vector(to_unsigned(2,8) ,
36621	 => std_logic_vector(to_unsigned(0,8) ,
36622	 => std_logic_vector(to_unsigned(0,8) ,
36623	 => std_logic_vector(to_unsigned(1,8) ,
36624	 => std_logic_vector(to_unsigned(0,8) ,
36625	 => std_logic_vector(to_unsigned(1,8) ,
36626	 => std_logic_vector(to_unsigned(2,8) ,
36627	 => std_logic_vector(to_unsigned(2,8) ,
36628	 => std_logic_vector(to_unsigned(2,8) ,
36629	 => std_logic_vector(to_unsigned(3,8) ,
36630	 => std_logic_vector(to_unsigned(3,8) ,
36631	 => std_logic_vector(to_unsigned(2,8) ,
36632	 => std_logic_vector(to_unsigned(4,8) ,
36633	 => std_logic_vector(to_unsigned(5,8) ,
36634	 => std_logic_vector(to_unsigned(7,8) ,
36635	 => std_logic_vector(to_unsigned(11,8) ,
36636	 => std_logic_vector(to_unsigned(5,8) ,
36637	 => std_logic_vector(to_unsigned(2,8) ,
36638	 => std_logic_vector(to_unsigned(1,8) ,
36639	 => std_logic_vector(to_unsigned(4,8) ,
36640	 => std_logic_vector(to_unsigned(13,8) ,
36641	 => std_logic_vector(to_unsigned(6,8) ,
36642	 => std_logic_vector(to_unsigned(4,8) ,
36643	 => std_logic_vector(to_unsigned(4,8) ,
36644	 => std_logic_vector(to_unsigned(5,8) ,
36645	 => std_logic_vector(to_unsigned(6,8) ,
36646	 => std_logic_vector(to_unsigned(3,8) ,
36647	 => std_logic_vector(to_unsigned(0,8) ,
36648	 => std_logic_vector(to_unsigned(0,8) ,
36649	 => std_logic_vector(to_unsigned(0,8) ,
36650	 => std_logic_vector(to_unsigned(1,8) ,
36651	 => std_logic_vector(to_unsigned(0,8) ,
36652	 => std_logic_vector(to_unsigned(1,8) ,
36653	 => std_logic_vector(to_unsigned(1,8) ,
36654	 => std_logic_vector(to_unsigned(2,8) ,
36655	 => std_logic_vector(to_unsigned(2,8) ,
36656	 => std_logic_vector(to_unsigned(2,8) ,
36657	 => std_logic_vector(to_unsigned(5,8) ,
36658	 => std_logic_vector(to_unsigned(6,8) ,
36659	 => std_logic_vector(to_unsigned(7,8) ,
36660	 => std_logic_vector(to_unsigned(3,8) ,
36661	 => std_logic_vector(to_unsigned(0,8) ,
36662	 => std_logic_vector(to_unsigned(2,8) ,
36663	 => std_logic_vector(to_unsigned(6,8) ,
36664	 => std_logic_vector(to_unsigned(2,8) ,
36665	 => std_logic_vector(to_unsigned(3,8) ,
36666	 => std_logic_vector(to_unsigned(3,8) ,
36667	 => std_logic_vector(to_unsigned(2,8) ,
36668	 => std_logic_vector(to_unsigned(2,8) ,
36669	 => std_logic_vector(to_unsigned(2,8) ,
36670	 => std_logic_vector(to_unsigned(1,8) ,
36671	 => std_logic_vector(to_unsigned(1,8) ,
36672	 => std_logic_vector(to_unsigned(0,8) ,
36673	 => std_logic_vector(to_unsigned(0,8) ,
36674	 => std_logic_vector(to_unsigned(0,8) ,
36675	 => std_logic_vector(to_unsigned(0,8) ,
36676	 => std_logic_vector(to_unsigned(0,8) ,
36677	 => std_logic_vector(to_unsigned(0,8) ,
36678	 => std_logic_vector(to_unsigned(0,8) ,
36679	 => std_logic_vector(to_unsigned(0,8) ,
36680	 => std_logic_vector(to_unsigned(1,8) ,
36681	 => std_logic_vector(to_unsigned(1,8) ,
36682	 => std_logic_vector(to_unsigned(1,8) ,
36683	 => std_logic_vector(to_unsigned(1,8) ,
36684	 => std_logic_vector(to_unsigned(2,8) ,
36685	 => std_logic_vector(to_unsigned(2,8) ,
36686	 => std_logic_vector(to_unsigned(2,8) ,
36687	 => std_logic_vector(to_unsigned(1,8) ,
36688	 => std_logic_vector(to_unsigned(1,8) ,
36689	 => std_logic_vector(to_unsigned(3,8) ,
36690	 => std_logic_vector(to_unsigned(4,8) ,
36691	 => std_logic_vector(to_unsigned(4,8) ,
36692	 => std_logic_vector(to_unsigned(1,8) ,
36693	 => std_logic_vector(to_unsigned(9,8) ,
36694	 => std_logic_vector(to_unsigned(18,8) ,
36695	 => std_logic_vector(to_unsigned(12,8) ,
36696	 => std_logic_vector(to_unsigned(8,8) ,
36697	 => std_logic_vector(to_unsigned(14,8) ,
36698	 => std_logic_vector(to_unsigned(15,8) ,
36699	 => std_logic_vector(to_unsigned(9,8) ,
36700	 => std_logic_vector(to_unsigned(6,8) ,
36701	 => std_logic_vector(to_unsigned(6,8) ,
36702	 => std_logic_vector(to_unsigned(0,8) ,
36703	 => std_logic_vector(to_unsigned(0,8) ,
36704	 => std_logic_vector(to_unsigned(2,8) ,
36705	 => std_logic_vector(to_unsigned(1,8) ,
36706	 => std_logic_vector(to_unsigned(0,8) ,
36707	 => std_logic_vector(to_unsigned(2,8) ,
36708	 => std_logic_vector(to_unsigned(9,8) ,
36709	 => std_logic_vector(to_unsigned(16,8) ,
36710	 => std_logic_vector(to_unsigned(41,8) ,
36711	 => std_logic_vector(to_unsigned(59,8) ,
36712	 => std_logic_vector(to_unsigned(50,8) ,
36713	 => std_logic_vector(to_unsigned(40,8) ,
36714	 => std_logic_vector(to_unsigned(25,8) ,
36715	 => std_logic_vector(to_unsigned(9,8) ,
36716	 => std_logic_vector(to_unsigned(2,8) ,
36717	 => std_logic_vector(to_unsigned(3,8) ,
36718	 => std_logic_vector(to_unsigned(5,8) ,
36719	 => std_logic_vector(to_unsigned(4,8) ,
36720	 => std_logic_vector(to_unsigned(3,8) ,
36721	 => std_logic_vector(to_unsigned(1,8) ,
36722	 => std_logic_vector(to_unsigned(1,8) ,
36723	 => std_logic_vector(to_unsigned(1,8) ,
36724	 => std_logic_vector(to_unsigned(23,8) ,
36725	 => std_logic_vector(to_unsigned(35,8) ,
36726	 => std_logic_vector(to_unsigned(10,8) ,
36727	 => std_logic_vector(to_unsigned(1,8) ,
36728	 => std_logic_vector(to_unsigned(2,8) ,
36729	 => std_logic_vector(to_unsigned(2,8) ,
36730	 => std_logic_vector(to_unsigned(1,8) ,
36731	 => std_logic_vector(to_unsigned(1,8) ,
36732	 => std_logic_vector(to_unsigned(1,8) ,
36733	 => std_logic_vector(to_unsigned(1,8) ,
36734	 => std_logic_vector(to_unsigned(1,8) ,
36735	 => std_logic_vector(to_unsigned(1,8) ,
36736	 => std_logic_vector(to_unsigned(2,8) ,
36737	 => std_logic_vector(to_unsigned(2,8) ,
36738	 => std_logic_vector(to_unsigned(2,8) ,
36739	 => std_logic_vector(to_unsigned(2,8) ,
36740	 => std_logic_vector(to_unsigned(3,8) ,
36741	 => std_logic_vector(to_unsigned(3,8) ,
36742	 => std_logic_vector(to_unsigned(9,8) ,
36743	 => std_logic_vector(to_unsigned(29,8) ,
36744	 => std_logic_vector(to_unsigned(30,8) ,
36745	 => std_logic_vector(to_unsigned(23,8) ,
36746	 => std_logic_vector(to_unsigned(9,8) ,
36747	 => std_logic_vector(to_unsigned(14,8) ,
36748	 => std_logic_vector(to_unsigned(37,8) ,
36749	 => std_logic_vector(to_unsigned(82,8) ,
36750	 => std_logic_vector(to_unsigned(35,8) ,
36751	 => std_logic_vector(to_unsigned(43,8) ,
36752	 => std_logic_vector(to_unsigned(31,8) ,
36753	 => std_logic_vector(to_unsigned(45,8) ,
36754	 => std_logic_vector(to_unsigned(4,8) ,
36755	 => std_logic_vector(to_unsigned(21,8) ,
36756	 => std_logic_vector(to_unsigned(24,8) ,
36757	 => std_logic_vector(to_unsigned(15,8) ,
36758	 => std_logic_vector(to_unsigned(13,8) ,
36759	 => std_logic_vector(to_unsigned(2,8) ,
36760	 => std_logic_vector(to_unsigned(10,8) ,
36761	 => std_logic_vector(to_unsigned(8,8) ,
36762	 => std_logic_vector(to_unsigned(4,8) ,
36763	 => std_logic_vector(to_unsigned(3,8) ,
36764	 => std_logic_vector(to_unsigned(4,8) ,
36765	 => std_logic_vector(to_unsigned(6,8) ,
36766	 => std_logic_vector(to_unsigned(9,8) ,
36767	 => std_logic_vector(to_unsigned(16,8) ,
36768	 => std_logic_vector(to_unsigned(21,8) ,
36769	 => std_logic_vector(to_unsigned(13,8) ,
36770	 => std_logic_vector(to_unsigned(8,8) ,
36771	 => std_logic_vector(to_unsigned(14,8) ,
36772	 => std_logic_vector(to_unsigned(24,8) ,
36773	 => std_logic_vector(to_unsigned(9,8) ,
36774	 => std_logic_vector(to_unsigned(6,8) ,
36775	 => std_logic_vector(to_unsigned(62,8) ,
36776	 => std_logic_vector(to_unsigned(20,8) ,
36777	 => std_logic_vector(to_unsigned(4,8) ,
36778	 => std_logic_vector(to_unsigned(4,8) ,
36779	 => std_logic_vector(to_unsigned(0,8) ,
36780	 => std_logic_vector(to_unsigned(51,8) ,
36781	 => std_logic_vector(to_unsigned(168,8) ,
36782	 => std_logic_vector(to_unsigned(149,8) ,
36783	 => std_logic_vector(to_unsigned(147,8) ,
36784	 => std_logic_vector(to_unsigned(134,8) ,
36785	 => std_logic_vector(to_unsigned(136,8) ,
36786	 => std_logic_vector(to_unsigned(154,8) ,
36787	 => std_logic_vector(to_unsigned(163,8) ,
36788	 => std_logic_vector(to_unsigned(166,8) ,
36789	 => std_logic_vector(to_unsigned(164,8) ,
36790	 => std_logic_vector(to_unsigned(161,8) ,
36791	 => std_logic_vector(to_unsigned(152,8) ,
36792	 => std_logic_vector(to_unsigned(147,8) ,
36793	 => std_logic_vector(to_unsigned(151,8) ,
36794	 => std_logic_vector(to_unsigned(163,8) ,
36795	 => std_logic_vector(to_unsigned(152,8) ,
36796	 => std_logic_vector(to_unsigned(133,8) ,
36797	 => std_logic_vector(to_unsigned(131,8) ,
36798	 => std_logic_vector(to_unsigned(131,8) ,
36799	 => std_logic_vector(to_unsigned(122,8) ,
36800	 => std_logic_vector(to_unsigned(131,8) ,
36801	 => std_logic_vector(to_unsigned(147,8) ,
36802	 => std_logic_vector(to_unsigned(138,8) ,
36803	 => std_logic_vector(to_unsigned(130,8) ,
36804	 => std_logic_vector(to_unsigned(111,8) ,
36805	 => std_logic_vector(to_unsigned(95,8) ,
36806	 => std_logic_vector(to_unsigned(53,8) ,
36807	 => std_logic_vector(to_unsigned(11,8) ,
36808	 => std_logic_vector(to_unsigned(6,8) ,
36809	 => std_logic_vector(to_unsigned(4,8) ,
36810	 => std_logic_vector(to_unsigned(1,8) ,
36811	 => std_logic_vector(to_unsigned(1,8) ,
36812	 => std_logic_vector(to_unsigned(2,8) ,
36813	 => std_logic_vector(to_unsigned(2,8) ,
36814	 => std_logic_vector(to_unsigned(1,8) ,
36815	 => std_logic_vector(to_unsigned(0,8) ,
36816	 => std_logic_vector(to_unsigned(0,8) ,
36817	 => std_logic_vector(to_unsigned(1,8) ,
36818	 => std_logic_vector(to_unsigned(1,8) ,
36819	 => std_logic_vector(to_unsigned(0,8) ,
36820	 => std_logic_vector(to_unsigned(0,8) ,
36821	 => std_logic_vector(to_unsigned(0,8) ,
36822	 => std_logic_vector(to_unsigned(0,8) ,
36823	 => std_logic_vector(to_unsigned(0,8) ,
36824	 => std_logic_vector(to_unsigned(0,8) ,
36825	 => std_logic_vector(to_unsigned(0,8) ,
36826	 => std_logic_vector(to_unsigned(0,8) ,
36827	 => std_logic_vector(to_unsigned(1,8) ,
36828	 => std_logic_vector(to_unsigned(1,8) ,
36829	 => std_logic_vector(to_unsigned(1,8) ,
36830	 => std_logic_vector(to_unsigned(1,8) ,
36831	 => std_logic_vector(to_unsigned(6,8) ,
36832	 => std_logic_vector(to_unsigned(20,8) ,
36833	 => std_logic_vector(to_unsigned(10,8) ,
36834	 => std_logic_vector(to_unsigned(9,8) ,
36835	 => std_logic_vector(to_unsigned(7,8) ,
36836	 => std_logic_vector(to_unsigned(7,8) ,
36837	 => std_logic_vector(to_unsigned(8,8) ,
36838	 => std_logic_vector(to_unsigned(4,8) ,
36839	 => std_logic_vector(to_unsigned(4,8) ,
36840	 => std_logic_vector(to_unsigned(2,8) ,
36841	 => std_logic_vector(to_unsigned(3,8) ,
36842	 => std_logic_vector(to_unsigned(3,8) ,
36843	 => std_logic_vector(to_unsigned(2,8) ,
36844	 => std_logic_vector(to_unsigned(3,8) ,
36845	 => std_logic_vector(to_unsigned(1,8) ,
36846	 => std_logic_vector(to_unsigned(1,8) ,
36847	 => std_logic_vector(to_unsigned(2,8) ,
36848	 => std_logic_vector(to_unsigned(2,8) ,
36849	 => std_logic_vector(to_unsigned(2,8) ,
36850	 => std_logic_vector(to_unsigned(1,8) ,
36851	 => std_logic_vector(to_unsigned(0,8) ,
36852	 => std_logic_vector(to_unsigned(1,8) ,
36853	 => std_logic_vector(to_unsigned(1,8) ,
36854	 => std_logic_vector(to_unsigned(1,8) ,
36855	 => std_logic_vector(to_unsigned(2,8) ,
36856	 => std_logic_vector(to_unsigned(8,8) ,
36857	 => std_logic_vector(to_unsigned(9,8) ,
36858	 => std_logic_vector(to_unsigned(6,8) ,
36859	 => std_logic_vector(to_unsigned(8,8) ,
36860	 => std_logic_vector(to_unsigned(5,8) ,
36861	 => std_logic_vector(to_unsigned(3,8) ,
36862	 => std_logic_vector(to_unsigned(2,8) ,
36863	 => std_logic_vector(to_unsigned(2,8) ,
36864	 => std_logic_vector(to_unsigned(3,8) ,
36865	 => std_logic_vector(to_unsigned(4,8) ,
36866	 => std_logic_vector(to_unsigned(1,8) ,
36867	 => std_logic_vector(to_unsigned(0,8) ,
36868	 => std_logic_vector(to_unsigned(1,8) ,
36869	 => std_logic_vector(to_unsigned(1,8) ,
36870	 => std_logic_vector(to_unsigned(9,8) ,
36871	 => std_logic_vector(to_unsigned(32,8) ,
36872	 => std_logic_vector(to_unsigned(18,8) ,
36873	 => std_logic_vector(to_unsigned(6,8) ,
36874	 => std_logic_vector(to_unsigned(1,8) ,
36875	 => std_logic_vector(to_unsigned(0,8) ,
36876	 => std_logic_vector(to_unsigned(1,8) ,
36877	 => std_logic_vector(to_unsigned(9,8) ,
36878	 => std_logic_vector(to_unsigned(9,8) ,
36879	 => std_logic_vector(to_unsigned(4,8) ,
36880	 => std_logic_vector(to_unsigned(5,8) ,
36881	 => std_logic_vector(to_unsigned(5,8) ,
36882	 => std_logic_vector(to_unsigned(8,8) ,
36883	 => std_logic_vector(to_unsigned(6,8) ,
36884	 => std_logic_vector(to_unsigned(2,8) ,
36885	 => std_logic_vector(to_unsigned(2,8) ,
36886	 => std_logic_vector(to_unsigned(5,8) ,
36887	 => std_logic_vector(to_unsigned(1,8) ,
36888	 => std_logic_vector(to_unsigned(0,8) ,
36889	 => std_logic_vector(to_unsigned(0,8) ,
36890	 => std_logic_vector(to_unsigned(0,8) ,
36891	 => std_logic_vector(to_unsigned(0,8) ,
36892	 => std_logic_vector(to_unsigned(6,8) ,
36893	 => std_logic_vector(to_unsigned(13,8) ,
36894	 => std_logic_vector(to_unsigned(7,8) ,
36895	 => std_logic_vector(to_unsigned(10,8) ,
36896	 => std_logic_vector(to_unsigned(9,8) ,
36897	 => std_logic_vector(to_unsigned(7,8) ,
36898	 => std_logic_vector(to_unsigned(7,8) ,
36899	 => std_logic_vector(to_unsigned(2,8) ,
36900	 => std_logic_vector(to_unsigned(7,8) ,
36901	 => std_logic_vector(to_unsigned(17,8) ,
36902	 => std_logic_vector(to_unsigned(5,8) ,
36903	 => std_logic_vector(to_unsigned(5,8) ,
36904	 => std_logic_vector(to_unsigned(7,8) ,
36905	 => std_logic_vector(to_unsigned(6,8) ,
36906	 => std_logic_vector(to_unsigned(3,8) ,
36907	 => std_logic_vector(to_unsigned(1,8) ,
36908	 => std_logic_vector(to_unsigned(1,8) ,
36909	 => std_logic_vector(to_unsigned(2,8) ,
36910	 => std_logic_vector(to_unsigned(6,8) ,
36911	 => std_logic_vector(to_unsigned(111,8) ,
36912	 => std_logic_vector(to_unsigned(183,8) ,
36913	 => std_logic_vector(to_unsigned(147,8) ,
36914	 => std_logic_vector(to_unsigned(170,8) ,
36915	 => std_logic_vector(to_unsigned(70,8) ,
36916	 => std_logic_vector(to_unsigned(1,8) ,
36917	 => std_logic_vector(to_unsigned(0,8) ,
36918	 => std_logic_vector(to_unsigned(1,8) ,
36919	 => std_logic_vector(to_unsigned(0,8) ,
36920	 => std_logic_vector(to_unsigned(1,8) ,
36921	 => std_logic_vector(to_unsigned(0,8) ,
36922	 => std_logic_vector(to_unsigned(1,8) ,
36923	 => std_logic_vector(to_unsigned(4,8) ,
36924	 => std_logic_vector(to_unsigned(4,8) ,
36925	 => std_logic_vector(to_unsigned(8,8) ,
36926	 => std_logic_vector(to_unsigned(3,8) ,
36927	 => std_logic_vector(to_unsigned(4,8) ,
36928	 => std_logic_vector(to_unsigned(4,8) ,
36929	 => std_logic_vector(to_unsigned(2,8) ,
36930	 => std_logic_vector(to_unsigned(0,8) ,
36931	 => std_logic_vector(to_unsigned(2,8) ,
36932	 => std_logic_vector(to_unsigned(6,8) ,
36933	 => std_logic_vector(to_unsigned(4,8) ,
36934	 => std_logic_vector(to_unsigned(4,8) ,
36935	 => std_logic_vector(to_unsigned(4,8) ,
36936	 => std_logic_vector(to_unsigned(4,8) ,
36937	 => std_logic_vector(to_unsigned(2,8) ,
36938	 => std_logic_vector(to_unsigned(2,8) ,
36939	 => std_logic_vector(to_unsigned(2,8) ,
36940	 => std_logic_vector(to_unsigned(2,8) ,
36941	 => std_logic_vector(to_unsigned(1,8) ,
36942	 => std_logic_vector(to_unsigned(0,8) ,
36943	 => std_logic_vector(to_unsigned(1,8) ,
36944	 => std_logic_vector(to_unsigned(1,8) ,
36945	 => std_logic_vector(to_unsigned(1,8) ,
36946	 => std_logic_vector(to_unsigned(2,8) ,
36947	 => std_logic_vector(to_unsigned(2,8) ,
36948	 => std_logic_vector(to_unsigned(2,8) ,
36949	 => std_logic_vector(to_unsigned(2,8) ,
36950	 => std_logic_vector(to_unsigned(3,8) ,
36951	 => std_logic_vector(to_unsigned(3,8) ,
36952	 => std_logic_vector(to_unsigned(5,8) ,
36953	 => std_logic_vector(to_unsigned(5,8) ,
36954	 => std_logic_vector(to_unsigned(7,8) ,
36955	 => std_logic_vector(to_unsigned(12,8) ,
36956	 => std_logic_vector(to_unsigned(5,8) ,
36957	 => std_logic_vector(to_unsigned(2,8) ,
36958	 => std_logic_vector(to_unsigned(1,8) ,
36959	 => std_logic_vector(to_unsigned(3,8) ,
36960	 => std_logic_vector(to_unsigned(12,8) ,
36961	 => std_logic_vector(to_unsigned(5,8) ,
36962	 => std_logic_vector(to_unsigned(4,8) ,
36963	 => std_logic_vector(to_unsigned(3,8) ,
36964	 => std_logic_vector(to_unsigned(3,8) ,
36965	 => std_logic_vector(to_unsigned(6,8) ,
36966	 => std_logic_vector(to_unsigned(2,8) ,
36967	 => std_logic_vector(to_unsigned(0,8) ,
36968	 => std_logic_vector(to_unsigned(0,8) ,
36969	 => std_logic_vector(to_unsigned(0,8) ,
36970	 => std_logic_vector(to_unsigned(0,8) ,
36971	 => std_logic_vector(to_unsigned(0,8) ,
36972	 => std_logic_vector(to_unsigned(1,8) ,
36973	 => std_logic_vector(to_unsigned(1,8) ,
36974	 => std_logic_vector(to_unsigned(2,8) ,
36975	 => std_logic_vector(to_unsigned(2,8) ,
36976	 => std_logic_vector(to_unsigned(2,8) ,
36977	 => std_logic_vector(to_unsigned(5,8) ,
36978	 => std_logic_vector(to_unsigned(5,8) ,
36979	 => std_logic_vector(to_unsigned(6,8) ,
36980	 => std_logic_vector(to_unsigned(4,8) ,
36981	 => std_logic_vector(to_unsigned(0,8) ,
36982	 => std_logic_vector(to_unsigned(1,8) ,
36983	 => std_logic_vector(to_unsigned(4,8) ,
36984	 => std_logic_vector(to_unsigned(2,8) ,
36985	 => std_logic_vector(to_unsigned(3,8) ,
36986	 => std_logic_vector(to_unsigned(2,8) ,
36987	 => std_logic_vector(to_unsigned(2,8) ,
36988	 => std_logic_vector(to_unsigned(2,8) ,
36989	 => std_logic_vector(to_unsigned(2,8) ,
36990	 => std_logic_vector(to_unsigned(2,8) ,
36991	 => std_logic_vector(to_unsigned(0,8) ,
36992	 => std_logic_vector(to_unsigned(0,8) ,
36993	 => std_logic_vector(to_unsigned(0,8) ,
36994	 => std_logic_vector(to_unsigned(0,8) ,
36995	 => std_logic_vector(to_unsigned(0,8) ,
36996	 => std_logic_vector(to_unsigned(0,8) ,
36997	 => std_logic_vector(to_unsigned(0,8) ,
36998	 => std_logic_vector(to_unsigned(0,8) ,
36999	 => std_logic_vector(to_unsigned(0,8) ,
37000	 => std_logic_vector(to_unsigned(1,8) ,
37001	 => std_logic_vector(to_unsigned(1,8) ,
37002	 => std_logic_vector(to_unsigned(0,8) ,
37003	 => std_logic_vector(to_unsigned(0,8) ,
37004	 => std_logic_vector(to_unsigned(0,8) ,
37005	 => std_logic_vector(to_unsigned(1,8) ,
37006	 => std_logic_vector(to_unsigned(2,8) ,
37007	 => std_logic_vector(to_unsigned(2,8) ,
37008	 => std_logic_vector(to_unsigned(2,8) ,
37009	 => std_logic_vector(to_unsigned(3,8) ,
37010	 => std_logic_vector(to_unsigned(4,8) ,
37011	 => std_logic_vector(to_unsigned(6,8) ,
37012	 => std_logic_vector(to_unsigned(2,8) ,
37013	 => std_logic_vector(to_unsigned(11,8) ,
37014	 => std_logic_vector(to_unsigned(14,8) ,
37015	 => std_logic_vector(to_unsigned(11,8) ,
37016	 => std_logic_vector(to_unsigned(18,8) ,
37017	 => std_logic_vector(to_unsigned(26,8) ,
37018	 => std_logic_vector(to_unsigned(17,8) ,
37019	 => std_logic_vector(to_unsigned(13,8) ,
37020	 => std_logic_vector(to_unsigned(11,8) ,
37021	 => std_logic_vector(to_unsigned(8,8) ,
37022	 => std_logic_vector(to_unsigned(1,8) ,
37023	 => std_logic_vector(to_unsigned(1,8) ,
37024	 => std_logic_vector(to_unsigned(2,8) ,
37025	 => std_logic_vector(to_unsigned(2,8) ,
37026	 => std_logic_vector(to_unsigned(3,8) ,
37027	 => std_logic_vector(to_unsigned(3,8) ,
37028	 => std_logic_vector(to_unsigned(8,8) ,
37029	 => std_logic_vector(to_unsigned(15,8) ,
37030	 => std_logic_vector(to_unsigned(22,8) ,
37031	 => std_logic_vector(to_unsigned(69,8) ,
37032	 => std_logic_vector(to_unsigned(77,8) ,
37033	 => std_logic_vector(to_unsigned(44,8) ,
37034	 => std_logic_vector(to_unsigned(22,8) ,
37035	 => std_logic_vector(to_unsigned(7,8) ,
37036	 => std_logic_vector(to_unsigned(1,8) ,
37037	 => std_logic_vector(to_unsigned(3,8) ,
37038	 => std_logic_vector(to_unsigned(3,8) ,
37039	 => std_logic_vector(to_unsigned(2,8) ,
37040	 => std_logic_vector(to_unsigned(1,8) ,
37041	 => std_logic_vector(to_unsigned(1,8) ,
37042	 => std_logic_vector(to_unsigned(1,8) ,
37043	 => std_logic_vector(to_unsigned(1,8) ,
37044	 => std_logic_vector(to_unsigned(17,8) ,
37045	 => std_logic_vector(to_unsigned(26,8) ,
37046	 => std_logic_vector(to_unsigned(12,8) ,
37047	 => std_logic_vector(to_unsigned(1,8) ,
37048	 => std_logic_vector(to_unsigned(1,8) ,
37049	 => std_logic_vector(to_unsigned(2,8) ,
37050	 => std_logic_vector(to_unsigned(2,8) ,
37051	 => std_logic_vector(to_unsigned(1,8) ,
37052	 => std_logic_vector(to_unsigned(1,8) ,
37053	 => std_logic_vector(to_unsigned(1,8) ,
37054	 => std_logic_vector(to_unsigned(0,8) ,
37055	 => std_logic_vector(to_unsigned(0,8) ,
37056	 => std_logic_vector(to_unsigned(2,8) ,
37057	 => std_logic_vector(to_unsigned(2,8) ,
37058	 => std_logic_vector(to_unsigned(2,8) ,
37059	 => std_logic_vector(to_unsigned(3,8) ,
37060	 => std_logic_vector(to_unsigned(2,8) ,
37061	 => std_logic_vector(to_unsigned(6,8) ,
37062	 => std_logic_vector(to_unsigned(13,8) ,
37063	 => std_logic_vector(to_unsigned(22,8) ,
37064	 => std_logic_vector(to_unsigned(18,8) ,
37065	 => std_logic_vector(to_unsigned(23,8) ,
37066	 => std_logic_vector(to_unsigned(11,8) ,
37067	 => std_logic_vector(to_unsigned(11,8) ,
37068	 => std_logic_vector(to_unsigned(22,8) ,
37069	 => std_logic_vector(to_unsigned(76,8) ,
37070	 => std_logic_vector(to_unsigned(73,8) ,
37071	 => std_logic_vector(to_unsigned(40,8) ,
37072	 => std_logic_vector(to_unsigned(38,8) ,
37073	 => std_logic_vector(to_unsigned(38,8) ,
37074	 => std_logic_vector(to_unsigned(21,8) ,
37075	 => std_logic_vector(to_unsigned(3,8) ,
37076	 => std_logic_vector(to_unsigned(11,8) ,
37077	 => std_logic_vector(to_unsigned(20,8) ,
37078	 => std_logic_vector(to_unsigned(25,8) ,
37079	 => std_logic_vector(to_unsigned(5,8) ,
37080	 => std_logic_vector(to_unsigned(7,8) ,
37081	 => std_logic_vector(to_unsigned(8,8) ,
37082	 => std_logic_vector(to_unsigned(5,8) ,
37083	 => std_logic_vector(to_unsigned(12,8) ,
37084	 => std_logic_vector(to_unsigned(7,8) ,
37085	 => std_logic_vector(to_unsigned(4,8) ,
37086	 => std_logic_vector(to_unsigned(4,8) ,
37087	 => std_logic_vector(to_unsigned(17,8) ,
37088	 => std_logic_vector(to_unsigned(25,8) ,
37089	 => std_logic_vector(to_unsigned(17,8) ,
37090	 => std_logic_vector(to_unsigned(9,8) ,
37091	 => std_logic_vector(to_unsigned(12,8) ,
37092	 => std_logic_vector(to_unsigned(8,8) ,
37093	 => std_logic_vector(to_unsigned(11,8) ,
37094	 => std_logic_vector(to_unsigned(29,8) ,
37095	 => std_logic_vector(to_unsigned(63,8) ,
37096	 => std_logic_vector(to_unsigned(17,8) ,
37097	 => std_logic_vector(to_unsigned(2,8) ,
37098	 => std_logic_vector(to_unsigned(3,8) ,
37099	 => std_logic_vector(to_unsigned(3,8) ,
37100	 => std_logic_vector(to_unsigned(114,8) ,
37101	 => std_logic_vector(to_unsigned(175,8) ,
37102	 => std_logic_vector(to_unsigned(159,8) ,
37103	 => std_logic_vector(to_unsigned(161,8) ,
37104	 => std_logic_vector(to_unsigned(161,8) ,
37105	 => std_logic_vector(to_unsigned(156,8) ,
37106	 => std_logic_vector(to_unsigned(156,8) ,
37107	 => std_logic_vector(to_unsigned(159,8) ,
37108	 => std_logic_vector(to_unsigned(157,8) ,
37109	 => std_logic_vector(to_unsigned(159,8) ,
37110	 => std_logic_vector(to_unsigned(166,8) ,
37111	 => std_logic_vector(to_unsigned(159,8) ,
37112	 => std_logic_vector(to_unsigned(156,8) ,
37113	 => std_logic_vector(to_unsigned(157,8) ,
37114	 => std_logic_vector(to_unsigned(159,8) ,
37115	 => std_logic_vector(to_unsigned(161,8) ,
37116	 => std_logic_vector(to_unsigned(149,8) ,
37117	 => std_logic_vector(to_unsigned(139,8) ,
37118	 => std_logic_vector(to_unsigned(131,8) ,
37119	 => std_logic_vector(to_unsigned(128,8) ,
37120	 => std_logic_vector(to_unsigned(139,8) ,
37121	 => std_logic_vector(to_unsigned(136,8) ,
37122	 => std_logic_vector(to_unsigned(138,8) ,
37123	 => std_logic_vector(to_unsigned(141,8) ,
37124	 => std_logic_vector(to_unsigned(141,8) ,
37125	 => std_logic_vector(to_unsigned(157,8) ,
37126	 => std_logic_vector(to_unsigned(136,8) ,
37127	 => std_logic_vector(to_unsigned(16,8) ,
37128	 => std_logic_vector(to_unsigned(1,8) ,
37129	 => std_logic_vector(to_unsigned(1,8) ,
37130	 => std_logic_vector(to_unsigned(2,8) ,
37131	 => std_logic_vector(to_unsigned(8,8) ,
37132	 => std_logic_vector(to_unsigned(10,8) ,
37133	 => std_logic_vector(to_unsigned(31,8) ,
37134	 => std_logic_vector(to_unsigned(68,8) ,
37135	 => std_logic_vector(to_unsigned(10,8) ,
37136	 => std_logic_vector(to_unsigned(0,8) ,
37137	 => std_logic_vector(to_unsigned(3,8) ,
37138	 => std_logic_vector(to_unsigned(2,8) ,
37139	 => std_logic_vector(to_unsigned(0,8) ,
37140	 => std_logic_vector(to_unsigned(3,8) ,
37141	 => std_logic_vector(to_unsigned(3,8) ,
37142	 => std_logic_vector(to_unsigned(1,8) ,
37143	 => std_logic_vector(to_unsigned(1,8) ,
37144	 => std_logic_vector(to_unsigned(0,8) ,
37145	 => std_logic_vector(to_unsigned(0,8) ,
37146	 => std_logic_vector(to_unsigned(0,8) ,
37147	 => std_logic_vector(to_unsigned(0,8) ,
37148	 => std_logic_vector(to_unsigned(0,8) ,
37149	 => std_logic_vector(to_unsigned(0,8) ,
37150	 => std_logic_vector(to_unsigned(0,8) ,
37151	 => std_logic_vector(to_unsigned(6,8) ,
37152	 => std_logic_vector(to_unsigned(20,8) ,
37153	 => std_logic_vector(to_unsigned(7,8) ,
37154	 => std_logic_vector(to_unsigned(8,8) ,
37155	 => std_logic_vector(to_unsigned(5,8) ,
37156	 => std_logic_vector(to_unsigned(4,8) ,
37157	 => std_logic_vector(to_unsigned(3,8) ,
37158	 => std_logic_vector(to_unsigned(3,8) ,
37159	 => std_logic_vector(to_unsigned(3,8) ,
37160	 => std_logic_vector(to_unsigned(2,8) ,
37161	 => std_logic_vector(to_unsigned(8,8) ,
37162	 => std_logic_vector(to_unsigned(8,8) ,
37163	 => std_logic_vector(to_unsigned(6,8) ,
37164	 => std_logic_vector(to_unsigned(2,8) ,
37165	 => std_logic_vector(to_unsigned(1,8) ,
37166	 => std_logic_vector(to_unsigned(1,8) ,
37167	 => std_logic_vector(to_unsigned(2,8) ,
37168	 => std_logic_vector(to_unsigned(5,8) ,
37169	 => std_logic_vector(to_unsigned(4,8) ,
37170	 => std_logic_vector(to_unsigned(1,8) ,
37171	 => std_logic_vector(to_unsigned(1,8) ,
37172	 => std_logic_vector(to_unsigned(1,8) ,
37173	 => std_logic_vector(to_unsigned(1,8) ,
37174	 => std_logic_vector(to_unsigned(1,8) ,
37175	 => std_logic_vector(to_unsigned(1,8) ,
37176	 => std_logic_vector(to_unsigned(4,8) ,
37177	 => std_logic_vector(to_unsigned(7,8) ,
37178	 => std_logic_vector(to_unsigned(5,8) ,
37179	 => std_logic_vector(to_unsigned(4,8) ,
37180	 => std_logic_vector(to_unsigned(2,8) ,
37181	 => std_logic_vector(to_unsigned(2,8) ,
37182	 => std_logic_vector(to_unsigned(2,8) ,
37183	 => std_logic_vector(to_unsigned(2,8) ,
37184	 => std_logic_vector(to_unsigned(2,8) ,
37185	 => std_logic_vector(to_unsigned(2,8) ,
37186	 => std_logic_vector(to_unsigned(1,8) ,
37187	 => std_logic_vector(to_unsigned(0,8) ,
37188	 => std_logic_vector(to_unsigned(1,8) ,
37189	 => std_logic_vector(to_unsigned(1,8) ,
37190	 => std_logic_vector(to_unsigned(1,8) ,
37191	 => std_logic_vector(to_unsigned(15,8) ,
37192	 => std_logic_vector(to_unsigned(30,8) ,
37193	 => std_logic_vector(to_unsigned(15,8) ,
37194	 => std_logic_vector(to_unsigned(5,8) ,
37195	 => std_logic_vector(to_unsigned(1,8) ,
37196	 => std_logic_vector(to_unsigned(1,8) ,
37197	 => std_logic_vector(to_unsigned(10,8) ,
37198	 => std_logic_vector(to_unsigned(8,8) ,
37199	 => std_logic_vector(to_unsigned(3,8) ,
37200	 => std_logic_vector(to_unsigned(4,8) ,
37201	 => std_logic_vector(to_unsigned(5,8) ,
37202	 => std_logic_vector(to_unsigned(6,8) ,
37203	 => std_logic_vector(to_unsigned(4,8) ,
37204	 => std_logic_vector(to_unsigned(1,8) ,
37205	 => std_logic_vector(to_unsigned(3,8) ,
37206	 => std_logic_vector(to_unsigned(4,8) ,
37207	 => std_logic_vector(to_unsigned(0,8) ,
37208	 => std_logic_vector(to_unsigned(0,8) ,
37209	 => std_logic_vector(to_unsigned(0,8) ,
37210	 => std_logic_vector(to_unsigned(0,8) ,
37211	 => std_logic_vector(to_unsigned(0,8) ,
37212	 => std_logic_vector(to_unsigned(4,8) ,
37213	 => std_logic_vector(to_unsigned(12,8) ,
37214	 => std_logic_vector(to_unsigned(6,8) ,
37215	 => std_logic_vector(to_unsigned(8,8) ,
37216	 => std_logic_vector(to_unsigned(7,8) ,
37217	 => std_logic_vector(to_unsigned(6,8) ,
37218	 => std_logic_vector(to_unsigned(6,8) ,
37219	 => std_logic_vector(to_unsigned(2,8) ,
37220	 => std_logic_vector(to_unsigned(3,8) ,
37221	 => std_logic_vector(to_unsigned(7,8) ,
37222	 => std_logic_vector(to_unsigned(2,8) ,
37223	 => std_logic_vector(to_unsigned(8,8) ,
37224	 => std_logic_vector(to_unsigned(8,8) ,
37225	 => std_logic_vector(to_unsigned(5,8) ,
37226	 => std_logic_vector(to_unsigned(4,8) ,
37227	 => std_logic_vector(to_unsigned(2,8) ,
37228	 => std_logic_vector(to_unsigned(2,8) ,
37229	 => std_logic_vector(to_unsigned(2,8) ,
37230	 => std_logic_vector(to_unsigned(2,8) ,
37231	 => std_logic_vector(to_unsigned(27,8) ,
37232	 => std_logic_vector(to_unsigned(168,8) ,
37233	 => std_logic_vector(to_unsigned(157,8) ,
37234	 => std_logic_vector(to_unsigned(151,8) ,
37235	 => std_logic_vector(to_unsigned(170,8) ,
37236	 => std_logic_vector(to_unsigned(30,8) ,
37237	 => std_logic_vector(to_unsigned(0,8) ,
37238	 => std_logic_vector(to_unsigned(1,8) ,
37239	 => std_logic_vector(to_unsigned(1,8) ,
37240	 => std_logic_vector(to_unsigned(1,8) ,
37241	 => std_logic_vector(to_unsigned(0,8) ,
37242	 => std_logic_vector(to_unsigned(1,8) ,
37243	 => std_logic_vector(to_unsigned(3,8) ,
37244	 => std_logic_vector(to_unsigned(4,8) ,
37245	 => std_logic_vector(to_unsigned(9,8) ,
37246	 => std_logic_vector(to_unsigned(3,8) ,
37247	 => std_logic_vector(to_unsigned(2,8) ,
37248	 => std_logic_vector(to_unsigned(3,8) ,
37249	 => std_logic_vector(to_unsigned(1,8) ,
37250	 => std_logic_vector(to_unsigned(0,8) ,
37251	 => std_logic_vector(to_unsigned(3,8) ,
37252	 => std_logic_vector(to_unsigned(5,8) ,
37253	 => std_logic_vector(to_unsigned(4,8) ,
37254	 => std_logic_vector(to_unsigned(5,8) ,
37255	 => std_logic_vector(to_unsigned(5,8) ,
37256	 => std_logic_vector(to_unsigned(5,8) ,
37257	 => std_logic_vector(to_unsigned(3,8) ,
37258	 => std_logic_vector(to_unsigned(2,8) ,
37259	 => std_logic_vector(to_unsigned(3,8) ,
37260	 => std_logic_vector(to_unsigned(3,8) ,
37261	 => std_logic_vector(to_unsigned(3,8) ,
37262	 => std_logic_vector(to_unsigned(0,8) ,
37263	 => std_logic_vector(to_unsigned(0,8) ,
37264	 => std_logic_vector(to_unsigned(2,8) ,
37265	 => std_logic_vector(to_unsigned(2,8) ,
37266	 => std_logic_vector(to_unsigned(2,8) ,
37267	 => std_logic_vector(to_unsigned(3,8) ,
37268	 => std_logic_vector(to_unsigned(3,8) ,
37269	 => std_logic_vector(to_unsigned(3,8) ,
37270	 => std_logic_vector(to_unsigned(4,8) ,
37271	 => std_logic_vector(to_unsigned(3,8) ,
37272	 => std_logic_vector(to_unsigned(4,8) ,
37273	 => std_logic_vector(to_unsigned(5,8) ,
37274	 => std_logic_vector(to_unsigned(10,8) ,
37275	 => std_logic_vector(to_unsigned(12,8) ,
37276	 => std_logic_vector(to_unsigned(5,8) ,
37277	 => std_logic_vector(to_unsigned(1,8) ,
37278	 => std_logic_vector(to_unsigned(0,8) ,
37279	 => std_logic_vector(to_unsigned(3,8) ,
37280	 => std_logic_vector(to_unsigned(11,8) ,
37281	 => std_logic_vector(to_unsigned(9,8) ,
37282	 => std_logic_vector(to_unsigned(6,8) ,
37283	 => std_logic_vector(to_unsigned(3,8) ,
37284	 => std_logic_vector(to_unsigned(3,8) ,
37285	 => std_logic_vector(to_unsigned(4,8) ,
37286	 => std_logic_vector(to_unsigned(1,8) ,
37287	 => std_logic_vector(to_unsigned(0,8) ,
37288	 => std_logic_vector(to_unsigned(0,8) ,
37289	 => std_logic_vector(to_unsigned(1,8) ,
37290	 => std_logic_vector(to_unsigned(0,8) ,
37291	 => std_logic_vector(to_unsigned(1,8) ,
37292	 => std_logic_vector(to_unsigned(1,8) ,
37293	 => std_logic_vector(to_unsigned(1,8) ,
37294	 => std_logic_vector(to_unsigned(2,8) ,
37295	 => std_logic_vector(to_unsigned(2,8) ,
37296	 => std_logic_vector(to_unsigned(3,8) ,
37297	 => std_logic_vector(to_unsigned(6,8) ,
37298	 => std_logic_vector(to_unsigned(6,8) ,
37299	 => std_logic_vector(to_unsigned(6,8) ,
37300	 => std_logic_vector(to_unsigned(3,8) ,
37301	 => std_logic_vector(to_unsigned(0,8) ,
37302	 => std_logic_vector(to_unsigned(2,8) ,
37303	 => std_logic_vector(to_unsigned(6,8) ,
37304	 => std_logic_vector(to_unsigned(3,8) ,
37305	 => std_logic_vector(to_unsigned(3,8) ,
37306	 => std_logic_vector(to_unsigned(3,8) ,
37307	 => std_logic_vector(to_unsigned(2,8) ,
37308	 => std_logic_vector(to_unsigned(2,8) ,
37309	 => std_logic_vector(to_unsigned(2,8) ,
37310	 => std_logic_vector(to_unsigned(2,8) ,
37311	 => std_logic_vector(to_unsigned(0,8) ,
37312	 => std_logic_vector(to_unsigned(0,8) ,
37313	 => std_logic_vector(to_unsigned(0,8) ,
37314	 => std_logic_vector(to_unsigned(0,8) ,
37315	 => std_logic_vector(to_unsigned(0,8) ,
37316	 => std_logic_vector(to_unsigned(0,8) ,
37317	 => std_logic_vector(to_unsigned(1,8) ,
37318	 => std_logic_vector(to_unsigned(1,8) ,
37319	 => std_logic_vector(to_unsigned(1,8) ,
37320	 => std_logic_vector(to_unsigned(1,8) ,
37321	 => std_logic_vector(to_unsigned(2,8) ,
37322	 => std_logic_vector(to_unsigned(1,8) ,
37323	 => std_logic_vector(to_unsigned(1,8) ,
37324	 => std_logic_vector(to_unsigned(1,8) ,
37325	 => std_logic_vector(to_unsigned(1,8) ,
37326	 => std_logic_vector(to_unsigned(2,8) ,
37327	 => std_logic_vector(to_unsigned(2,8) ,
37328	 => std_logic_vector(to_unsigned(1,8) ,
37329	 => std_logic_vector(to_unsigned(2,8) ,
37330	 => std_logic_vector(to_unsigned(3,8) ,
37331	 => std_logic_vector(to_unsigned(4,8) ,
37332	 => std_logic_vector(to_unsigned(2,8) ,
37333	 => std_logic_vector(to_unsigned(8,8) ,
37334	 => std_logic_vector(to_unsigned(13,8) ,
37335	 => std_logic_vector(to_unsigned(17,8) ,
37336	 => std_logic_vector(to_unsigned(37,8) ,
37337	 => std_logic_vector(to_unsigned(31,8) ,
37338	 => std_logic_vector(to_unsigned(30,8) ,
37339	 => std_logic_vector(to_unsigned(32,8) ,
37340	 => std_logic_vector(to_unsigned(20,8) ,
37341	 => std_logic_vector(to_unsigned(8,8) ,
37342	 => std_logic_vector(to_unsigned(1,8) ,
37343	 => std_logic_vector(to_unsigned(0,8) ,
37344	 => std_logic_vector(to_unsigned(1,8) ,
37345	 => std_logic_vector(to_unsigned(1,8) ,
37346	 => std_logic_vector(to_unsigned(1,8) ,
37347	 => std_logic_vector(to_unsigned(1,8) ,
37348	 => std_logic_vector(to_unsigned(1,8) ,
37349	 => std_logic_vector(to_unsigned(8,8) ,
37350	 => std_logic_vector(to_unsigned(32,8) ,
37351	 => std_logic_vector(to_unsigned(85,8) ,
37352	 => std_logic_vector(to_unsigned(86,8) ,
37353	 => std_logic_vector(to_unsigned(45,8) ,
37354	 => std_logic_vector(to_unsigned(20,8) ,
37355	 => std_logic_vector(to_unsigned(7,8) ,
37356	 => std_logic_vector(to_unsigned(2,8) ,
37357	 => std_logic_vector(to_unsigned(2,8) ,
37358	 => std_logic_vector(to_unsigned(2,8) ,
37359	 => std_logic_vector(to_unsigned(1,8) ,
37360	 => std_logic_vector(to_unsigned(2,8) ,
37361	 => std_logic_vector(to_unsigned(1,8) ,
37362	 => std_logic_vector(to_unsigned(1,8) ,
37363	 => std_logic_vector(to_unsigned(1,8) ,
37364	 => std_logic_vector(to_unsigned(14,8) ,
37365	 => std_logic_vector(to_unsigned(41,8) ,
37366	 => std_logic_vector(to_unsigned(23,8) ,
37367	 => std_logic_vector(to_unsigned(1,8) ,
37368	 => std_logic_vector(to_unsigned(1,8) ,
37369	 => std_logic_vector(to_unsigned(1,8) ,
37370	 => std_logic_vector(to_unsigned(1,8) ,
37371	 => std_logic_vector(to_unsigned(1,8) ,
37372	 => std_logic_vector(to_unsigned(1,8) ,
37373	 => std_logic_vector(to_unsigned(1,8) ,
37374	 => std_logic_vector(to_unsigned(1,8) ,
37375	 => std_logic_vector(to_unsigned(0,8) ,
37376	 => std_logic_vector(to_unsigned(2,8) ,
37377	 => std_logic_vector(to_unsigned(4,8) ,
37378	 => std_logic_vector(to_unsigned(4,8) ,
37379	 => std_logic_vector(to_unsigned(3,8) ,
37380	 => std_logic_vector(to_unsigned(2,8) ,
37381	 => std_logic_vector(to_unsigned(7,8) ,
37382	 => std_logic_vector(to_unsigned(13,8) ,
37383	 => std_logic_vector(to_unsigned(10,8) ,
37384	 => std_logic_vector(to_unsigned(6,8) ,
37385	 => std_logic_vector(to_unsigned(18,8) ,
37386	 => std_logic_vector(to_unsigned(21,8) ,
37387	 => std_logic_vector(to_unsigned(9,8) ,
37388	 => std_logic_vector(to_unsigned(15,8) ,
37389	 => std_logic_vector(to_unsigned(52,8) ,
37390	 => std_logic_vector(to_unsigned(58,8) ,
37391	 => std_logic_vector(to_unsigned(32,8) ,
37392	 => std_logic_vector(to_unsigned(40,8) ,
37393	 => std_logic_vector(to_unsigned(24,8) ,
37394	 => std_logic_vector(to_unsigned(33,8) ,
37395	 => std_logic_vector(to_unsigned(20,8) ,
37396	 => std_logic_vector(to_unsigned(12,8) ,
37397	 => std_logic_vector(to_unsigned(17,8) ,
37398	 => std_logic_vector(to_unsigned(25,8) ,
37399	 => std_logic_vector(to_unsigned(10,8) ,
37400	 => std_logic_vector(to_unsigned(3,8) ,
37401	 => std_logic_vector(to_unsigned(7,8) ,
37402	 => std_logic_vector(to_unsigned(3,8) ,
37403	 => std_logic_vector(to_unsigned(5,8) ,
37404	 => std_logic_vector(to_unsigned(3,8) ,
37405	 => std_logic_vector(to_unsigned(1,8) ,
37406	 => std_logic_vector(to_unsigned(6,8) ,
37407	 => std_logic_vector(to_unsigned(49,8) ,
37408	 => std_logic_vector(to_unsigned(85,8) ,
37409	 => std_logic_vector(to_unsigned(55,8) ,
37410	 => std_logic_vector(to_unsigned(24,8) ,
37411	 => std_logic_vector(to_unsigned(8,8) ,
37412	 => std_logic_vector(to_unsigned(10,8) ,
37413	 => std_logic_vector(to_unsigned(16,8) ,
37414	 => std_logic_vector(to_unsigned(8,8) ,
37415	 => std_logic_vector(to_unsigned(46,8) ,
37416	 => std_logic_vector(to_unsigned(23,8) ,
37417	 => std_logic_vector(to_unsigned(2,8) ,
37418	 => std_logic_vector(to_unsigned(1,8) ,
37419	 => std_logic_vector(to_unsigned(12,8) ,
37420	 => std_logic_vector(to_unsigned(119,8) ,
37421	 => std_logic_vector(to_unsigned(122,8) ,
37422	 => std_logic_vector(to_unsigned(131,8) ,
37423	 => std_logic_vector(to_unsigned(136,8) ,
37424	 => std_logic_vector(to_unsigned(152,8) ,
37425	 => std_logic_vector(to_unsigned(163,8) ,
37426	 => std_logic_vector(to_unsigned(164,8) ,
37427	 => std_logic_vector(to_unsigned(163,8) ,
37428	 => std_logic_vector(to_unsigned(166,8) ,
37429	 => std_logic_vector(to_unsigned(179,8) ,
37430	 => std_logic_vector(to_unsigned(175,8) ,
37431	 => std_logic_vector(to_unsigned(166,8) ,
37432	 => std_logic_vector(to_unsigned(173,8) ,
37433	 => std_logic_vector(to_unsigned(171,8) ,
37434	 => std_logic_vector(to_unsigned(168,8) ,
37435	 => std_logic_vector(to_unsigned(171,8) ,
37436	 => std_logic_vector(to_unsigned(170,8) ,
37437	 => std_logic_vector(to_unsigned(164,8) ,
37438	 => std_logic_vector(to_unsigned(157,8) ,
37439	 => std_logic_vector(to_unsigned(157,8) ,
37440	 => std_logic_vector(to_unsigned(156,8) ,
37441	 => std_logic_vector(to_unsigned(131,8) ,
37442	 => std_logic_vector(to_unsigned(133,8) ,
37443	 => std_logic_vector(to_unsigned(125,8) ,
37444	 => std_logic_vector(to_unsigned(130,8) ,
37445	 => std_logic_vector(to_unsigned(128,8) ,
37446	 => std_logic_vector(to_unsigned(144,8) ,
37447	 => std_logic_vector(to_unsigned(112,8) ,
37448	 => std_logic_vector(to_unsigned(50,8) ,
37449	 => std_logic_vector(to_unsigned(42,8) ,
37450	 => std_logic_vector(to_unsigned(82,8) ,
37451	 => std_logic_vector(to_unsigned(124,8) ,
37452	 => std_logic_vector(to_unsigned(124,8) ,
37453	 => std_logic_vector(to_unsigned(142,8) ,
37454	 => std_logic_vector(to_unsigned(168,8) ,
37455	 => std_logic_vector(to_unsigned(52,8) ,
37456	 => std_logic_vector(to_unsigned(1,8) ,
37457	 => std_logic_vector(to_unsigned(6,8) ,
37458	 => std_logic_vector(to_unsigned(3,8) ,
37459	 => std_logic_vector(to_unsigned(1,8) ,
37460	 => std_logic_vector(to_unsigned(69,8) ,
37461	 => std_logic_vector(to_unsigned(127,8) ,
37462	 => std_logic_vector(to_unsigned(82,8) ,
37463	 => std_logic_vector(to_unsigned(73,8) ,
37464	 => std_logic_vector(to_unsigned(58,8) ,
37465	 => std_logic_vector(to_unsigned(44,8) ,
37466	 => std_logic_vector(to_unsigned(35,8) ,
37467	 => std_logic_vector(to_unsigned(23,8) ,
37468	 => std_logic_vector(to_unsigned(13,8) ,
37469	 => std_logic_vector(to_unsigned(6,8) ,
37470	 => std_logic_vector(to_unsigned(4,8) ,
37471	 => std_logic_vector(to_unsigned(8,8) ,
37472	 => std_logic_vector(to_unsigned(13,8) ,
37473	 => std_logic_vector(to_unsigned(4,8) ,
37474	 => std_logic_vector(to_unsigned(3,8) ,
37475	 => std_logic_vector(to_unsigned(6,8) ,
37476	 => std_logic_vector(to_unsigned(4,8) ,
37477	 => std_logic_vector(to_unsigned(4,8) ,
37478	 => std_logic_vector(to_unsigned(5,8) ,
37479	 => std_logic_vector(to_unsigned(3,8) ,
37480	 => std_logic_vector(to_unsigned(3,8) ,
37481	 => std_logic_vector(to_unsigned(9,8) ,
37482	 => std_logic_vector(to_unsigned(11,8) ,
37483	 => std_logic_vector(to_unsigned(8,8) ,
37484	 => std_logic_vector(to_unsigned(1,8) ,
37485	 => std_logic_vector(to_unsigned(0,8) ,
37486	 => std_logic_vector(to_unsigned(2,8) ,
37487	 => std_logic_vector(to_unsigned(8,8) ,
37488	 => std_logic_vector(to_unsigned(8,8) ,
37489	 => std_logic_vector(to_unsigned(1,8) ,
37490	 => std_logic_vector(to_unsigned(0,8) ,
37491	 => std_logic_vector(to_unsigned(1,8) ,
37492	 => std_logic_vector(to_unsigned(1,8) ,
37493	 => std_logic_vector(to_unsigned(2,8) ,
37494	 => std_logic_vector(to_unsigned(2,8) ,
37495	 => std_logic_vector(to_unsigned(2,8) ,
37496	 => std_logic_vector(to_unsigned(3,8) ,
37497	 => std_logic_vector(to_unsigned(7,8) ,
37498	 => std_logic_vector(to_unsigned(7,8) ,
37499	 => std_logic_vector(to_unsigned(3,8) ,
37500	 => std_logic_vector(to_unsigned(5,8) ,
37501	 => std_logic_vector(to_unsigned(4,8) ,
37502	 => std_logic_vector(to_unsigned(3,8) ,
37503	 => std_logic_vector(to_unsigned(3,8) ,
37504	 => std_logic_vector(to_unsigned(2,8) ,
37505	 => std_logic_vector(to_unsigned(2,8) ,
37506	 => std_logic_vector(to_unsigned(1,8) ,
37507	 => std_logic_vector(to_unsigned(0,8) ,
37508	 => std_logic_vector(to_unsigned(2,8) ,
37509	 => std_logic_vector(to_unsigned(6,8) ,
37510	 => std_logic_vector(to_unsigned(1,8) ,
37511	 => std_logic_vector(to_unsigned(1,8) ,
37512	 => std_logic_vector(to_unsigned(6,8) ,
37513	 => std_logic_vector(to_unsigned(5,8) ,
37514	 => std_logic_vector(to_unsigned(3,8) ,
37515	 => std_logic_vector(to_unsigned(1,8) ,
37516	 => std_logic_vector(to_unsigned(1,8) ,
37517	 => std_logic_vector(to_unsigned(9,8) ,
37518	 => std_logic_vector(to_unsigned(8,8) ,
37519	 => std_logic_vector(to_unsigned(4,8) ,
37520	 => std_logic_vector(to_unsigned(4,8) ,
37521	 => std_logic_vector(to_unsigned(5,8) ,
37522	 => std_logic_vector(to_unsigned(6,8) ,
37523	 => std_logic_vector(to_unsigned(2,8) ,
37524	 => std_logic_vector(to_unsigned(2,8) ,
37525	 => std_logic_vector(to_unsigned(8,8) ,
37526	 => std_logic_vector(to_unsigned(3,8) ,
37527	 => std_logic_vector(to_unsigned(0,8) ,
37528	 => std_logic_vector(to_unsigned(0,8) ,
37529	 => std_logic_vector(to_unsigned(0,8) ,
37530	 => std_logic_vector(to_unsigned(0,8) ,
37531	 => std_logic_vector(to_unsigned(0,8) ,
37532	 => std_logic_vector(to_unsigned(3,8) ,
37533	 => std_logic_vector(to_unsigned(14,8) ,
37534	 => std_logic_vector(to_unsigned(7,8) ,
37535	 => std_logic_vector(to_unsigned(6,8) ,
37536	 => std_logic_vector(to_unsigned(6,8) ,
37537	 => std_logic_vector(to_unsigned(6,8) ,
37538	 => std_logic_vector(to_unsigned(7,8) ,
37539	 => std_logic_vector(to_unsigned(2,8) ,
37540	 => std_logic_vector(to_unsigned(2,8) ,
37541	 => std_logic_vector(to_unsigned(4,8) ,
37542	 => std_logic_vector(to_unsigned(2,8) ,
37543	 => std_logic_vector(to_unsigned(9,8) ,
37544	 => std_logic_vector(to_unsigned(7,8) ,
37545	 => std_logic_vector(to_unsigned(4,8) ,
37546	 => std_logic_vector(to_unsigned(5,8) ,
37547	 => std_logic_vector(to_unsigned(3,8) ,
37548	 => std_logic_vector(to_unsigned(2,8) ,
37549	 => std_logic_vector(to_unsigned(2,8) ,
37550	 => std_logic_vector(to_unsigned(1,8) ,
37551	 => std_logic_vector(to_unsigned(1,8) ,
37552	 => std_logic_vector(to_unsigned(71,8) ,
37553	 => std_logic_vector(to_unsigned(175,8) ,
37554	 => std_logic_vector(to_unsigned(144,8) ,
37555	 => std_logic_vector(to_unsigned(159,8) ,
37556	 => std_logic_vector(to_unsigned(133,8) ,
37557	 => std_logic_vector(to_unsigned(12,8) ,
37558	 => std_logic_vector(to_unsigned(0,8) ,
37559	 => std_logic_vector(to_unsigned(1,8) ,
37560	 => std_logic_vector(to_unsigned(1,8) ,
37561	 => std_logic_vector(to_unsigned(0,8) ,
37562	 => std_logic_vector(to_unsigned(1,8) ,
37563	 => std_logic_vector(to_unsigned(3,8) ,
37564	 => std_logic_vector(to_unsigned(6,8) ,
37565	 => std_logic_vector(to_unsigned(8,8) ,
37566	 => std_logic_vector(to_unsigned(3,8) ,
37567	 => std_logic_vector(to_unsigned(2,8) ,
37568	 => std_logic_vector(to_unsigned(3,8) ,
37569	 => std_logic_vector(to_unsigned(2,8) ,
37570	 => std_logic_vector(to_unsigned(0,8) ,
37571	 => std_logic_vector(to_unsigned(3,8) ,
37572	 => std_logic_vector(to_unsigned(7,8) ,
37573	 => std_logic_vector(to_unsigned(4,8) ,
37574	 => std_logic_vector(to_unsigned(4,8) ,
37575	 => std_logic_vector(to_unsigned(4,8) ,
37576	 => std_logic_vector(to_unsigned(4,8) ,
37577	 => std_logic_vector(to_unsigned(5,8) ,
37578	 => std_logic_vector(to_unsigned(4,8) ,
37579	 => std_logic_vector(to_unsigned(2,8) ,
37580	 => std_logic_vector(to_unsigned(3,8) ,
37581	 => std_logic_vector(to_unsigned(4,8) ,
37582	 => std_logic_vector(to_unsigned(1,8) ,
37583	 => std_logic_vector(to_unsigned(0,8) ,
37584	 => std_logic_vector(to_unsigned(1,8) ,
37585	 => std_logic_vector(to_unsigned(1,8) ,
37586	 => std_logic_vector(to_unsigned(2,8) ,
37587	 => std_logic_vector(to_unsigned(3,8) ,
37588	 => std_logic_vector(to_unsigned(3,8) ,
37589	 => std_logic_vector(to_unsigned(4,8) ,
37590	 => std_logic_vector(to_unsigned(4,8) ,
37591	 => std_logic_vector(to_unsigned(3,8) ,
37592	 => std_logic_vector(to_unsigned(3,8) ,
37593	 => std_logic_vector(to_unsigned(7,8) ,
37594	 => std_logic_vector(to_unsigned(11,8) ,
37595	 => std_logic_vector(to_unsigned(10,8) ,
37596	 => std_logic_vector(to_unsigned(5,8) ,
37597	 => std_logic_vector(to_unsigned(1,8) ,
37598	 => std_logic_vector(to_unsigned(0,8) ,
37599	 => std_logic_vector(to_unsigned(4,8) ,
37600	 => std_logic_vector(to_unsigned(10,8) ,
37601	 => std_logic_vector(to_unsigned(8,8) ,
37602	 => std_logic_vector(to_unsigned(7,8) ,
37603	 => std_logic_vector(to_unsigned(4,8) ,
37604	 => std_logic_vector(to_unsigned(2,8) ,
37605	 => std_logic_vector(to_unsigned(4,8) ,
37606	 => std_logic_vector(to_unsigned(1,8) ,
37607	 => std_logic_vector(to_unsigned(0,8) ,
37608	 => std_logic_vector(to_unsigned(0,8) ,
37609	 => std_logic_vector(to_unsigned(0,8) ,
37610	 => std_logic_vector(to_unsigned(1,8) ,
37611	 => std_logic_vector(to_unsigned(1,8) ,
37612	 => std_logic_vector(to_unsigned(1,8) ,
37613	 => std_logic_vector(to_unsigned(1,8) ,
37614	 => std_logic_vector(to_unsigned(2,8) ,
37615	 => std_logic_vector(to_unsigned(1,8) ,
37616	 => std_logic_vector(to_unsigned(4,8) ,
37617	 => std_logic_vector(to_unsigned(9,8) ,
37618	 => std_logic_vector(to_unsigned(6,8) ,
37619	 => std_logic_vector(to_unsigned(7,8) ,
37620	 => std_logic_vector(to_unsigned(3,8) ,
37621	 => std_logic_vector(to_unsigned(0,8) ,
37622	 => std_logic_vector(to_unsigned(2,8) ,
37623	 => std_logic_vector(to_unsigned(7,8) ,
37624	 => std_logic_vector(to_unsigned(4,8) ,
37625	 => std_logic_vector(to_unsigned(3,8) ,
37626	 => std_logic_vector(to_unsigned(3,8) ,
37627	 => std_logic_vector(to_unsigned(2,8) ,
37628	 => std_logic_vector(to_unsigned(2,8) ,
37629	 => std_logic_vector(to_unsigned(2,8) ,
37630	 => std_logic_vector(to_unsigned(1,8) ,
37631	 => std_logic_vector(to_unsigned(0,8) ,
37632	 => std_logic_vector(to_unsigned(0,8) ,
37633	 => std_logic_vector(to_unsigned(0,8) ,
37634	 => std_logic_vector(to_unsigned(0,8) ,
37635	 => std_logic_vector(to_unsigned(0,8) ,
37636	 => std_logic_vector(to_unsigned(0,8) ,
37637	 => std_logic_vector(to_unsigned(1,8) ,
37638	 => std_logic_vector(to_unsigned(1,8) ,
37639	 => std_logic_vector(to_unsigned(1,8) ,
37640	 => std_logic_vector(to_unsigned(0,8) ,
37641	 => std_logic_vector(to_unsigned(1,8) ,
37642	 => std_logic_vector(to_unsigned(1,8) ,
37643	 => std_logic_vector(to_unsigned(1,8) ,
37644	 => std_logic_vector(to_unsigned(1,8) ,
37645	 => std_logic_vector(to_unsigned(1,8) ,
37646	 => std_logic_vector(to_unsigned(2,8) ,
37647	 => std_logic_vector(to_unsigned(2,8) ,
37648	 => std_logic_vector(to_unsigned(2,8) ,
37649	 => std_logic_vector(to_unsigned(2,8) ,
37650	 => std_logic_vector(to_unsigned(3,8) ,
37651	 => std_logic_vector(to_unsigned(5,8) ,
37652	 => std_logic_vector(to_unsigned(1,8) ,
37653	 => std_logic_vector(to_unsigned(8,8) ,
37654	 => std_logic_vector(to_unsigned(14,8) ,
37655	 => std_logic_vector(to_unsigned(19,8) ,
37656	 => std_logic_vector(to_unsigned(41,8) ,
37657	 => std_logic_vector(to_unsigned(35,8) ,
37658	 => std_logic_vector(to_unsigned(35,8) ,
37659	 => std_logic_vector(to_unsigned(25,8) ,
37660	 => std_logic_vector(to_unsigned(23,8) ,
37661	 => std_logic_vector(to_unsigned(8,8) ,
37662	 => std_logic_vector(to_unsigned(0,8) ,
37663	 => std_logic_vector(to_unsigned(0,8) ,
37664	 => std_logic_vector(to_unsigned(0,8) ,
37665	 => std_logic_vector(to_unsigned(0,8) ,
37666	 => std_logic_vector(to_unsigned(0,8) ,
37667	 => std_logic_vector(to_unsigned(1,8) ,
37668	 => std_logic_vector(to_unsigned(0,8) ,
37669	 => std_logic_vector(to_unsigned(8,8) ,
37670	 => std_logic_vector(to_unsigned(62,8) ,
37671	 => std_logic_vector(to_unsigned(91,8) ,
37672	 => std_logic_vector(to_unsigned(73,8) ,
37673	 => std_logic_vector(to_unsigned(42,8) ,
37674	 => std_logic_vector(to_unsigned(29,8) ,
37675	 => std_logic_vector(to_unsigned(13,8) ,
37676	 => std_logic_vector(to_unsigned(3,8) ,
37677	 => std_logic_vector(to_unsigned(2,8) ,
37678	 => std_logic_vector(to_unsigned(2,8) ,
37679	 => std_logic_vector(to_unsigned(2,8) ,
37680	 => std_logic_vector(to_unsigned(2,8) ,
37681	 => std_logic_vector(to_unsigned(1,8) ,
37682	 => std_logic_vector(to_unsigned(2,8) ,
37683	 => std_logic_vector(to_unsigned(1,8) ,
37684	 => std_logic_vector(to_unsigned(8,8) ,
37685	 => std_logic_vector(to_unsigned(43,8) ,
37686	 => std_logic_vector(to_unsigned(30,8) ,
37687	 => std_logic_vector(to_unsigned(3,8) ,
37688	 => std_logic_vector(to_unsigned(1,8) ,
37689	 => std_logic_vector(to_unsigned(3,8) ,
37690	 => std_logic_vector(to_unsigned(4,8) ,
37691	 => std_logic_vector(to_unsigned(5,8) ,
37692	 => std_logic_vector(to_unsigned(5,8) ,
37693	 => std_logic_vector(to_unsigned(5,8) ,
37694	 => std_logic_vector(to_unsigned(4,8) ,
37695	 => std_logic_vector(to_unsigned(3,8) ,
37696	 => std_logic_vector(to_unsigned(4,8) ,
37697	 => std_logic_vector(to_unsigned(4,8) ,
37698	 => std_logic_vector(to_unsigned(4,8) ,
37699	 => std_logic_vector(to_unsigned(3,8) ,
37700	 => std_logic_vector(to_unsigned(3,8) ,
37701	 => std_logic_vector(to_unsigned(8,8) ,
37702	 => std_logic_vector(to_unsigned(11,8) ,
37703	 => std_logic_vector(to_unsigned(6,8) ,
37704	 => std_logic_vector(to_unsigned(10,8) ,
37705	 => std_logic_vector(to_unsigned(38,8) ,
37706	 => std_logic_vector(to_unsigned(29,8) ,
37707	 => std_logic_vector(to_unsigned(7,8) ,
37708	 => std_logic_vector(to_unsigned(13,8) ,
37709	 => std_logic_vector(to_unsigned(41,8) ,
37710	 => std_logic_vector(to_unsigned(65,8) ,
37711	 => std_logic_vector(to_unsigned(60,8) ,
37712	 => std_logic_vector(to_unsigned(42,8) ,
37713	 => std_logic_vector(to_unsigned(34,8) ,
37714	 => std_logic_vector(to_unsigned(27,8) ,
37715	 => std_logic_vector(to_unsigned(17,8) ,
37716	 => std_logic_vector(to_unsigned(13,8) ,
37717	 => std_logic_vector(to_unsigned(14,8) ,
37718	 => std_logic_vector(to_unsigned(17,8) ,
37719	 => std_logic_vector(to_unsigned(17,8) ,
37720	 => std_logic_vector(to_unsigned(7,8) ,
37721	 => std_logic_vector(to_unsigned(6,8) ,
37722	 => std_logic_vector(to_unsigned(2,8) ,
37723	 => std_logic_vector(to_unsigned(1,8) ,
37724	 => std_logic_vector(to_unsigned(4,8) ,
37725	 => std_logic_vector(to_unsigned(2,8) ,
37726	 => std_logic_vector(to_unsigned(13,8) ,
37727	 => std_logic_vector(to_unsigned(108,8) ,
37728	 => std_logic_vector(to_unsigned(119,8) ,
37729	 => std_logic_vector(to_unsigned(80,8) ,
37730	 => std_logic_vector(to_unsigned(51,8) ,
37731	 => std_logic_vector(to_unsigned(12,8) ,
37732	 => std_logic_vector(to_unsigned(2,8) ,
37733	 => std_logic_vector(to_unsigned(4,8) ,
37734	 => std_logic_vector(to_unsigned(9,8) ,
37735	 => std_logic_vector(to_unsigned(14,8) ,
37736	 => std_logic_vector(to_unsigned(7,8) ,
37737	 => std_logic_vector(to_unsigned(3,8) ,
37738	 => std_logic_vector(to_unsigned(1,8) ,
37739	 => std_logic_vector(to_unsigned(2,8) ,
37740	 => std_logic_vector(to_unsigned(5,8) ,
37741	 => std_logic_vector(to_unsigned(5,8) ,
37742	 => std_logic_vector(to_unsigned(8,8) ,
37743	 => std_logic_vector(to_unsigned(13,8) ,
37744	 => std_logic_vector(to_unsigned(20,8) ,
37745	 => std_logic_vector(to_unsigned(32,8) ,
37746	 => std_logic_vector(to_unsigned(45,8) ,
37747	 => std_logic_vector(to_unsigned(53,8) ,
37748	 => std_logic_vector(to_unsigned(72,8) ,
37749	 => std_logic_vector(to_unsigned(96,8) ,
37750	 => std_logic_vector(to_unsigned(105,8) ,
37751	 => std_logic_vector(to_unsigned(127,8) ,
37752	 => std_logic_vector(to_unsigned(144,8) ,
37753	 => std_logic_vector(to_unsigned(152,8) ,
37754	 => std_logic_vector(to_unsigned(161,8) ,
37755	 => std_logic_vector(to_unsigned(168,8) ,
37756	 => std_logic_vector(to_unsigned(171,8) ,
37757	 => std_logic_vector(to_unsigned(177,8) ,
37758	 => std_logic_vector(to_unsigned(177,8) ,
37759	 => std_logic_vector(to_unsigned(184,8) ,
37760	 => std_logic_vector(to_unsigned(184,8) ,
37761	 => std_logic_vector(to_unsigned(136,8) ,
37762	 => std_logic_vector(to_unsigned(141,8) ,
37763	 => std_logic_vector(to_unsigned(142,8) ,
37764	 => std_logic_vector(to_unsigned(142,8) ,
37765	 => std_logic_vector(to_unsigned(139,8) ,
37766	 => std_logic_vector(to_unsigned(130,8) ,
37767	 => std_logic_vector(to_unsigned(142,8) ,
37768	 => std_logic_vector(to_unsigned(156,8) ,
37769	 => std_logic_vector(to_unsigned(154,8) ,
37770	 => std_logic_vector(to_unsigned(156,8) ,
37771	 => std_logic_vector(to_unsigned(149,8) ,
37772	 => std_logic_vector(to_unsigned(141,8) ,
37773	 => std_logic_vector(to_unsigned(136,8) ,
37774	 => std_logic_vector(to_unsigned(154,8) ,
37775	 => std_logic_vector(to_unsigned(52,8) ,
37776	 => std_logic_vector(to_unsigned(1,8) ,
37777	 => std_logic_vector(to_unsigned(8,8) ,
37778	 => std_logic_vector(to_unsigned(5,8) ,
37779	 => std_logic_vector(to_unsigned(1,8) ,
37780	 => std_logic_vector(to_unsigned(76,8) ,
37781	 => std_logic_vector(to_unsigned(192,8) ,
37782	 => std_logic_vector(to_unsigned(157,8) ,
37783	 => std_logic_vector(to_unsigned(168,8) ,
37784	 => std_logic_vector(to_unsigned(166,8) ,
37785	 => std_logic_vector(to_unsigned(163,8) ,
37786	 => std_logic_vector(to_unsigned(168,8) ,
37787	 => std_logic_vector(to_unsigned(166,8) ,
37788	 => std_logic_vector(to_unsigned(141,8) ,
37789	 => std_logic_vector(to_unsigned(133,8) ,
37790	 => std_logic_vector(to_unsigned(86,8) ,
37791	 => std_logic_vector(to_unsigned(8,8) ,
37792	 => std_logic_vector(to_unsigned(6,8) ,
37793	 => std_logic_vector(to_unsigned(9,8) ,
37794	 => std_logic_vector(to_unsigned(8,8) ,
37795	 => std_logic_vector(to_unsigned(7,8) ,
37796	 => std_logic_vector(to_unsigned(8,8) ,
37797	 => std_logic_vector(to_unsigned(6,8) ,
37798	 => std_logic_vector(to_unsigned(5,8) ,
37799	 => std_logic_vector(to_unsigned(4,8) ,
37800	 => std_logic_vector(to_unsigned(5,8) ,
37801	 => std_logic_vector(to_unsigned(8,8) ,
37802	 => std_logic_vector(to_unsigned(10,8) ,
37803	 => std_logic_vector(to_unsigned(4,8) ,
37804	 => std_logic_vector(to_unsigned(0,8) ,
37805	 => std_logic_vector(to_unsigned(1,8) ,
37806	 => std_logic_vector(to_unsigned(3,8) ,
37807	 => std_logic_vector(to_unsigned(4,8) ,
37808	 => std_logic_vector(to_unsigned(1,8) ,
37809	 => std_logic_vector(to_unsigned(0,8) ,
37810	 => std_logic_vector(to_unsigned(1,8) ,
37811	 => std_logic_vector(to_unsigned(3,8) ,
37812	 => std_logic_vector(to_unsigned(3,8) ,
37813	 => std_logic_vector(to_unsigned(3,8) ,
37814	 => std_logic_vector(to_unsigned(4,8) ,
37815	 => std_logic_vector(to_unsigned(3,8) ,
37816	 => std_logic_vector(to_unsigned(4,8) ,
37817	 => std_logic_vector(to_unsigned(6,8) ,
37818	 => std_logic_vector(to_unsigned(8,8) ,
37819	 => std_logic_vector(to_unsigned(7,8) ,
37820	 => std_logic_vector(to_unsigned(11,8) ,
37821	 => std_logic_vector(to_unsigned(14,8) ,
37822	 => std_logic_vector(to_unsigned(7,8) ,
37823	 => std_logic_vector(to_unsigned(5,8) ,
37824	 => std_logic_vector(to_unsigned(5,8) ,
37825	 => std_logic_vector(to_unsigned(5,8) ,
37826	 => std_logic_vector(to_unsigned(1,8) ,
37827	 => std_logic_vector(to_unsigned(1,8) ,
37828	 => std_logic_vector(to_unsigned(3,8) ,
37829	 => std_logic_vector(to_unsigned(6,8) ,
37830	 => std_logic_vector(to_unsigned(1,8) ,
37831	 => std_logic_vector(to_unsigned(0,8) ,
37832	 => std_logic_vector(to_unsigned(0,8) ,
37833	 => std_logic_vector(to_unsigned(0,8) ,
37834	 => std_logic_vector(to_unsigned(0,8) ,
37835	 => std_logic_vector(to_unsigned(0,8) ,
37836	 => std_logic_vector(to_unsigned(1,8) ,
37837	 => std_logic_vector(to_unsigned(9,8) ,
37838	 => std_logic_vector(to_unsigned(7,8) ,
37839	 => std_logic_vector(to_unsigned(3,8) ,
37840	 => std_logic_vector(to_unsigned(4,8) ,
37841	 => std_logic_vector(to_unsigned(6,8) ,
37842	 => std_logic_vector(to_unsigned(6,8) ,
37843	 => std_logic_vector(to_unsigned(3,8) ,
37844	 => std_logic_vector(to_unsigned(5,8) ,
37845	 => std_logic_vector(to_unsigned(10,8) ,
37846	 => std_logic_vector(to_unsigned(2,8) ,
37847	 => std_logic_vector(to_unsigned(0,8) ,
37848	 => std_logic_vector(to_unsigned(0,8) ,
37849	 => std_logic_vector(to_unsigned(0,8) ,
37850	 => std_logic_vector(to_unsigned(0,8) ,
37851	 => std_logic_vector(to_unsigned(0,8) ,
37852	 => std_logic_vector(to_unsigned(4,8) ,
37853	 => std_logic_vector(to_unsigned(13,8) ,
37854	 => std_logic_vector(to_unsigned(6,8) ,
37855	 => std_logic_vector(to_unsigned(6,8) ,
37856	 => std_logic_vector(to_unsigned(7,8) ,
37857	 => std_logic_vector(to_unsigned(6,8) ,
37858	 => std_logic_vector(to_unsigned(6,8) ,
37859	 => std_logic_vector(to_unsigned(3,8) ,
37860	 => std_logic_vector(to_unsigned(2,8) ,
37861	 => std_logic_vector(to_unsigned(2,8) ,
37862	 => std_logic_vector(to_unsigned(2,8) ,
37863	 => std_logic_vector(to_unsigned(9,8) ,
37864	 => std_logic_vector(to_unsigned(6,8) ,
37865	 => std_logic_vector(to_unsigned(5,8) ,
37866	 => std_logic_vector(to_unsigned(5,8) ,
37867	 => std_logic_vector(to_unsigned(3,8) ,
37868	 => std_logic_vector(to_unsigned(2,8) ,
37869	 => std_logic_vector(to_unsigned(2,8) ,
37870	 => std_logic_vector(to_unsigned(1,8) ,
37871	 => std_logic_vector(to_unsigned(0,8) ,
37872	 => std_logic_vector(to_unsigned(11,8) ,
37873	 => std_logic_vector(to_unsigned(147,8) ,
37874	 => std_logic_vector(to_unsigned(161,8) ,
37875	 => std_logic_vector(to_unsigned(146,8) ,
37876	 => std_logic_vector(to_unsigned(163,8) ,
37877	 => std_logic_vector(to_unsigned(66,8) ,
37878	 => std_logic_vector(to_unsigned(1,8) ,
37879	 => std_logic_vector(to_unsigned(1,8) ,
37880	 => std_logic_vector(to_unsigned(1,8) ,
37881	 => std_logic_vector(to_unsigned(0,8) ,
37882	 => std_logic_vector(to_unsigned(1,8) ,
37883	 => std_logic_vector(to_unsigned(2,8) ,
37884	 => std_logic_vector(to_unsigned(6,8) ,
37885	 => std_logic_vector(to_unsigned(7,8) ,
37886	 => std_logic_vector(to_unsigned(3,8) ,
37887	 => std_logic_vector(to_unsigned(3,8) ,
37888	 => std_logic_vector(to_unsigned(4,8) ,
37889	 => std_logic_vector(to_unsigned(2,8) ,
37890	 => std_logic_vector(to_unsigned(0,8) ,
37891	 => std_logic_vector(to_unsigned(3,8) ,
37892	 => std_logic_vector(to_unsigned(7,8) ,
37893	 => std_logic_vector(to_unsigned(4,8) ,
37894	 => std_logic_vector(to_unsigned(4,8) ,
37895	 => std_logic_vector(to_unsigned(6,8) ,
37896	 => std_logic_vector(to_unsigned(5,8) ,
37897	 => std_logic_vector(to_unsigned(4,8) ,
37898	 => std_logic_vector(to_unsigned(5,8) ,
37899	 => std_logic_vector(to_unsigned(3,8) ,
37900	 => std_logic_vector(to_unsigned(3,8) ,
37901	 => std_logic_vector(to_unsigned(4,8) ,
37902	 => std_logic_vector(to_unsigned(2,8) ,
37903	 => std_logic_vector(to_unsigned(1,8) ,
37904	 => std_logic_vector(to_unsigned(0,8) ,
37905	 => std_logic_vector(to_unsigned(1,8) ,
37906	 => std_logic_vector(to_unsigned(2,8) ,
37907	 => std_logic_vector(to_unsigned(3,8) ,
37908	 => std_logic_vector(to_unsigned(4,8) ,
37909	 => std_logic_vector(to_unsigned(3,8) ,
37910	 => std_logic_vector(to_unsigned(3,8) ,
37911	 => std_logic_vector(to_unsigned(2,8) ,
37912	 => std_logic_vector(to_unsigned(3,8) ,
37913	 => std_logic_vector(to_unsigned(9,8) ,
37914	 => std_logic_vector(to_unsigned(9,8) ,
37915	 => std_logic_vector(to_unsigned(8,8) ,
37916	 => std_logic_vector(to_unsigned(5,8) ,
37917	 => std_logic_vector(to_unsigned(1,8) ,
37918	 => std_logic_vector(to_unsigned(0,8) ,
37919	 => std_logic_vector(to_unsigned(6,8) ,
37920	 => std_logic_vector(to_unsigned(10,8) ,
37921	 => std_logic_vector(to_unsigned(6,8) ,
37922	 => std_logic_vector(to_unsigned(7,8) ,
37923	 => std_logic_vector(to_unsigned(6,8) ,
37924	 => std_logic_vector(to_unsigned(2,8) ,
37925	 => std_logic_vector(to_unsigned(2,8) ,
37926	 => std_logic_vector(to_unsigned(1,8) ,
37927	 => std_logic_vector(to_unsigned(0,8) ,
37928	 => std_logic_vector(to_unsigned(0,8) ,
37929	 => std_logic_vector(to_unsigned(0,8) ,
37930	 => std_logic_vector(to_unsigned(1,8) ,
37931	 => std_logic_vector(to_unsigned(1,8) ,
37932	 => std_logic_vector(to_unsigned(1,8) ,
37933	 => std_logic_vector(to_unsigned(2,8) ,
37934	 => std_logic_vector(to_unsigned(2,8) ,
37935	 => std_logic_vector(to_unsigned(1,8) ,
37936	 => std_logic_vector(to_unsigned(3,8) ,
37937	 => std_logic_vector(to_unsigned(7,8) ,
37938	 => std_logic_vector(to_unsigned(4,8) ,
37939	 => std_logic_vector(to_unsigned(5,8) ,
37940	 => std_logic_vector(to_unsigned(4,8) ,
37941	 => std_logic_vector(to_unsigned(0,8) ,
37942	 => std_logic_vector(to_unsigned(1,8) ,
37943	 => std_logic_vector(to_unsigned(6,8) ,
37944	 => std_logic_vector(to_unsigned(4,8) ,
37945	 => std_logic_vector(to_unsigned(4,8) ,
37946	 => std_logic_vector(to_unsigned(3,8) ,
37947	 => std_logic_vector(to_unsigned(2,8) ,
37948	 => std_logic_vector(to_unsigned(2,8) ,
37949	 => std_logic_vector(to_unsigned(2,8) ,
37950	 => std_logic_vector(to_unsigned(2,8) ,
37951	 => std_logic_vector(to_unsigned(0,8) ,
37952	 => std_logic_vector(to_unsigned(0,8) ,
37953	 => std_logic_vector(to_unsigned(0,8) ,
37954	 => std_logic_vector(to_unsigned(0,8) ,
37955	 => std_logic_vector(to_unsigned(0,8) ,
37956	 => std_logic_vector(to_unsigned(1,8) ,
37957	 => std_logic_vector(to_unsigned(1,8) ,
37958	 => std_logic_vector(to_unsigned(1,8) ,
37959	 => std_logic_vector(to_unsigned(1,8) ,
37960	 => std_logic_vector(to_unsigned(1,8) ,
37961	 => std_logic_vector(to_unsigned(2,8) ,
37962	 => std_logic_vector(to_unsigned(1,8) ,
37963	 => std_logic_vector(to_unsigned(1,8) ,
37964	 => std_logic_vector(to_unsigned(1,8) ,
37965	 => std_logic_vector(to_unsigned(1,8) ,
37966	 => std_logic_vector(to_unsigned(1,8) ,
37967	 => std_logic_vector(to_unsigned(2,8) ,
37968	 => std_logic_vector(to_unsigned(3,8) ,
37969	 => std_logic_vector(to_unsigned(3,8) ,
37970	 => std_logic_vector(to_unsigned(3,8) ,
37971	 => std_logic_vector(to_unsigned(6,8) ,
37972	 => std_logic_vector(to_unsigned(1,8) ,
37973	 => std_logic_vector(to_unsigned(5,8) ,
37974	 => std_logic_vector(to_unsigned(17,8) ,
37975	 => std_logic_vector(to_unsigned(28,8) ,
37976	 => std_logic_vector(to_unsigned(47,8) ,
37977	 => std_logic_vector(to_unsigned(39,8) ,
37978	 => std_logic_vector(to_unsigned(29,8) ,
37979	 => std_logic_vector(to_unsigned(22,8) ,
37980	 => std_logic_vector(to_unsigned(24,8) ,
37981	 => std_logic_vector(to_unsigned(6,8) ,
37982	 => std_logic_vector(to_unsigned(0,8) ,
37983	 => std_logic_vector(to_unsigned(1,8) ,
37984	 => std_logic_vector(to_unsigned(0,8) ,
37985	 => std_logic_vector(to_unsigned(0,8) ,
37986	 => std_logic_vector(to_unsigned(1,8) ,
37987	 => std_logic_vector(to_unsigned(1,8) ,
37988	 => std_logic_vector(to_unsigned(1,8) ,
37989	 => std_logic_vector(to_unsigned(5,8) ,
37990	 => std_logic_vector(to_unsigned(46,8) ,
37991	 => std_logic_vector(to_unsigned(90,8) ,
37992	 => std_logic_vector(to_unsigned(86,8) ,
37993	 => std_logic_vector(to_unsigned(48,8) ,
37994	 => std_logic_vector(to_unsigned(33,8) ,
37995	 => std_logic_vector(to_unsigned(17,8) ,
37996	 => std_logic_vector(to_unsigned(3,8) ,
37997	 => std_logic_vector(to_unsigned(2,8) ,
37998	 => std_logic_vector(to_unsigned(2,8) ,
37999	 => std_logic_vector(to_unsigned(2,8) ,
38000	 => std_logic_vector(to_unsigned(3,8) ,
38001	 => std_logic_vector(to_unsigned(1,8) ,
38002	 => std_logic_vector(to_unsigned(2,8) ,
38003	 => std_logic_vector(to_unsigned(2,8) ,
38004	 => std_logic_vector(to_unsigned(4,8) ,
38005	 => std_logic_vector(to_unsigned(31,8) ,
38006	 => std_logic_vector(to_unsigned(35,8) ,
38007	 => std_logic_vector(to_unsigned(4,8) ,
38008	 => std_logic_vector(to_unsigned(0,8) ,
38009	 => std_logic_vector(to_unsigned(1,8) ,
38010	 => std_logic_vector(to_unsigned(2,8) ,
38011	 => std_logic_vector(to_unsigned(4,8) ,
38012	 => std_logic_vector(to_unsigned(4,8) ,
38013	 => std_logic_vector(to_unsigned(4,8) ,
38014	 => std_logic_vector(to_unsigned(4,8) ,
38015	 => std_logic_vector(to_unsigned(5,8) ,
38016	 => std_logic_vector(to_unsigned(4,8) ,
38017	 => std_logic_vector(to_unsigned(2,8) ,
38018	 => std_logic_vector(to_unsigned(3,8) ,
38019	 => std_logic_vector(to_unsigned(3,8) ,
38020	 => std_logic_vector(to_unsigned(3,8) ,
38021	 => std_logic_vector(to_unsigned(6,8) ,
38022	 => std_logic_vector(to_unsigned(6,8) ,
38023	 => std_logic_vector(to_unsigned(4,8) ,
38024	 => std_logic_vector(to_unsigned(14,8) ,
38025	 => std_logic_vector(to_unsigned(37,8) ,
38026	 => std_logic_vector(to_unsigned(23,8) ,
38027	 => std_logic_vector(to_unsigned(11,8) ,
38028	 => std_logic_vector(to_unsigned(10,8) ,
38029	 => std_logic_vector(to_unsigned(29,8) ,
38030	 => std_logic_vector(to_unsigned(70,8) ,
38031	 => std_logic_vector(to_unsigned(62,8) ,
38032	 => std_logic_vector(to_unsigned(56,8) ,
38033	 => std_logic_vector(to_unsigned(23,8) ,
38034	 => std_logic_vector(to_unsigned(25,8) ,
38035	 => std_logic_vector(to_unsigned(33,8) ,
38036	 => std_logic_vector(to_unsigned(21,8) ,
38037	 => std_logic_vector(to_unsigned(13,8) ,
38038	 => std_logic_vector(to_unsigned(12,8) ,
38039	 => std_logic_vector(to_unsigned(18,8) ,
38040	 => std_logic_vector(to_unsigned(12,8) ,
38041	 => std_logic_vector(to_unsigned(3,8) ,
38042	 => std_logic_vector(to_unsigned(1,8) ,
38043	 => std_logic_vector(to_unsigned(2,8) ,
38044	 => std_logic_vector(to_unsigned(4,8) ,
38045	 => std_logic_vector(to_unsigned(6,8) ,
38046	 => std_logic_vector(to_unsigned(8,8) ,
38047	 => std_logic_vector(to_unsigned(16,8) ,
38048	 => std_logic_vector(to_unsigned(35,8) ,
38049	 => std_logic_vector(to_unsigned(51,8) ,
38050	 => std_logic_vector(to_unsigned(22,8) ,
38051	 => std_logic_vector(to_unsigned(10,8) ,
38052	 => std_logic_vector(to_unsigned(4,8) ,
38053	 => std_logic_vector(to_unsigned(2,8) ,
38054	 => std_logic_vector(to_unsigned(6,8) ,
38055	 => std_logic_vector(to_unsigned(10,8) ,
38056	 => std_logic_vector(to_unsigned(6,8) ,
38057	 => std_logic_vector(to_unsigned(2,8) ,
38058	 => std_logic_vector(to_unsigned(2,8) ,
38059	 => std_logic_vector(to_unsigned(2,8) ,
38060	 => std_logic_vector(to_unsigned(2,8) ,
38061	 => std_logic_vector(to_unsigned(2,8) ,
38062	 => std_logic_vector(to_unsigned(1,8) ,
38063	 => std_logic_vector(to_unsigned(1,8) ,
38064	 => std_logic_vector(to_unsigned(0,8) ,
38065	 => std_logic_vector(to_unsigned(0,8) ,
38066	 => std_logic_vector(to_unsigned(0,8) ,
38067	 => std_logic_vector(to_unsigned(0,8) ,
38068	 => std_logic_vector(to_unsigned(0,8) ,
38069	 => std_logic_vector(to_unsigned(1,8) ,
38070	 => std_logic_vector(to_unsigned(2,8) ,
38071	 => std_logic_vector(to_unsigned(5,8) ,
38072	 => std_logic_vector(to_unsigned(8,8) ,
38073	 => std_logic_vector(to_unsigned(11,8) ,
38074	 => std_logic_vector(to_unsigned(17,8) ,
38075	 => std_logic_vector(to_unsigned(22,8) ,
38076	 => std_logic_vector(to_unsigned(30,8) ,
38077	 => std_logic_vector(to_unsigned(35,8) ,
38078	 => std_logic_vector(to_unsigned(45,8) ,
38079	 => std_logic_vector(to_unsigned(54,8) ,
38080	 => std_logic_vector(to_unsigned(71,8) ,
38081	 => std_logic_vector(to_unsigned(138,8) ,
38082	 => std_logic_vector(to_unsigned(142,8) ,
38083	 => std_logic_vector(to_unsigned(142,8) ,
38084	 => std_logic_vector(to_unsigned(139,8) ,
38085	 => std_logic_vector(to_unsigned(136,8) ,
38086	 => std_logic_vector(to_unsigned(138,8) ,
38087	 => std_logic_vector(to_unsigned(130,8) ,
38088	 => std_logic_vector(to_unsigned(133,8) ,
38089	 => std_logic_vector(to_unsigned(127,8) ,
38090	 => std_logic_vector(to_unsigned(127,8) ,
38091	 => std_logic_vector(to_unsigned(131,8) ,
38092	 => std_logic_vector(to_unsigned(136,8) ,
38093	 => std_logic_vector(to_unsigned(136,8) ,
38094	 => std_logic_vector(to_unsigned(152,8) ,
38095	 => std_logic_vector(to_unsigned(41,8) ,
38096	 => std_logic_vector(to_unsigned(1,8) ,
38097	 => std_logic_vector(to_unsigned(9,8) ,
38098	 => std_logic_vector(to_unsigned(13,8) ,
38099	 => std_logic_vector(to_unsigned(1,8) ,
38100	 => std_logic_vector(to_unsigned(25,8) ,
38101	 => std_logic_vector(to_unsigned(164,8) ,
38102	 => std_logic_vector(to_unsigned(152,8) ,
38103	 => std_logic_vector(to_unsigned(146,8) ,
38104	 => std_logic_vector(to_unsigned(144,8) ,
38105	 => std_logic_vector(to_unsigned(144,8) ,
38106	 => std_logic_vector(to_unsigned(152,8) ,
38107	 => std_logic_vector(to_unsigned(166,8) ,
38108	 => std_logic_vector(to_unsigned(157,8) ,
38109	 => std_logic_vector(to_unsigned(171,8) ,
38110	 => std_logic_vector(to_unsigned(100,8) ,
38111	 => std_logic_vector(to_unsigned(8,8) ,
38112	 => std_logic_vector(to_unsigned(6,8) ,
38113	 => std_logic_vector(to_unsigned(6,8) ,
38114	 => std_logic_vector(to_unsigned(5,8) ,
38115	 => std_logic_vector(to_unsigned(3,8) ,
38116	 => std_logic_vector(to_unsigned(3,8) ,
38117	 => std_logic_vector(to_unsigned(4,8) ,
38118	 => std_logic_vector(to_unsigned(3,8) ,
38119	 => std_logic_vector(to_unsigned(4,8) ,
38120	 => std_logic_vector(to_unsigned(7,8) ,
38121	 => std_logic_vector(to_unsigned(9,8) ,
38122	 => std_logic_vector(to_unsigned(9,8) ,
38123	 => std_logic_vector(to_unsigned(2,8) ,
38124	 => std_logic_vector(to_unsigned(1,8) ,
38125	 => std_logic_vector(to_unsigned(5,8) ,
38126	 => std_logic_vector(to_unsigned(16,8) ,
38127	 => std_logic_vector(to_unsigned(7,8) ,
38128	 => std_logic_vector(to_unsigned(3,8) ,
38129	 => std_logic_vector(to_unsigned(3,8) ,
38130	 => std_logic_vector(to_unsigned(3,8) ,
38131	 => std_logic_vector(to_unsigned(2,8) ,
38132	 => std_logic_vector(to_unsigned(1,8) ,
38133	 => std_logic_vector(to_unsigned(2,8) ,
38134	 => std_logic_vector(to_unsigned(2,8) ,
38135	 => std_logic_vector(to_unsigned(2,8) ,
38136	 => std_logic_vector(to_unsigned(2,8) ,
38137	 => std_logic_vector(to_unsigned(1,8) ,
38138	 => std_logic_vector(to_unsigned(3,8) ,
38139	 => std_logic_vector(to_unsigned(7,8) ,
38140	 => std_logic_vector(to_unsigned(13,8) ,
38141	 => std_logic_vector(to_unsigned(10,8) ,
38142	 => std_logic_vector(to_unsigned(2,8) ,
38143	 => std_logic_vector(to_unsigned(6,8) ,
38144	 => std_logic_vector(to_unsigned(8,8) ,
38145	 => std_logic_vector(to_unsigned(1,8) ,
38146	 => std_logic_vector(to_unsigned(0,8) ,
38147	 => std_logic_vector(to_unsigned(1,8) ,
38148	 => std_logic_vector(to_unsigned(3,8) ,
38149	 => std_logic_vector(to_unsigned(4,8) ,
38150	 => std_logic_vector(to_unsigned(6,8) ,
38151	 => std_logic_vector(to_unsigned(3,8) ,
38152	 => std_logic_vector(to_unsigned(0,8) ,
38153	 => std_logic_vector(to_unsigned(0,8) ,
38154	 => std_logic_vector(to_unsigned(0,8) ,
38155	 => std_logic_vector(to_unsigned(0,8) ,
38156	 => std_logic_vector(to_unsigned(1,8) ,
38157	 => std_logic_vector(to_unsigned(9,8) ,
38158	 => std_logic_vector(to_unsigned(7,8) ,
38159	 => std_logic_vector(to_unsigned(2,8) ,
38160	 => std_logic_vector(to_unsigned(4,8) ,
38161	 => std_logic_vector(to_unsigned(6,8) ,
38162	 => std_logic_vector(to_unsigned(6,8) ,
38163	 => std_logic_vector(to_unsigned(4,8) ,
38164	 => std_logic_vector(to_unsigned(8,8) ,
38165	 => std_logic_vector(to_unsigned(8,8) ,
38166	 => std_logic_vector(to_unsigned(1,8) ,
38167	 => std_logic_vector(to_unsigned(0,8) ,
38168	 => std_logic_vector(to_unsigned(0,8) ,
38169	 => std_logic_vector(to_unsigned(0,8) ,
38170	 => std_logic_vector(to_unsigned(0,8) ,
38171	 => std_logic_vector(to_unsigned(0,8) ,
38172	 => std_logic_vector(to_unsigned(3,8) ,
38173	 => std_logic_vector(to_unsigned(9,8) ,
38174	 => std_logic_vector(to_unsigned(6,8) ,
38175	 => std_logic_vector(to_unsigned(5,8) ,
38176	 => std_logic_vector(to_unsigned(5,8) ,
38177	 => std_logic_vector(to_unsigned(5,8) ,
38178	 => std_logic_vector(to_unsigned(7,8) ,
38179	 => std_logic_vector(to_unsigned(2,8) ,
38180	 => std_logic_vector(to_unsigned(1,8) ,
38181	 => std_logic_vector(to_unsigned(1,8) ,
38182	 => std_logic_vector(to_unsigned(1,8) ,
38183	 => std_logic_vector(to_unsigned(7,8) ,
38184	 => std_logic_vector(to_unsigned(7,8) ,
38185	 => std_logic_vector(to_unsigned(6,8) ,
38186	 => std_logic_vector(to_unsigned(5,8) ,
38187	 => std_logic_vector(to_unsigned(3,8) ,
38188	 => std_logic_vector(to_unsigned(2,8) ,
38189	 => std_logic_vector(to_unsigned(1,8) ,
38190	 => std_logic_vector(to_unsigned(1,8) ,
38191	 => std_logic_vector(to_unsigned(1,8) ,
38192	 => std_logic_vector(to_unsigned(0,8) ,
38193	 => std_logic_vector(to_unsigned(65,8) ,
38194	 => std_logic_vector(to_unsigned(186,8) ,
38195	 => std_logic_vector(to_unsigned(152,8) ,
38196	 => std_logic_vector(to_unsigned(157,8) ,
38197	 => std_logic_vector(to_unsigned(136,8) ,
38198	 => std_logic_vector(to_unsigned(14,8) ,
38199	 => std_logic_vector(to_unsigned(0,8) ,
38200	 => std_logic_vector(to_unsigned(1,8) ,
38201	 => std_logic_vector(to_unsigned(1,8) ,
38202	 => std_logic_vector(to_unsigned(1,8) ,
38203	 => std_logic_vector(to_unsigned(1,8) ,
38204	 => std_logic_vector(to_unsigned(8,8) ,
38205	 => std_logic_vector(to_unsigned(8,8) ,
38206	 => std_logic_vector(to_unsigned(4,8) ,
38207	 => std_logic_vector(to_unsigned(4,8) ,
38208	 => std_logic_vector(to_unsigned(4,8) ,
38209	 => std_logic_vector(to_unsigned(2,8) ,
38210	 => std_logic_vector(to_unsigned(0,8) ,
38211	 => std_logic_vector(to_unsigned(3,8) ,
38212	 => std_logic_vector(to_unsigned(8,8) ,
38213	 => std_logic_vector(to_unsigned(5,8) ,
38214	 => std_logic_vector(to_unsigned(3,8) ,
38215	 => std_logic_vector(to_unsigned(4,8) ,
38216	 => std_logic_vector(to_unsigned(7,8) ,
38217	 => std_logic_vector(to_unsigned(5,8) ,
38218	 => std_logic_vector(to_unsigned(4,8) ,
38219	 => std_logic_vector(to_unsigned(2,8) ,
38220	 => std_logic_vector(to_unsigned(3,8) ,
38221	 => std_logic_vector(to_unsigned(3,8) ,
38222	 => std_logic_vector(to_unsigned(3,8) ,
38223	 => std_logic_vector(to_unsigned(2,8) ,
38224	 => std_logic_vector(to_unsigned(0,8) ,
38225	 => std_logic_vector(to_unsigned(1,8) ,
38226	 => std_logic_vector(to_unsigned(1,8) ,
38227	 => std_logic_vector(to_unsigned(2,8) ,
38228	 => std_logic_vector(to_unsigned(2,8) ,
38229	 => std_logic_vector(to_unsigned(2,8) ,
38230	 => std_logic_vector(to_unsigned(2,8) ,
38231	 => std_logic_vector(to_unsigned(2,8) ,
38232	 => std_logic_vector(to_unsigned(4,8) ,
38233	 => std_logic_vector(to_unsigned(7,8) ,
38234	 => std_logic_vector(to_unsigned(7,8) ,
38235	 => std_logic_vector(to_unsigned(6,8) ,
38236	 => std_logic_vector(to_unsigned(4,8) ,
38237	 => std_logic_vector(to_unsigned(1,8) ,
38238	 => std_logic_vector(to_unsigned(0,8) ,
38239	 => std_logic_vector(to_unsigned(6,8) ,
38240	 => std_logic_vector(to_unsigned(7,8) ,
38241	 => std_logic_vector(to_unsigned(6,8) ,
38242	 => std_logic_vector(to_unsigned(5,8) ,
38243	 => std_logic_vector(to_unsigned(6,8) ,
38244	 => std_logic_vector(to_unsigned(4,8) ,
38245	 => std_logic_vector(to_unsigned(2,8) ,
38246	 => std_logic_vector(to_unsigned(2,8) ,
38247	 => std_logic_vector(to_unsigned(1,8) ,
38248	 => std_logic_vector(to_unsigned(1,8) ,
38249	 => std_logic_vector(to_unsigned(1,8) ,
38250	 => std_logic_vector(to_unsigned(1,8) ,
38251	 => std_logic_vector(to_unsigned(1,8) ,
38252	 => std_logic_vector(to_unsigned(1,8) ,
38253	 => std_logic_vector(to_unsigned(1,8) ,
38254	 => std_logic_vector(to_unsigned(2,8) ,
38255	 => std_logic_vector(to_unsigned(1,8) ,
38256	 => std_logic_vector(to_unsigned(3,8) ,
38257	 => std_logic_vector(to_unsigned(6,8) ,
38258	 => std_logic_vector(to_unsigned(6,8) ,
38259	 => std_logic_vector(to_unsigned(4,8) ,
38260	 => std_logic_vector(to_unsigned(3,8) ,
38261	 => std_logic_vector(to_unsigned(1,8) ,
38262	 => std_logic_vector(to_unsigned(1,8) ,
38263	 => std_logic_vector(to_unsigned(6,8) ,
38264	 => std_logic_vector(to_unsigned(4,8) ,
38265	 => std_logic_vector(to_unsigned(3,8) ,
38266	 => std_logic_vector(to_unsigned(3,8) ,
38267	 => std_logic_vector(to_unsigned(4,8) ,
38268	 => std_logic_vector(to_unsigned(2,8) ,
38269	 => std_logic_vector(to_unsigned(2,8) ,
38270	 => std_logic_vector(to_unsigned(2,8) ,
38271	 => std_logic_vector(to_unsigned(0,8) ,
38272	 => std_logic_vector(to_unsigned(0,8) ,
38273	 => std_logic_vector(to_unsigned(0,8) ,
38274	 => std_logic_vector(to_unsigned(0,8) ,
38275	 => std_logic_vector(to_unsigned(0,8) ,
38276	 => std_logic_vector(to_unsigned(1,8) ,
38277	 => std_logic_vector(to_unsigned(1,8) ,
38278	 => std_logic_vector(to_unsigned(1,8) ,
38279	 => std_logic_vector(to_unsigned(1,8) ,
38280	 => std_logic_vector(to_unsigned(1,8) ,
38281	 => std_logic_vector(to_unsigned(2,8) ,
38282	 => std_logic_vector(to_unsigned(1,8) ,
38283	 => std_logic_vector(to_unsigned(1,8) ,
38284	 => std_logic_vector(to_unsigned(2,8) ,
38285	 => std_logic_vector(to_unsigned(1,8) ,
38286	 => std_logic_vector(to_unsigned(2,8) ,
38287	 => std_logic_vector(to_unsigned(3,8) ,
38288	 => std_logic_vector(to_unsigned(4,8) ,
38289	 => std_logic_vector(to_unsigned(3,8) ,
38290	 => std_logic_vector(to_unsigned(6,8) ,
38291	 => std_logic_vector(to_unsigned(8,8) ,
38292	 => std_logic_vector(to_unsigned(2,8) ,
38293	 => std_logic_vector(to_unsigned(3,8) ,
38294	 => std_logic_vector(to_unsigned(27,8) ,
38295	 => std_logic_vector(to_unsigned(51,8) ,
38296	 => std_logic_vector(to_unsigned(58,8) ,
38297	 => std_logic_vector(to_unsigned(44,8) ,
38298	 => std_logic_vector(to_unsigned(39,8) ,
38299	 => std_logic_vector(to_unsigned(30,8) ,
38300	 => std_logic_vector(to_unsigned(27,8) ,
38301	 => std_logic_vector(to_unsigned(5,8) ,
38302	 => std_logic_vector(to_unsigned(0,8) ,
38303	 => std_logic_vector(to_unsigned(1,8) ,
38304	 => std_logic_vector(to_unsigned(0,8) ,
38305	 => std_logic_vector(to_unsigned(0,8) ,
38306	 => std_logic_vector(to_unsigned(1,8) ,
38307	 => std_logic_vector(to_unsigned(2,8) ,
38308	 => std_logic_vector(to_unsigned(2,8) ,
38309	 => std_logic_vector(to_unsigned(4,8) ,
38310	 => std_logic_vector(to_unsigned(48,8) ,
38311	 => std_logic_vector(to_unsigned(111,8) ,
38312	 => std_logic_vector(to_unsigned(127,8) ,
38313	 => std_logic_vector(to_unsigned(74,8) ,
38314	 => std_logic_vector(to_unsigned(37,8) ,
38315	 => std_logic_vector(to_unsigned(25,8) ,
38316	 => std_logic_vector(to_unsigned(5,8) ,
38317	 => std_logic_vector(to_unsigned(1,8) ,
38318	 => std_logic_vector(to_unsigned(1,8) ,
38319	 => std_logic_vector(to_unsigned(2,8) ,
38320	 => std_logic_vector(to_unsigned(5,8) ,
38321	 => std_logic_vector(to_unsigned(1,8) ,
38322	 => std_logic_vector(to_unsigned(1,8) ,
38323	 => std_logic_vector(to_unsigned(2,8) ,
38324	 => std_logic_vector(to_unsigned(1,8) ,
38325	 => std_logic_vector(to_unsigned(23,8) ,
38326	 => std_logic_vector(to_unsigned(42,8) ,
38327	 => std_logic_vector(to_unsigned(6,8) ,
38328	 => std_logic_vector(to_unsigned(0,8) ,
38329	 => std_logic_vector(to_unsigned(1,8) ,
38330	 => std_logic_vector(to_unsigned(1,8) ,
38331	 => std_logic_vector(to_unsigned(1,8) ,
38332	 => std_logic_vector(to_unsigned(1,8) ,
38333	 => std_logic_vector(to_unsigned(2,8) ,
38334	 => std_logic_vector(to_unsigned(2,8) ,
38335	 => std_logic_vector(to_unsigned(2,8) ,
38336	 => std_logic_vector(to_unsigned(3,8) ,
38337	 => std_logic_vector(to_unsigned(3,8) ,
38338	 => std_logic_vector(to_unsigned(3,8) ,
38339	 => std_logic_vector(to_unsigned(4,8) ,
38340	 => std_logic_vector(to_unsigned(3,8) ,
38341	 => std_logic_vector(to_unsigned(6,8) ,
38342	 => std_logic_vector(to_unsigned(4,8) ,
38343	 => std_logic_vector(to_unsigned(8,8) ,
38344	 => std_logic_vector(to_unsigned(14,8) ,
38345	 => std_logic_vector(to_unsigned(15,8) ,
38346	 => std_logic_vector(to_unsigned(32,8) ,
38347	 => std_logic_vector(to_unsigned(23,8) ,
38348	 => std_logic_vector(to_unsigned(5,8) ,
38349	 => std_logic_vector(to_unsigned(24,8) ,
38350	 => std_logic_vector(to_unsigned(70,8) ,
38351	 => std_logic_vector(to_unsigned(101,8) ,
38352	 => std_logic_vector(to_unsigned(152,8) ,
38353	 => std_logic_vector(to_unsigned(37,8) ,
38354	 => std_logic_vector(to_unsigned(1,8) ,
38355	 => std_logic_vector(to_unsigned(6,8) ,
38356	 => std_logic_vector(to_unsigned(18,8) ,
38357	 => std_logic_vector(to_unsigned(20,8) ,
38358	 => std_logic_vector(to_unsigned(12,8) ,
38359	 => std_logic_vector(to_unsigned(16,8) ,
38360	 => std_logic_vector(to_unsigned(18,8) ,
38361	 => std_logic_vector(to_unsigned(7,8) ,
38362	 => std_logic_vector(to_unsigned(2,8) ,
38363	 => std_logic_vector(to_unsigned(3,8) ,
38364	 => std_logic_vector(to_unsigned(9,8) ,
38365	 => std_logic_vector(to_unsigned(6,8) ,
38366	 => std_logic_vector(to_unsigned(3,8) ,
38367	 => std_logic_vector(to_unsigned(5,8) ,
38368	 => std_logic_vector(to_unsigned(15,8) ,
38369	 => std_logic_vector(to_unsigned(18,8) ,
38370	 => std_logic_vector(to_unsigned(18,8) ,
38371	 => std_logic_vector(to_unsigned(14,8) ,
38372	 => std_logic_vector(to_unsigned(15,8) ,
38373	 => std_logic_vector(to_unsigned(10,8) ,
38374	 => std_logic_vector(to_unsigned(9,8) ,
38375	 => std_logic_vector(to_unsigned(11,8) ,
38376	 => std_logic_vector(to_unsigned(7,8) ,
38377	 => std_logic_vector(to_unsigned(6,8) ,
38378	 => std_logic_vector(to_unsigned(10,8) ,
38379	 => std_logic_vector(to_unsigned(36,8) ,
38380	 => std_logic_vector(to_unsigned(78,8) ,
38381	 => std_logic_vector(to_unsigned(80,8) ,
38382	 => std_logic_vector(to_unsigned(85,8) ,
38383	 => std_logic_vector(to_unsigned(76,8) ,
38384	 => std_logic_vector(to_unsigned(60,8) ,
38385	 => std_logic_vector(to_unsigned(43,8) ,
38386	 => std_logic_vector(to_unsigned(38,8) ,
38387	 => std_logic_vector(to_unsigned(36,8) ,
38388	 => std_logic_vector(to_unsigned(29,8) ,
38389	 => std_logic_vector(to_unsigned(18,8) ,
38390	 => std_logic_vector(to_unsigned(10,8) ,
38391	 => std_logic_vector(to_unsigned(6,8) ,
38392	 => std_logic_vector(to_unsigned(4,8) ,
38393	 => std_logic_vector(to_unsigned(1,8) ,
38394	 => std_logic_vector(to_unsigned(0,8) ,
38395	 => std_logic_vector(to_unsigned(0,8) ,
38396	 => std_logic_vector(to_unsigned(0,8) ,
38397	 => std_logic_vector(to_unsigned(0,8) ,
38398	 => std_logic_vector(to_unsigned(0,8) ,
38399	 => std_logic_vector(to_unsigned(0,8) ,
38400	 => std_logic_vector(to_unsigned(0,8) ,
38401	 => std_logic_vector(to_unsigned(136,8) ,
38402	 => std_logic_vector(to_unsigned(146,8) ,
38403	 => std_logic_vector(to_unsigned(149,8) ,
38404	 => std_logic_vector(to_unsigned(144,8) ,
38405	 => std_logic_vector(to_unsigned(141,8) ,
38406	 => std_logic_vector(to_unsigned(142,8) ,
38407	 => std_logic_vector(to_unsigned(139,8) ,
38408	 => std_logic_vector(to_unsigned(138,8) ,
38409	 => std_logic_vector(to_unsigned(134,8) ,
38410	 => std_logic_vector(to_unsigned(136,8) ,
38411	 => std_logic_vector(to_unsigned(146,8) ,
38412	 => std_logic_vector(to_unsigned(147,8) ,
38413	 => std_logic_vector(to_unsigned(141,8) ,
38414	 => std_logic_vector(to_unsigned(151,8) ,
38415	 => std_logic_vector(to_unsigned(43,8) ,
38416	 => std_logic_vector(to_unsigned(4,8) ,
38417	 => std_logic_vector(to_unsigned(12,8) ,
38418	 => std_logic_vector(to_unsigned(13,8) ,
38419	 => std_logic_vector(to_unsigned(2,8) ,
38420	 => std_logic_vector(to_unsigned(5,8) ,
38421	 => std_logic_vector(to_unsigned(128,8) ,
38422	 => std_logic_vector(to_unsigned(173,8) ,
38423	 => std_logic_vector(to_unsigned(152,8) ,
38424	 => std_logic_vector(to_unsigned(159,8) ,
38425	 => std_logic_vector(to_unsigned(161,8) ,
38426	 => std_logic_vector(to_unsigned(157,8) ,
38427	 => std_logic_vector(to_unsigned(157,8) ,
38428	 => std_logic_vector(to_unsigned(147,8) ,
38429	 => std_logic_vector(to_unsigned(166,8) ,
38430	 => std_logic_vector(to_unsigned(52,8) ,
38431	 => std_logic_vector(to_unsigned(1,8) ,
38432	 => std_logic_vector(to_unsigned(3,8) ,
38433	 => std_logic_vector(to_unsigned(4,8) ,
38434	 => std_logic_vector(to_unsigned(4,8) ,
38435	 => std_logic_vector(to_unsigned(2,8) ,
38436	 => std_logic_vector(to_unsigned(2,8) ,
38437	 => std_logic_vector(to_unsigned(3,8) ,
38438	 => std_logic_vector(to_unsigned(4,8) ,
38439	 => std_logic_vector(to_unsigned(6,8) ,
38440	 => std_logic_vector(to_unsigned(8,8) ,
38441	 => std_logic_vector(to_unsigned(12,8) ,
38442	 => std_logic_vector(to_unsigned(5,8) ,
38443	 => std_logic_vector(to_unsigned(1,8) ,
38444	 => std_logic_vector(to_unsigned(1,8) ,
38445	 => std_logic_vector(to_unsigned(26,8) ,
38446	 => std_logic_vector(to_unsigned(144,8) ,
38447	 => std_logic_vector(to_unsigned(142,8) ,
38448	 => std_logic_vector(to_unsigned(114,8) ,
38449	 => std_logic_vector(to_unsigned(103,8) ,
38450	 => std_logic_vector(to_unsigned(84,8) ,
38451	 => std_logic_vector(to_unsigned(70,8) ,
38452	 => std_logic_vector(to_unsigned(54,8) ,
38453	 => std_logic_vector(to_unsigned(48,8) ,
38454	 => std_logic_vector(to_unsigned(35,8) ,
38455	 => std_logic_vector(to_unsigned(24,8) ,
38456	 => std_logic_vector(to_unsigned(15,8) ,
38457	 => std_logic_vector(to_unsigned(10,8) ,
38458	 => std_logic_vector(to_unsigned(3,8) ,
38459	 => std_logic_vector(to_unsigned(2,8) ,
38460	 => std_logic_vector(to_unsigned(7,8) ,
38461	 => std_logic_vector(to_unsigned(2,8) ,
38462	 => std_logic_vector(to_unsigned(4,8) ,
38463	 => std_logic_vector(to_unsigned(11,8) ,
38464	 => std_logic_vector(to_unsigned(2,8) ,
38465	 => std_logic_vector(to_unsigned(0,8) ,
38466	 => std_logic_vector(to_unsigned(0,8) ,
38467	 => std_logic_vector(to_unsigned(0,8) ,
38468	 => std_logic_vector(to_unsigned(1,8) ,
38469	 => std_logic_vector(to_unsigned(5,8) ,
38470	 => std_logic_vector(to_unsigned(5,8) ,
38471	 => std_logic_vector(to_unsigned(2,8) ,
38472	 => std_logic_vector(to_unsigned(1,8) ,
38473	 => std_logic_vector(to_unsigned(0,8) ,
38474	 => std_logic_vector(to_unsigned(0,8) ,
38475	 => std_logic_vector(to_unsigned(0,8) ,
38476	 => std_logic_vector(to_unsigned(1,8) ,
38477	 => std_logic_vector(to_unsigned(6,8) ,
38478	 => std_logic_vector(to_unsigned(4,8) ,
38479	 => std_logic_vector(to_unsigned(3,8) ,
38480	 => std_logic_vector(to_unsigned(4,8) ,
38481	 => std_logic_vector(to_unsigned(4,8) ,
38482	 => std_logic_vector(to_unsigned(5,8) ,
38483	 => std_logic_vector(to_unsigned(6,8) ,
38484	 => std_logic_vector(to_unsigned(10,8) ,
38485	 => std_logic_vector(to_unsigned(5,8) ,
38486	 => std_logic_vector(to_unsigned(1,8) ,
38487	 => std_logic_vector(to_unsigned(0,8) ,
38488	 => std_logic_vector(to_unsigned(0,8) ,
38489	 => std_logic_vector(to_unsigned(0,8) ,
38490	 => std_logic_vector(to_unsigned(0,8) ,
38491	 => std_logic_vector(to_unsigned(0,8) ,
38492	 => std_logic_vector(to_unsigned(2,8) ,
38493	 => std_logic_vector(to_unsigned(7,8) ,
38494	 => std_logic_vector(to_unsigned(5,8) ,
38495	 => std_logic_vector(to_unsigned(4,8) ,
38496	 => std_logic_vector(to_unsigned(5,8) ,
38497	 => std_logic_vector(to_unsigned(6,8) ,
38498	 => std_logic_vector(to_unsigned(7,8) ,
38499	 => std_logic_vector(to_unsigned(1,8) ,
38500	 => std_logic_vector(to_unsigned(0,8) ,
38501	 => std_logic_vector(to_unsigned(2,8) ,
38502	 => std_logic_vector(to_unsigned(1,8) ,
38503	 => std_logic_vector(to_unsigned(6,8) ,
38504	 => std_logic_vector(to_unsigned(11,8) ,
38505	 => std_logic_vector(to_unsigned(5,8) ,
38506	 => std_logic_vector(to_unsigned(3,8) ,
38507	 => std_logic_vector(to_unsigned(2,8) ,
38508	 => std_logic_vector(to_unsigned(1,8) ,
38509	 => std_logic_vector(to_unsigned(1,8) ,
38510	 => std_logic_vector(to_unsigned(0,8) ,
38511	 => std_logic_vector(to_unsigned(1,8) ,
38512	 => std_logic_vector(to_unsigned(0,8) ,
38513	 => std_logic_vector(to_unsigned(6,8) ,
38514	 => std_logic_vector(to_unsigned(107,8) ,
38515	 => std_logic_vector(to_unsigned(161,8) ,
38516	 => std_logic_vector(to_unsigned(149,8) ,
38517	 => std_logic_vector(to_unsigned(159,8) ,
38518	 => std_logic_vector(to_unsigned(52,8) ,
38519	 => std_logic_vector(to_unsigned(1,8) ,
38520	 => std_logic_vector(to_unsigned(0,8) ,
38521	 => std_logic_vector(to_unsigned(1,8) ,
38522	 => std_logic_vector(to_unsigned(0,8) ,
38523	 => std_logic_vector(to_unsigned(1,8) ,
38524	 => std_logic_vector(to_unsigned(9,8) ,
38525	 => std_logic_vector(to_unsigned(7,8) ,
38526	 => std_logic_vector(to_unsigned(3,8) ,
38527	 => std_logic_vector(to_unsigned(4,8) ,
38528	 => std_logic_vector(to_unsigned(4,8) ,
38529	 => std_logic_vector(to_unsigned(2,8) ,
38530	 => std_logic_vector(to_unsigned(0,8) ,
38531	 => std_logic_vector(to_unsigned(2,8) ,
38532	 => std_logic_vector(to_unsigned(7,8) ,
38533	 => std_logic_vector(to_unsigned(5,8) ,
38534	 => std_logic_vector(to_unsigned(4,8) ,
38535	 => std_logic_vector(to_unsigned(5,8) ,
38536	 => std_logic_vector(to_unsigned(8,8) ,
38537	 => std_logic_vector(to_unsigned(7,8) ,
38538	 => std_logic_vector(to_unsigned(4,8) ,
38539	 => std_logic_vector(to_unsigned(4,8) ,
38540	 => std_logic_vector(to_unsigned(3,8) ,
38541	 => std_logic_vector(to_unsigned(5,8) ,
38542	 => std_logic_vector(to_unsigned(5,8) ,
38543	 => std_logic_vector(to_unsigned(1,8) ,
38544	 => std_logic_vector(to_unsigned(0,8) ,
38545	 => std_logic_vector(to_unsigned(0,8) ,
38546	 => std_logic_vector(to_unsigned(1,8) ,
38547	 => std_logic_vector(to_unsigned(1,8) ,
38548	 => std_logic_vector(to_unsigned(2,8) ,
38549	 => std_logic_vector(to_unsigned(3,8) ,
38550	 => std_logic_vector(to_unsigned(3,8) ,
38551	 => std_logic_vector(to_unsigned(2,8) ,
38552	 => std_logic_vector(to_unsigned(4,8) ,
38553	 => std_logic_vector(to_unsigned(8,8) ,
38554	 => std_logic_vector(to_unsigned(8,8) ,
38555	 => std_logic_vector(to_unsigned(6,8) ,
38556	 => std_logic_vector(to_unsigned(3,8) ,
38557	 => std_logic_vector(to_unsigned(0,8) ,
38558	 => std_logic_vector(to_unsigned(1,8) ,
38559	 => std_logic_vector(to_unsigned(6,8) ,
38560	 => std_logic_vector(to_unsigned(8,8) ,
38561	 => std_logic_vector(to_unsigned(6,8) ,
38562	 => std_logic_vector(to_unsigned(5,8) ,
38563	 => std_logic_vector(to_unsigned(5,8) ,
38564	 => std_logic_vector(to_unsigned(4,8) ,
38565	 => std_logic_vector(to_unsigned(2,8) ,
38566	 => std_logic_vector(to_unsigned(2,8) ,
38567	 => std_logic_vector(to_unsigned(0,8) ,
38568	 => std_logic_vector(to_unsigned(1,8) ,
38569	 => std_logic_vector(to_unsigned(1,8) ,
38570	 => std_logic_vector(to_unsigned(1,8) ,
38571	 => std_logic_vector(to_unsigned(1,8) ,
38572	 => std_logic_vector(to_unsigned(1,8) ,
38573	 => std_logic_vector(to_unsigned(2,8) ,
38574	 => std_logic_vector(to_unsigned(2,8) ,
38575	 => std_logic_vector(to_unsigned(2,8) ,
38576	 => std_logic_vector(to_unsigned(4,8) ,
38577	 => std_logic_vector(to_unsigned(6,8) ,
38578	 => std_logic_vector(to_unsigned(3,8) ,
38579	 => std_logic_vector(to_unsigned(2,8) ,
38580	 => std_logic_vector(to_unsigned(3,8) ,
38581	 => std_logic_vector(to_unsigned(1,8) ,
38582	 => std_logic_vector(to_unsigned(1,8) ,
38583	 => std_logic_vector(to_unsigned(10,8) ,
38584	 => std_logic_vector(to_unsigned(6,8) ,
38585	 => std_logic_vector(to_unsigned(3,8) ,
38586	 => std_logic_vector(to_unsigned(2,8) ,
38587	 => std_logic_vector(to_unsigned(3,8) ,
38588	 => std_logic_vector(to_unsigned(2,8) ,
38589	 => std_logic_vector(to_unsigned(1,8) ,
38590	 => std_logic_vector(to_unsigned(1,8) ,
38591	 => std_logic_vector(to_unsigned(1,8) ,
38592	 => std_logic_vector(to_unsigned(0,8) ,
38593	 => std_logic_vector(to_unsigned(0,8) ,
38594	 => std_logic_vector(to_unsigned(0,8) ,
38595	 => std_logic_vector(to_unsigned(0,8) ,
38596	 => std_logic_vector(to_unsigned(1,8) ,
38597	 => std_logic_vector(to_unsigned(1,8) ,
38598	 => std_logic_vector(to_unsigned(2,8) ,
38599	 => std_logic_vector(to_unsigned(1,8) ,
38600	 => std_logic_vector(to_unsigned(1,8) ,
38601	 => std_logic_vector(to_unsigned(2,8) ,
38602	 => std_logic_vector(to_unsigned(2,8) ,
38603	 => std_logic_vector(to_unsigned(1,8) ,
38604	 => std_logic_vector(to_unsigned(2,8) ,
38605	 => std_logic_vector(to_unsigned(1,8) ,
38606	 => std_logic_vector(to_unsigned(1,8) ,
38607	 => std_logic_vector(to_unsigned(3,8) ,
38608	 => std_logic_vector(to_unsigned(3,8) ,
38609	 => std_logic_vector(to_unsigned(4,8) ,
38610	 => std_logic_vector(to_unsigned(9,8) ,
38611	 => std_logic_vector(to_unsigned(7,8) ,
38612	 => std_logic_vector(to_unsigned(2,8) ,
38613	 => std_logic_vector(to_unsigned(2,8) ,
38614	 => std_logic_vector(to_unsigned(25,8) ,
38615	 => std_logic_vector(to_unsigned(68,8) ,
38616	 => std_logic_vector(to_unsigned(82,8) ,
38617	 => std_logic_vector(to_unsigned(53,8) ,
38618	 => std_logic_vector(to_unsigned(32,8) ,
38619	 => std_logic_vector(to_unsigned(23,8) ,
38620	 => std_logic_vector(to_unsigned(28,8) ,
38621	 => std_logic_vector(to_unsigned(7,8) ,
38622	 => std_logic_vector(to_unsigned(0,8) ,
38623	 => std_logic_vector(to_unsigned(0,8) ,
38624	 => std_logic_vector(to_unsigned(0,8) ,
38625	 => std_logic_vector(to_unsigned(1,8) ,
38626	 => std_logic_vector(to_unsigned(1,8) ,
38627	 => std_logic_vector(to_unsigned(2,8) ,
38628	 => std_logic_vector(to_unsigned(1,8) ,
38629	 => std_logic_vector(to_unsigned(3,8) ,
38630	 => std_logic_vector(to_unsigned(59,8) ,
38631	 => std_logic_vector(to_unsigned(116,8) ,
38632	 => std_logic_vector(to_unsigned(133,8) ,
38633	 => std_logic_vector(to_unsigned(99,8) ,
38634	 => std_logic_vector(to_unsigned(50,8) ,
38635	 => std_logic_vector(to_unsigned(32,8) ,
38636	 => std_logic_vector(to_unsigned(7,8) ,
38637	 => std_logic_vector(to_unsigned(1,8) ,
38638	 => std_logic_vector(to_unsigned(2,8) ,
38639	 => std_logic_vector(to_unsigned(2,8) ,
38640	 => std_logic_vector(to_unsigned(6,8) ,
38641	 => std_logic_vector(to_unsigned(2,8) ,
38642	 => std_logic_vector(to_unsigned(1,8) ,
38643	 => std_logic_vector(to_unsigned(2,8) ,
38644	 => std_logic_vector(to_unsigned(1,8) ,
38645	 => std_logic_vector(to_unsigned(15,8) ,
38646	 => std_logic_vector(to_unsigned(35,8) ,
38647	 => std_logic_vector(to_unsigned(13,8) ,
38648	 => std_logic_vector(to_unsigned(0,8) ,
38649	 => std_logic_vector(to_unsigned(1,8) ,
38650	 => std_logic_vector(to_unsigned(1,8) ,
38651	 => std_logic_vector(to_unsigned(2,8) ,
38652	 => std_logic_vector(to_unsigned(2,8) ,
38653	 => std_logic_vector(to_unsigned(3,8) ,
38654	 => std_logic_vector(to_unsigned(3,8) ,
38655	 => std_logic_vector(to_unsigned(2,8) ,
38656	 => std_logic_vector(to_unsigned(2,8) ,
38657	 => std_logic_vector(to_unsigned(3,8) ,
38658	 => std_logic_vector(to_unsigned(4,8) ,
38659	 => std_logic_vector(to_unsigned(3,8) ,
38660	 => std_logic_vector(to_unsigned(5,8) ,
38661	 => std_logic_vector(to_unsigned(5,8) ,
38662	 => std_logic_vector(to_unsigned(8,8) ,
38663	 => std_logic_vector(to_unsigned(22,8) ,
38664	 => std_logic_vector(to_unsigned(21,8) ,
38665	 => std_logic_vector(to_unsigned(35,8) ,
38666	 => std_logic_vector(to_unsigned(39,8) ,
38667	 => std_logic_vector(to_unsigned(30,8) ,
38668	 => std_logic_vector(to_unsigned(6,8) ,
38669	 => std_logic_vector(to_unsigned(18,8) ,
38670	 => std_logic_vector(to_unsigned(41,8) ,
38671	 => std_logic_vector(to_unsigned(116,8) ,
38672	 => std_logic_vector(to_unsigned(186,8) ,
38673	 => std_logic_vector(to_unsigned(142,8) ,
38674	 => std_logic_vector(to_unsigned(45,8) ,
38675	 => std_logic_vector(to_unsigned(13,8) ,
38676	 => std_logic_vector(to_unsigned(7,8) ,
38677	 => std_logic_vector(to_unsigned(7,8) ,
38678	 => std_logic_vector(to_unsigned(11,8) ,
38679	 => std_logic_vector(to_unsigned(18,8) ,
38680	 => std_logic_vector(to_unsigned(17,8) ,
38681	 => std_logic_vector(to_unsigned(7,8) ,
38682	 => std_logic_vector(to_unsigned(2,8) ,
38683	 => std_logic_vector(to_unsigned(3,8) ,
38684	 => std_logic_vector(to_unsigned(14,8) ,
38685	 => std_logic_vector(to_unsigned(17,8) ,
38686	 => std_logic_vector(to_unsigned(13,8) ,
38687	 => std_logic_vector(to_unsigned(24,8) ,
38688	 => std_logic_vector(to_unsigned(27,8) ,
38689	 => std_logic_vector(to_unsigned(28,8) ,
38690	 => std_logic_vector(to_unsigned(34,8) ,
38691	 => std_logic_vector(to_unsigned(19,8) ,
38692	 => std_logic_vector(to_unsigned(18,8) ,
38693	 => std_logic_vector(to_unsigned(17,8) ,
38694	 => std_logic_vector(to_unsigned(10,8) ,
38695	 => std_logic_vector(to_unsigned(9,8) ,
38696	 => std_logic_vector(to_unsigned(7,8) ,
38697	 => std_logic_vector(to_unsigned(8,8) ,
38698	 => std_logic_vector(to_unsigned(16,8) ,
38699	 => std_logic_vector(to_unsigned(58,8) ,
38700	 => std_logic_vector(to_unsigned(156,8) ,
38701	 => std_logic_vector(to_unsigned(175,8) ,
38702	 => std_logic_vector(to_unsigned(181,8) ,
38703	 => std_logic_vector(to_unsigned(184,8) ,
38704	 => std_logic_vector(to_unsigned(154,8) ,
38705	 => std_logic_vector(to_unsigned(149,8) ,
38706	 => std_logic_vector(to_unsigned(171,8) ,
38707	 => std_logic_vector(to_unsigned(157,8) ,
38708	 => std_logic_vector(to_unsigned(156,8) ,
38709	 => std_logic_vector(to_unsigned(159,8) ,
38710	 => std_logic_vector(to_unsigned(141,8) ,
38711	 => std_logic_vector(to_unsigned(128,8) ,
38712	 => std_logic_vector(to_unsigned(125,8) ,
38713	 => std_logic_vector(to_unsigned(109,8) ,
38714	 => std_logic_vector(to_unsigned(92,8) ,
38715	 => std_logic_vector(to_unsigned(78,8) ,
38716	 => std_logic_vector(to_unsigned(64,8) ,
38717	 => std_logic_vector(to_unsigned(56,8) ,
38718	 => std_logic_vector(to_unsigned(39,8) ,
38719	 => std_logic_vector(to_unsigned(25,8) ,
38720	 => std_logic_vector(to_unsigned(21,8) ,
38721	 => std_logic_vector(to_unsigned(144,8) ,
38722	 => std_logic_vector(to_unsigned(147,8) ,
38723	 => std_logic_vector(to_unsigned(146,8) ,
38724	 => std_logic_vector(to_unsigned(139,8) ,
38725	 => std_logic_vector(to_unsigned(139,8) ,
38726	 => std_logic_vector(to_unsigned(138,8) ,
38727	 => std_logic_vector(to_unsigned(136,8) ,
38728	 => std_logic_vector(to_unsigned(134,8) ,
38729	 => std_logic_vector(to_unsigned(133,8) ,
38730	 => std_logic_vector(to_unsigned(130,8) ,
38731	 => std_logic_vector(to_unsigned(138,8) ,
38732	 => std_logic_vector(to_unsigned(144,8) ,
38733	 => std_logic_vector(to_unsigned(142,8) ,
38734	 => std_logic_vector(to_unsigned(149,8) ,
38735	 => std_logic_vector(to_unsigned(44,8) ,
38736	 => std_logic_vector(to_unsigned(16,8) ,
38737	 => std_logic_vector(to_unsigned(22,8) ,
38738	 => std_logic_vector(to_unsigned(17,8) ,
38739	 => std_logic_vector(to_unsigned(3,8) ,
38740	 => std_logic_vector(to_unsigned(2,8) ,
38741	 => std_logic_vector(to_unsigned(103,8) ,
38742	 => std_logic_vector(to_unsigned(177,8) ,
38743	 => std_logic_vector(to_unsigned(146,8) ,
38744	 => std_logic_vector(to_unsigned(152,8) ,
38745	 => std_logic_vector(to_unsigned(157,8) ,
38746	 => std_logic_vector(to_unsigned(156,8) ,
38747	 => std_logic_vector(to_unsigned(154,8) ,
38748	 => std_logic_vector(to_unsigned(149,8) ,
38749	 => std_logic_vector(to_unsigned(168,8) ,
38750	 => std_logic_vector(to_unsigned(93,8) ,
38751	 => std_logic_vector(to_unsigned(9,8) ,
38752	 => std_logic_vector(to_unsigned(2,8) ,
38753	 => std_logic_vector(to_unsigned(2,8) ,
38754	 => std_logic_vector(to_unsigned(7,8) ,
38755	 => std_logic_vector(to_unsigned(12,8) ,
38756	 => std_logic_vector(to_unsigned(8,8) ,
38757	 => std_logic_vector(to_unsigned(8,8) ,
38758	 => std_logic_vector(to_unsigned(8,8) ,
38759	 => std_logic_vector(to_unsigned(12,8) ,
38760	 => std_logic_vector(to_unsigned(13,8) ,
38761	 => std_logic_vector(to_unsigned(8,8) ,
38762	 => std_logic_vector(to_unsigned(3,8) ,
38763	 => std_logic_vector(to_unsigned(2,8) ,
38764	 => std_logic_vector(to_unsigned(5,8) ,
38765	 => std_logic_vector(to_unsigned(87,8) ,
38766	 => std_logic_vector(to_unsigned(190,8) ,
38767	 => std_logic_vector(to_unsigned(171,8) ,
38768	 => std_logic_vector(to_unsigned(179,8) ,
38769	 => std_logic_vector(to_unsigned(184,8) ,
38770	 => std_logic_vector(to_unsigned(184,8) ,
38771	 => std_logic_vector(to_unsigned(186,8) ,
38772	 => std_logic_vector(to_unsigned(179,8) ,
38773	 => std_logic_vector(to_unsigned(168,8) ,
38774	 => std_logic_vector(to_unsigned(164,8) ,
38775	 => std_logic_vector(to_unsigned(154,8) ,
38776	 => std_logic_vector(to_unsigned(141,8) ,
38777	 => std_logic_vector(to_unsigned(151,8) ,
38778	 => std_logic_vector(to_unsigned(64,8) ,
38779	 => std_logic_vector(to_unsigned(1,8) ,
38780	 => std_logic_vector(to_unsigned(1,8) ,
38781	 => std_logic_vector(to_unsigned(7,8) ,
38782	 => std_logic_vector(to_unsigned(12,8) ,
38783	 => std_logic_vector(to_unsigned(2,8) ,
38784	 => std_logic_vector(to_unsigned(1,8) ,
38785	 => std_logic_vector(to_unsigned(0,8) ,
38786	 => std_logic_vector(to_unsigned(1,8) ,
38787	 => std_logic_vector(to_unsigned(2,8) ,
38788	 => std_logic_vector(to_unsigned(2,8) ,
38789	 => std_logic_vector(to_unsigned(8,8) ,
38790	 => std_logic_vector(to_unsigned(3,8) ,
38791	 => std_logic_vector(to_unsigned(1,8) ,
38792	 => std_logic_vector(to_unsigned(1,8) ,
38793	 => std_logic_vector(to_unsigned(1,8) ,
38794	 => std_logic_vector(to_unsigned(0,8) ,
38795	 => std_logic_vector(to_unsigned(0,8) ,
38796	 => std_logic_vector(to_unsigned(2,8) ,
38797	 => std_logic_vector(to_unsigned(8,8) ,
38798	 => std_logic_vector(to_unsigned(3,8) ,
38799	 => std_logic_vector(to_unsigned(2,8) ,
38800	 => std_logic_vector(to_unsigned(4,8) ,
38801	 => std_logic_vector(to_unsigned(6,8) ,
38802	 => std_logic_vector(to_unsigned(5,8) ,
38803	 => std_logic_vector(to_unsigned(6,8) ,
38804	 => std_logic_vector(to_unsigned(6,8) ,
38805	 => std_logic_vector(to_unsigned(3,8) ,
38806	 => std_logic_vector(to_unsigned(1,8) ,
38807	 => std_logic_vector(to_unsigned(1,8) ,
38808	 => std_logic_vector(to_unsigned(0,8) ,
38809	 => std_logic_vector(to_unsigned(0,8) ,
38810	 => std_logic_vector(to_unsigned(1,8) ,
38811	 => std_logic_vector(to_unsigned(0,8) ,
38812	 => std_logic_vector(to_unsigned(2,8) ,
38813	 => std_logic_vector(to_unsigned(6,8) ,
38814	 => std_logic_vector(to_unsigned(6,8) ,
38815	 => std_logic_vector(to_unsigned(5,8) ,
38816	 => std_logic_vector(to_unsigned(6,8) ,
38817	 => std_logic_vector(to_unsigned(5,8) ,
38818	 => std_logic_vector(to_unsigned(5,8) ,
38819	 => std_logic_vector(to_unsigned(1,8) ,
38820	 => std_logic_vector(to_unsigned(1,8) ,
38821	 => std_logic_vector(to_unsigned(1,8) ,
38822	 => std_logic_vector(to_unsigned(0,8) ,
38823	 => std_logic_vector(to_unsigned(6,8) ,
38824	 => std_logic_vector(to_unsigned(10,8) ,
38825	 => std_logic_vector(to_unsigned(3,8) ,
38826	 => std_logic_vector(to_unsigned(3,8) ,
38827	 => std_logic_vector(to_unsigned(3,8) ,
38828	 => std_logic_vector(to_unsigned(3,8) ,
38829	 => std_logic_vector(to_unsigned(2,8) ,
38830	 => std_logic_vector(to_unsigned(0,8) ,
38831	 => std_logic_vector(to_unsigned(1,8) ,
38832	 => std_logic_vector(to_unsigned(1,8) ,
38833	 => std_logic_vector(to_unsigned(0,8) ,
38834	 => std_logic_vector(to_unsigned(15,8) ,
38835	 => std_logic_vector(to_unsigned(134,8) ,
38836	 => std_logic_vector(to_unsigned(139,8) ,
38837	 => std_logic_vector(to_unsigned(138,8) ,
38838	 => std_logic_vector(to_unsigned(105,8) ,
38839	 => std_logic_vector(to_unsigned(8,8) ,
38840	 => std_logic_vector(to_unsigned(0,8) ,
38841	 => std_logic_vector(to_unsigned(2,8) ,
38842	 => std_logic_vector(to_unsigned(1,8) ,
38843	 => std_logic_vector(to_unsigned(1,8) ,
38844	 => std_logic_vector(to_unsigned(8,8) ,
38845	 => std_logic_vector(to_unsigned(5,8) ,
38846	 => std_logic_vector(to_unsigned(3,8) ,
38847	 => std_logic_vector(to_unsigned(4,8) ,
38848	 => std_logic_vector(to_unsigned(5,8) ,
38849	 => std_logic_vector(to_unsigned(3,8) ,
38850	 => std_logic_vector(to_unsigned(0,8) ,
38851	 => std_logic_vector(to_unsigned(2,8) ,
38852	 => std_logic_vector(to_unsigned(8,8) ,
38853	 => std_logic_vector(to_unsigned(5,8) ,
38854	 => std_logic_vector(to_unsigned(4,8) ,
38855	 => std_logic_vector(to_unsigned(5,8) ,
38856	 => std_logic_vector(to_unsigned(8,8) ,
38857	 => std_logic_vector(to_unsigned(6,8) ,
38858	 => std_logic_vector(to_unsigned(4,8) ,
38859	 => std_logic_vector(to_unsigned(5,8) ,
38860	 => std_logic_vector(to_unsigned(5,8) ,
38861	 => std_logic_vector(to_unsigned(4,8) ,
38862	 => std_logic_vector(to_unsigned(3,8) ,
38863	 => std_logic_vector(to_unsigned(1,8) ,
38864	 => std_logic_vector(to_unsigned(0,8) ,
38865	 => std_logic_vector(to_unsigned(0,8) ,
38866	 => std_logic_vector(to_unsigned(1,8) ,
38867	 => std_logic_vector(to_unsigned(1,8) ,
38868	 => std_logic_vector(to_unsigned(2,8) ,
38869	 => std_logic_vector(to_unsigned(3,8) ,
38870	 => std_logic_vector(to_unsigned(3,8) ,
38871	 => std_logic_vector(to_unsigned(2,8) ,
38872	 => std_logic_vector(to_unsigned(3,8) ,
38873	 => std_logic_vector(to_unsigned(8,8) ,
38874	 => std_logic_vector(to_unsigned(8,8) ,
38875	 => std_logic_vector(to_unsigned(5,8) ,
38876	 => std_logic_vector(to_unsigned(3,8) ,
38877	 => std_logic_vector(to_unsigned(0,8) ,
38878	 => std_logic_vector(to_unsigned(2,8) ,
38879	 => std_logic_vector(to_unsigned(9,8) ,
38880	 => std_logic_vector(to_unsigned(11,8) ,
38881	 => std_logic_vector(to_unsigned(7,8) ,
38882	 => std_logic_vector(to_unsigned(5,8) ,
38883	 => std_logic_vector(to_unsigned(5,8) ,
38884	 => std_logic_vector(to_unsigned(6,8) ,
38885	 => std_logic_vector(to_unsigned(5,8) ,
38886	 => std_logic_vector(to_unsigned(2,8) ,
38887	 => std_logic_vector(to_unsigned(1,8) ,
38888	 => std_logic_vector(to_unsigned(1,8) ,
38889	 => std_logic_vector(to_unsigned(1,8) ,
38890	 => std_logic_vector(to_unsigned(1,8) ,
38891	 => std_logic_vector(to_unsigned(2,8) ,
38892	 => std_logic_vector(to_unsigned(2,8) ,
38893	 => std_logic_vector(to_unsigned(2,8) ,
38894	 => std_logic_vector(to_unsigned(2,8) ,
38895	 => std_logic_vector(to_unsigned(2,8) ,
38896	 => std_logic_vector(to_unsigned(4,8) ,
38897	 => std_logic_vector(to_unsigned(4,8) ,
38898	 => std_logic_vector(to_unsigned(2,8) ,
38899	 => std_logic_vector(to_unsigned(2,8) ,
38900	 => std_logic_vector(to_unsigned(4,8) ,
38901	 => std_logic_vector(to_unsigned(1,8) ,
38902	 => std_logic_vector(to_unsigned(1,8) ,
38903	 => std_logic_vector(to_unsigned(7,8) ,
38904	 => std_logic_vector(to_unsigned(6,8) ,
38905	 => std_logic_vector(to_unsigned(5,8) ,
38906	 => std_logic_vector(to_unsigned(2,8) ,
38907	 => std_logic_vector(to_unsigned(3,8) ,
38908	 => std_logic_vector(to_unsigned(3,8) ,
38909	 => std_logic_vector(to_unsigned(1,8) ,
38910	 => std_logic_vector(to_unsigned(1,8) ,
38911	 => std_logic_vector(to_unsigned(1,8) ,
38912	 => std_logic_vector(to_unsigned(0,8) ,
38913	 => std_logic_vector(to_unsigned(0,8) ,
38914	 => std_logic_vector(to_unsigned(1,8) ,
38915	 => std_logic_vector(to_unsigned(1,8) ,
38916	 => std_logic_vector(to_unsigned(1,8) ,
38917	 => std_logic_vector(to_unsigned(1,8) ,
38918	 => std_logic_vector(to_unsigned(2,8) ,
38919	 => std_logic_vector(to_unsigned(2,8) ,
38920	 => std_logic_vector(to_unsigned(2,8) ,
38921	 => std_logic_vector(to_unsigned(1,8) ,
38922	 => std_logic_vector(to_unsigned(1,8) ,
38923	 => std_logic_vector(to_unsigned(2,8) ,
38924	 => std_logic_vector(to_unsigned(1,8) ,
38925	 => std_logic_vector(to_unsigned(2,8) ,
38926	 => std_logic_vector(to_unsigned(1,8) ,
38927	 => std_logic_vector(to_unsigned(2,8) ,
38928	 => std_logic_vector(to_unsigned(3,8) ,
38929	 => std_logic_vector(to_unsigned(4,8) ,
38930	 => std_logic_vector(to_unsigned(8,8) ,
38931	 => std_logic_vector(to_unsigned(6,8) ,
38932	 => std_logic_vector(to_unsigned(2,8) ,
38933	 => std_logic_vector(to_unsigned(1,8) ,
38934	 => std_logic_vector(to_unsigned(20,8) ,
38935	 => std_logic_vector(to_unsigned(77,8) ,
38936	 => std_logic_vector(to_unsigned(93,8) ,
38937	 => std_logic_vector(to_unsigned(46,8) ,
38938	 => std_logic_vector(to_unsigned(18,8) ,
38939	 => std_logic_vector(to_unsigned(28,8) ,
38940	 => std_logic_vector(to_unsigned(29,8) ,
38941	 => std_logic_vector(to_unsigned(6,8) ,
38942	 => std_logic_vector(to_unsigned(0,8) ,
38943	 => std_logic_vector(to_unsigned(0,8) ,
38944	 => std_logic_vector(to_unsigned(1,8) ,
38945	 => std_logic_vector(to_unsigned(1,8) ,
38946	 => std_logic_vector(to_unsigned(1,8) ,
38947	 => std_logic_vector(to_unsigned(1,8) ,
38948	 => std_logic_vector(to_unsigned(1,8) ,
38949	 => std_logic_vector(to_unsigned(2,8) ,
38950	 => std_logic_vector(to_unsigned(52,8) ,
38951	 => std_logic_vector(to_unsigned(107,8) ,
38952	 => std_logic_vector(to_unsigned(128,8) ,
38953	 => std_logic_vector(to_unsigned(122,8) ,
38954	 => std_logic_vector(to_unsigned(51,8) ,
38955	 => std_logic_vector(to_unsigned(20,8) ,
38956	 => std_logic_vector(to_unsigned(12,8) ,
38957	 => std_logic_vector(to_unsigned(1,8) ,
38958	 => std_logic_vector(to_unsigned(1,8) ,
38959	 => std_logic_vector(to_unsigned(2,8) ,
38960	 => std_logic_vector(to_unsigned(4,8) ,
38961	 => std_logic_vector(to_unsigned(2,8) ,
38962	 => std_logic_vector(to_unsigned(1,8) ,
38963	 => std_logic_vector(to_unsigned(3,8) ,
38964	 => std_logic_vector(to_unsigned(3,8) ,
38965	 => std_logic_vector(to_unsigned(10,8) ,
38966	 => std_logic_vector(to_unsigned(32,8) ,
38967	 => std_logic_vector(to_unsigned(23,8) ,
38968	 => std_logic_vector(to_unsigned(1,8) ,
38969	 => std_logic_vector(to_unsigned(0,8) ,
38970	 => std_logic_vector(to_unsigned(1,8) ,
38971	 => std_logic_vector(to_unsigned(2,8) ,
38972	 => std_logic_vector(to_unsigned(4,8) ,
38973	 => std_logic_vector(to_unsigned(4,8) ,
38974	 => std_logic_vector(to_unsigned(2,8) ,
38975	 => std_logic_vector(to_unsigned(2,8) ,
38976	 => std_logic_vector(to_unsigned(2,8) ,
38977	 => std_logic_vector(to_unsigned(2,8) ,
38978	 => std_logic_vector(to_unsigned(3,8) ,
38979	 => std_logic_vector(to_unsigned(3,8) ,
38980	 => std_logic_vector(to_unsigned(6,8) ,
38981	 => std_logic_vector(to_unsigned(4,8) ,
38982	 => std_logic_vector(to_unsigned(11,8) ,
38983	 => std_logic_vector(to_unsigned(24,8) ,
38984	 => std_logic_vector(to_unsigned(20,8) ,
38985	 => std_logic_vector(to_unsigned(37,8) ,
38986	 => std_logic_vector(to_unsigned(30,8) ,
38987	 => std_logic_vector(to_unsigned(28,8) ,
38988	 => std_logic_vector(to_unsigned(18,8) ,
38989	 => std_logic_vector(to_unsigned(8,8) ,
38990	 => std_logic_vector(to_unsigned(46,8) ,
38991	 => std_logic_vector(to_unsigned(142,8) ,
38992	 => std_logic_vector(to_unsigned(138,8) ,
38993	 => std_logic_vector(to_unsigned(121,8) ,
38994	 => std_logic_vector(to_unsigned(146,8) ,
38995	 => std_logic_vector(to_unsigned(152,8) ,
38996	 => std_logic_vector(to_unsigned(74,8) ,
38997	 => std_logic_vector(to_unsigned(19,8) ,
38998	 => std_logic_vector(to_unsigned(3,8) ,
38999	 => std_logic_vector(to_unsigned(5,8) ,
39000	 => std_logic_vector(to_unsigned(3,8) ,
39001	 => std_logic_vector(to_unsigned(1,8) ,
39002	 => std_logic_vector(to_unsigned(1,8) ,
39003	 => std_logic_vector(to_unsigned(1,8) ,
39004	 => std_logic_vector(to_unsigned(1,8) ,
39005	 => std_logic_vector(to_unsigned(5,8) ,
39006	 => std_logic_vector(to_unsigned(19,8) ,
39007	 => std_logic_vector(to_unsigned(29,8) ,
39008	 => std_logic_vector(to_unsigned(20,8) ,
39009	 => std_logic_vector(to_unsigned(12,8) ,
39010	 => std_logic_vector(to_unsigned(17,8) ,
39011	 => std_logic_vector(to_unsigned(20,8) ,
39012	 => std_logic_vector(to_unsigned(18,8) ,
39013	 => std_logic_vector(to_unsigned(15,8) ,
39014	 => std_logic_vector(to_unsigned(12,8) ,
39015	 => std_logic_vector(to_unsigned(8,8) ,
39016	 => std_logic_vector(to_unsigned(3,8) ,
39017	 => std_logic_vector(to_unsigned(7,8) ,
39018	 => std_logic_vector(to_unsigned(8,8) ,
39019	 => std_logic_vector(to_unsigned(22,8) ,
39020	 => std_logic_vector(to_unsigned(76,8) ,
39021	 => std_logic_vector(to_unsigned(114,8) ,
39022	 => std_logic_vector(to_unsigned(125,8) ,
39023	 => std_logic_vector(to_unsigned(138,8) ,
39024	 => std_logic_vector(to_unsigned(108,8) ,
39025	 => std_logic_vector(to_unsigned(114,8) ,
39026	 => std_logic_vector(to_unsigned(146,8) ,
39027	 => std_logic_vector(to_unsigned(157,8) ,
39028	 => std_logic_vector(to_unsigned(161,8) ,
39029	 => std_logic_vector(to_unsigned(173,8) ,
39030	 => std_logic_vector(to_unsigned(175,8) ,
39031	 => std_logic_vector(to_unsigned(173,8) ,
39032	 => std_logic_vector(to_unsigned(171,8) ,
39033	 => std_logic_vector(to_unsigned(177,8) ,
39034	 => std_logic_vector(to_unsigned(186,8) ,
39035	 => std_logic_vector(to_unsigned(184,8) ,
39036	 => std_logic_vector(to_unsigned(184,8) ,
39037	 => std_logic_vector(to_unsigned(177,8) ,
39038	 => std_logic_vector(to_unsigned(173,8) ,
39039	 => std_logic_vector(to_unsigned(168,8) ,
39040	 => std_logic_vector(to_unsigned(163,8) ,
39041	 => std_logic_vector(to_unsigned(141,8) ,
39042	 => std_logic_vector(to_unsigned(139,8) ,
39043	 => std_logic_vector(to_unsigned(136,8) ,
39044	 => std_logic_vector(to_unsigned(138,8) ,
39045	 => std_logic_vector(to_unsigned(139,8) ,
39046	 => std_logic_vector(to_unsigned(139,8) ,
39047	 => std_logic_vector(to_unsigned(134,8) ,
39048	 => std_logic_vector(to_unsigned(131,8) ,
39049	 => std_logic_vector(to_unsigned(136,8) ,
39050	 => std_logic_vector(to_unsigned(136,8) ,
39051	 => std_logic_vector(to_unsigned(141,8) ,
39052	 => std_logic_vector(to_unsigned(144,8) ,
39053	 => std_logic_vector(to_unsigned(136,8) ,
39054	 => std_logic_vector(to_unsigned(152,8) ,
39055	 => std_logic_vector(to_unsigned(58,8) ,
39056	 => std_logic_vector(to_unsigned(22,8) ,
39057	 => std_logic_vector(to_unsigned(41,8) ,
39058	 => std_logic_vector(to_unsigned(19,8) ,
39059	 => std_logic_vector(to_unsigned(1,8) ,
39060	 => std_logic_vector(to_unsigned(5,8) ,
39061	 => std_logic_vector(to_unsigned(124,8) ,
39062	 => std_logic_vector(to_unsigned(168,8) ,
39063	 => std_logic_vector(to_unsigned(144,8) ,
39064	 => std_logic_vector(to_unsigned(144,8) ,
39065	 => std_logic_vector(to_unsigned(154,8) ,
39066	 => std_logic_vector(to_unsigned(159,8) ,
39067	 => std_logic_vector(to_unsigned(149,8) ,
39068	 => std_logic_vector(to_unsigned(154,8) ,
39069	 => std_logic_vector(to_unsigned(151,8) ,
39070	 => std_logic_vector(to_unsigned(157,8) ,
39071	 => std_logic_vector(to_unsigned(130,8) ,
39072	 => std_logic_vector(to_unsigned(60,8) ,
39073	 => std_logic_vector(to_unsigned(19,8) ,
39074	 => std_logic_vector(to_unsigned(6,8) ,
39075	 => std_logic_vector(to_unsigned(8,8) ,
39076	 => std_logic_vector(to_unsigned(11,8) ,
39077	 => std_logic_vector(to_unsigned(11,8) ,
39078	 => std_logic_vector(to_unsigned(13,8) ,
39079	 => std_logic_vector(to_unsigned(16,8) ,
39080	 => std_logic_vector(to_unsigned(6,8) ,
39081	 => std_logic_vector(to_unsigned(1,8) ,
39082	 => std_logic_vector(to_unsigned(3,8) ,
39083	 => std_logic_vector(to_unsigned(5,8) ,
39084	 => std_logic_vector(to_unsigned(37,8) ,
39085	 => std_logic_vector(to_unsigned(157,8) ,
39086	 => std_logic_vector(to_unsigned(164,8) ,
39087	 => std_logic_vector(to_unsigned(144,8) ,
39088	 => std_logic_vector(to_unsigned(156,8) ,
39089	 => std_logic_vector(to_unsigned(159,8) ,
39090	 => std_logic_vector(to_unsigned(157,8) ,
39091	 => std_logic_vector(to_unsigned(157,8) ,
39092	 => std_logic_vector(to_unsigned(156,8) ,
39093	 => std_logic_vector(to_unsigned(151,8) ,
39094	 => std_logic_vector(to_unsigned(156,8) ,
39095	 => std_logic_vector(to_unsigned(154,8) ,
39096	 => std_logic_vector(to_unsigned(156,8) ,
39097	 => std_logic_vector(to_unsigned(166,8) ,
39098	 => std_logic_vector(to_unsigned(134,8) ,
39099	 => std_logic_vector(to_unsigned(18,8) ,
39100	 => std_logic_vector(to_unsigned(4,8) ,
39101	 => std_logic_vector(to_unsigned(11,8) ,
39102	 => std_logic_vector(to_unsigned(2,8) ,
39103	 => std_logic_vector(to_unsigned(1,8) ,
39104	 => std_logic_vector(to_unsigned(2,8) ,
39105	 => std_logic_vector(to_unsigned(1,8) ,
39106	 => std_logic_vector(to_unsigned(30,8) ,
39107	 => std_logic_vector(to_unsigned(85,8) ,
39108	 => std_logic_vector(to_unsigned(8,8) ,
39109	 => std_logic_vector(to_unsigned(4,8) ,
39110	 => std_logic_vector(to_unsigned(16,8) ,
39111	 => std_logic_vector(to_unsigned(26,8) ,
39112	 => std_logic_vector(to_unsigned(5,8) ,
39113	 => std_logic_vector(to_unsigned(0,8) ,
39114	 => std_logic_vector(to_unsigned(4,8) ,
39115	 => std_logic_vector(to_unsigned(4,8) ,
39116	 => std_logic_vector(to_unsigned(5,8) ,
39117	 => std_logic_vector(to_unsigned(13,8) ,
39118	 => std_logic_vector(to_unsigned(8,8) ,
39119	 => std_logic_vector(to_unsigned(5,8) ,
39120	 => std_logic_vector(to_unsigned(5,8) ,
39121	 => std_logic_vector(to_unsigned(5,8) ,
39122	 => std_logic_vector(to_unsigned(5,8) ,
39123	 => std_logic_vector(to_unsigned(2,8) ,
39124	 => std_logic_vector(to_unsigned(1,8) ,
39125	 => std_logic_vector(to_unsigned(2,8) ,
39126	 => std_logic_vector(to_unsigned(1,8) ,
39127	 => std_logic_vector(to_unsigned(1,8) ,
39128	 => std_logic_vector(to_unsigned(0,8) ,
39129	 => std_logic_vector(to_unsigned(0,8) ,
39130	 => std_logic_vector(to_unsigned(1,8) ,
39131	 => std_logic_vector(to_unsigned(0,8) ,
39132	 => std_logic_vector(to_unsigned(2,8) ,
39133	 => std_logic_vector(to_unsigned(4,8) ,
39134	 => std_logic_vector(to_unsigned(5,8) ,
39135	 => std_logic_vector(to_unsigned(5,8) ,
39136	 => std_logic_vector(to_unsigned(6,8) ,
39137	 => std_logic_vector(to_unsigned(4,8) ,
39138	 => std_logic_vector(to_unsigned(6,8) ,
39139	 => std_logic_vector(to_unsigned(2,8) ,
39140	 => std_logic_vector(to_unsigned(1,8) ,
39141	 => std_logic_vector(to_unsigned(3,8) ,
39142	 => std_logic_vector(to_unsigned(0,8) ,
39143	 => std_logic_vector(to_unsigned(4,8) ,
39144	 => std_logic_vector(to_unsigned(11,8) ,
39145	 => std_logic_vector(to_unsigned(4,8) ,
39146	 => std_logic_vector(to_unsigned(5,8) ,
39147	 => std_logic_vector(to_unsigned(4,8) ,
39148	 => std_logic_vector(to_unsigned(1,8) ,
39149	 => std_logic_vector(to_unsigned(1,8) ,
39150	 => std_logic_vector(to_unsigned(1,8) ,
39151	 => std_logic_vector(to_unsigned(1,8) ,
39152	 => std_logic_vector(to_unsigned(1,8) ,
39153	 => std_logic_vector(to_unsigned(0,8) ,
39154	 => std_logic_vector(to_unsigned(1,8) ,
39155	 => std_logic_vector(to_unsigned(71,8) ,
39156	 => std_logic_vector(to_unsigned(151,8) ,
39157	 => std_logic_vector(to_unsigned(119,8) ,
39158	 => std_logic_vector(to_unsigned(131,8) ,
39159	 => std_logic_vector(to_unsigned(43,8) ,
39160	 => std_logic_vector(to_unsigned(1,8) ,
39161	 => std_logic_vector(to_unsigned(1,8) ,
39162	 => std_logic_vector(to_unsigned(1,8) ,
39163	 => std_logic_vector(to_unsigned(3,8) ,
39164	 => std_logic_vector(to_unsigned(7,8) ,
39165	 => std_logic_vector(to_unsigned(3,8) ,
39166	 => std_logic_vector(to_unsigned(3,8) ,
39167	 => std_logic_vector(to_unsigned(4,8) ,
39168	 => std_logic_vector(to_unsigned(4,8) ,
39169	 => std_logic_vector(to_unsigned(1,8) ,
39170	 => std_logic_vector(to_unsigned(0,8) ,
39171	 => std_logic_vector(to_unsigned(3,8) ,
39172	 => std_logic_vector(to_unsigned(8,8) ,
39173	 => std_logic_vector(to_unsigned(5,8) ,
39174	 => std_logic_vector(to_unsigned(3,8) ,
39175	 => std_logic_vector(to_unsigned(4,8) ,
39176	 => std_logic_vector(to_unsigned(5,8) ,
39177	 => std_logic_vector(to_unsigned(6,8) ,
39178	 => std_logic_vector(to_unsigned(6,8) ,
39179	 => std_logic_vector(to_unsigned(4,8) ,
39180	 => std_logic_vector(to_unsigned(5,8) ,
39181	 => std_logic_vector(to_unsigned(5,8) ,
39182	 => std_logic_vector(to_unsigned(4,8) ,
39183	 => std_logic_vector(to_unsigned(1,8) ,
39184	 => std_logic_vector(to_unsigned(0,8) ,
39185	 => std_logic_vector(to_unsigned(0,8) ,
39186	 => std_logic_vector(to_unsigned(1,8) ,
39187	 => std_logic_vector(to_unsigned(1,8) ,
39188	 => std_logic_vector(to_unsigned(1,8) ,
39189	 => std_logic_vector(to_unsigned(2,8) ,
39190	 => std_logic_vector(to_unsigned(2,8) ,
39191	 => std_logic_vector(to_unsigned(1,8) ,
39192	 => std_logic_vector(to_unsigned(4,8) ,
39193	 => std_logic_vector(to_unsigned(9,8) ,
39194	 => std_logic_vector(to_unsigned(8,8) ,
39195	 => std_logic_vector(to_unsigned(4,8) ,
39196	 => std_logic_vector(to_unsigned(2,8) ,
39197	 => std_logic_vector(to_unsigned(0,8) ,
39198	 => std_logic_vector(to_unsigned(2,8) ,
39199	 => std_logic_vector(to_unsigned(8,8) ,
39200	 => std_logic_vector(to_unsigned(8,8) ,
39201	 => std_logic_vector(to_unsigned(6,8) ,
39202	 => std_logic_vector(to_unsigned(7,8) ,
39203	 => std_logic_vector(to_unsigned(6,8) ,
39204	 => std_logic_vector(to_unsigned(6,8) ,
39205	 => std_logic_vector(to_unsigned(9,8) ,
39206	 => std_logic_vector(to_unsigned(4,8) ,
39207	 => std_logic_vector(to_unsigned(1,8) ,
39208	 => std_logic_vector(to_unsigned(1,8) ,
39209	 => std_logic_vector(to_unsigned(1,8) ,
39210	 => std_logic_vector(to_unsigned(1,8) ,
39211	 => std_logic_vector(to_unsigned(2,8) ,
39212	 => std_logic_vector(to_unsigned(1,8) ,
39213	 => std_logic_vector(to_unsigned(2,8) ,
39214	 => std_logic_vector(to_unsigned(1,8) ,
39215	 => std_logic_vector(to_unsigned(2,8) ,
39216	 => std_logic_vector(to_unsigned(5,8) ,
39217	 => std_logic_vector(to_unsigned(4,8) ,
39218	 => std_logic_vector(to_unsigned(2,8) ,
39219	 => std_logic_vector(to_unsigned(4,8) ,
39220	 => std_logic_vector(to_unsigned(5,8) ,
39221	 => std_logic_vector(to_unsigned(1,8) ,
39222	 => std_logic_vector(to_unsigned(1,8) ,
39223	 => std_logic_vector(to_unsigned(6,8) ,
39224	 => std_logic_vector(to_unsigned(5,8) ,
39225	 => std_logic_vector(to_unsigned(4,8) ,
39226	 => std_logic_vector(to_unsigned(2,8) ,
39227	 => std_logic_vector(to_unsigned(2,8) ,
39228	 => std_logic_vector(to_unsigned(3,8) ,
39229	 => std_logic_vector(to_unsigned(2,8) ,
39230	 => std_logic_vector(to_unsigned(1,8) ,
39231	 => std_logic_vector(to_unsigned(1,8) ,
39232	 => std_logic_vector(to_unsigned(0,8) ,
39233	 => std_logic_vector(to_unsigned(1,8) ,
39234	 => std_logic_vector(to_unsigned(0,8) ,
39235	 => std_logic_vector(to_unsigned(1,8) ,
39236	 => std_logic_vector(to_unsigned(1,8) ,
39237	 => std_logic_vector(to_unsigned(1,8) ,
39238	 => std_logic_vector(to_unsigned(1,8) ,
39239	 => std_logic_vector(to_unsigned(2,8) ,
39240	 => std_logic_vector(to_unsigned(2,8) ,
39241	 => std_logic_vector(to_unsigned(2,8) ,
39242	 => std_logic_vector(to_unsigned(2,8) ,
39243	 => std_logic_vector(to_unsigned(2,8) ,
39244	 => std_logic_vector(to_unsigned(2,8) ,
39245	 => std_logic_vector(to_unsigned(1,8) ,
39246	 => std_logic_vector(to_unsigned(2,8) ,
39247	 => std_logic_vector(to_unsigned(4,8) ,
39248	 => std_logic_vector(to_unsigned(4,8) ,
39249	 => std_logic_vector(to_unsigned(6,8) ,
39250	 => std_logic_vector(to_unsigned(8,8) ,
39251	 => std_logic_vector(to_unsigned(6,8) ,
39252	 => std_logic_vector(to_unsigned(4,8) ,
39253	 => std_logic_vector(to_unsigned(1,8) ,
39254	 => std_logic_vector(to_unsigned(25,8) ,
39255	 => std_logic_vector(to_unsigned(105,8) ,
39256	 => std_logic_vector(to_unsigned(93,8) ,
39257	 => std_logic_vector(to_unsigned(45,8) ,
39258	 => std_logic_vector(to_unsigned(30,8) ,
39259	 => std_logic_vector(to_unsigned(37,8) ,
39260	 => std_logic_vector(to_unsigned(19,8) ,
39261	 => std_logic_vector(to_unsigned(4,8) ,
39262	 => std_logic_vector(to_unsigned(0,8) ,
39263	 => std_logic_vector(to_unsigned(0,8) ,
39264	 => std_logic_vector(to_unsigned(0,8) ,
39265	 => std_logic_vector(to_unsigned(1,8) ,
39266	 => std_logic_vector(to_unsigned(1,8) ,
39267	 => std_logic_vector(to_unsigned(2,8) ,
39268	 => std_logic_vector(to_unsigned(1,8) ,
39269	 => std_logic_vector(to_unsigned(3,8) ,
39270	 => std_logic_vector(to_unsigned(66,8) ,
39271	 => std_logic_vector(to_unsigned(109,8) ,
39272	 => std_logic_vector(to_unsigned(124,8) ,
39273	 => std_logic_vector(to_unsigned(133,8) ,
39274	 => std_logic_vector(to_unsigned(54,8) ,
39275	 => std_logic_vector(to_unsigned(15,8) ,
39276	 => std_logic_vector(to_unsigned(11,8) ,
39277	 => std_logic_vector(to_unsigned(2,8) ,
39278	 => std_logic_vector(to_unsigned(1,8) ,
39279	 => std_logic_vector(to_unsigned(2,8) ,
39280	 => std_logic_vector(to_unsigned(5,8) ,
39281	 => std_logic_vector(to_unsigned(3,8) ,
39282	 => std_logic_vector(to_unsigned(1,8) ,
39283	 => std_logic_vector(to_unsigned(2,8) ,
39284	 => std_logic_vector(to_unsigned(3,8) ,
39285	 => std_logic_vector(to_unsigned(5,8) ,
39286	 => std_logic_vector(to_unsigned(23,8) ,
39287	 => std_logic_vector(to_unsigned(29,8) ,
39288	 => std_logic_vector(to_unsigned(4,8) ,
39289	 => std_logic_vector(to_unsigned(0,8) ,
39290	 => std_logic_vector(to_unsigned(1,8) ,
39291	 => std_logic_vector(to_unsigned(3,8) ,
39292	 => std_logic_vector(to_unsigned(3,8) ,
39293	 => std_logic_vector(to_unsigned(3,8) ,
39294	 => std_logic_vector(to_unsigned(2,8) ,
39295	 => std_logic_vector(to_unsigned(3,8) ,
39296	 => std_logic_vector(to_unsigned(4,8) ,
39297	 => std_logic_vector(to_unsigned(3,8) ,
39298	 => std_logic_vector(to_unsigned(2,8) ,
39299	 => std_logic_vector(to_unsigned(3,8) ,
39300	 => std_logic_vector(to_unsigned(6,8) ,
39301	 => std_logic_vector(to_unsigned(2,8) ,
39302	 => std_logic_vector(to_unsigned(6,8) ,
39303	 => std_logic_vector(to_unsigned(19,8) ,
39304	 => std_logic_vector(to_unsigned(18,8) ,
39305	 => std_logic_vector(to_unsigned(13,8) ,
39306	 => std_logic_vector(to_unsigned(25,8) ,
39307	 => std_logic_vector(to_unsigned(48,8) ,
39308	 => std_logic_vector(to_unsigned(30,8) ,
39309	 => std_logic_vector(to_unsigned(38,8) ,
39310	 => std_logic_vector(to_unsigned(116,8) ,
39311	 => std_logic_vector(to_unsigned(156,8) ,
39312	 => std_logic_vector(to_unsigned(108,8) ,
39313	 => std_logic_vector(to_unsigned(44,8) ,
39314	 => std_logic_vector(to_unsigned(31,8) ,
39315	 => std_logic_vector(to_unsigned(56,8) ,
39316	 => std_logic_vector(to_unsigned(58,8) ,
39317	 => std_logic_vector(to_unsigned(59,8) ,
39318	 => std_logic_vector(to_unsigned(3,8) ,
39319	 => std_logic_vector(to_unsigned(0,8) ,
39320	 => std_logic_vector(to_unsigned(1,8) ,
39321	 => std_logic_vector(to_unsigned(1,8) ,
39322	 => std_logic_vector(to_unsigned(1,8) ,
39323	 => std_logic_vector(to_unsigned(1,8) ,
39324	 => std_logic_vector(to_unsigned(0,8) ,
39325	 => std_logic_vector(to_unsigned(2,8) ,
39326	 => std_logic_vector(to_unsigned(16,8) ,
39327	 => std_logic_vector(to_unsigned(20,8) ,
39328	 => std_logic_vector(to_unsigned(13,8) ,
39329	 => std_logic_vector(to_unsigned(9,8) ,
39330	 => std_logic_vector(to_unsigned(10,8) ,
39331	 => std_logic_vector(to_unsigned(13,8) ,
39332	 => std_logic_vector(to_unsigned(16,8) ,
39333	 => std_logic_vector(to_unsigned(18,8) ,
39334	 => std_logic_vector(to_unsigned(14,8) ,
39335	 => std_logic_vector(to_unsigned(2,8) ,
39336	 => std_logic_vector(to_unsigned(0,8) ,
39337	 => std_logic_vector(to_unsigned(1,8) ,
39338	 => std_logic_vector(to_unsigned(1,8) ,
39339	 => std_logic_vector(to_unsigned(1,8) ,
39340	 => std_logic_vector(to_unsigned(1,8) ,
39341	 => std_logic_vector(to_unsigned(4,8) ,
39342	 => std_logic_vector(to_unsigned(6,8) ,
39343	 => std_logic_vector(to_unsigned(11,8) ,
39344	 => std_logic_vector(to_unsigned(15,8) ,
39345	 => std_logic_vector(to_unsigned(22,8) ,
39346	 => std_logic_vector(to_unsigned(29,8) ,
39347	 => std_logic_vector(to_unsigned(45,8) ,
39348	 => std_logic_vector(to_unsigned(59,8) ,
39349	 => std_logic_vector(to_unsigned(65,8) ,
39350	 => std_logic_vector(to_unsigned(71,8) ,
39351	 => std_logic_vector(to_unsigned(78,8) ,
39352	 => std_logic_vector(to_unsigned(92,8) ,
39353	 => std_logic_vector(to_unsigned(82,8) ,
39354	 => std_logic_vector(to_unsigned(96,8) ,
39355	 => std_logic_vector(to_unsigned(124,8) ,
39356	 => std_logic_vector(to_unsigned(130,8) ,
39357	 => std_logic_vector(to_unsigned(92,8) ,
39358	 => std_logic_vector(to_unsigned(138,8) ,
39359	 => std_logic_vector(to_unsigned(173,8) ,
39360	 => std_logic_vector(to_unsigned(177,8) ,
39361	 => std_logic_vector(to_unsigned(146,8) ,
39362	 => std_logic_vector(to_unsigned(142,8) ,
39363	 => std_logic_vector(to_unsigned(138,8) ,
39364	 => std_logic_vector(to_unsigned(134,8) ,
39365	 => std_logic_vector(to_unsigned(134,8) ,
39366	 => std_logic_vector(to_unsigned(131,8) ,
39367	 => std_logic_vector(to_unsigned(128,8) ,
39368	 => std_logic_vector(to_unsigned(125,8) ,
39369	 => std_logic_vector(to_unsigned(131,8) ,
39370	 => std_logic_vector(to_unsigned(136,8) ,
39371	 => std_logic_vector(to_unsigned(138,8) ,
39372	 => std_logic_vector(to_unsigned(141,8) ,
39373	 => std_logic_vector(to_unsigned(138,8) ,
39374	 => std_logic_vector(to_unsigned(152,8) ,
39375	 => std_logic_vector(to_unsigned(81,8) ,
39376	 => std_logic_vector(to_unsigned(13,8) ,
39377	 => std_logic_vector(to_unsigned(42,8) ,
39378	 => std_logic_vector(to_unsigned(25,8) ,
39379	 => std_logic_vector(to_unsigned(0,8) ,
39380	 => std_logic_vector(to_unsigned(18,8) ,
39381	 => std_logic_vector(to_unsigned(159,8) ,
39382	 => std_logic_vector(to_unsigned(159,8) ,
39383	 => std_logic_vector(to_unsigned(152,8) ,
39384	 => std_logic_vector(to_unsigned(159,8) ,
39385	 => std_logic_vector(to_unsigned(157,8) ,
39386	 => std_logic_vector(to_unsigned(157,8) ,
39387	 => std_logic_vector(to_unsigned(156,8) ,
39388	 => std_logic_vector(to_unsigned(151,8) ,
39389	 => std_logic_vector(to_unsigned(149,8) ,
39390	 => std_logic_vector(to_unsigned(152,8) ,
39391	 => std_logic_vector(to_unsigned(170,8) ,
39392	 => std_logic_vector(to_unsigned(161,8) ,
39393	 => std_logic_vector(to_unsigned(29,8) ,
39394	 => std_logic_vector(to_unsigned(1,8) ,
39395	 => std_logic_vector(to_unsigned(2,8) ,
39396	 => std_logic_vector(to_unsigned(4,8) ,
39397	 => std_logic_vector(to_unsigned(7,8) ,
39398	 => std_logic_vector(to_unsigned(8,8) ,
39399	 => std_logic_vector(to_unsigned(4,8) ,
39400	 => std_logic_vector(to_unsigned(2,8) ,
39401	 => std_logic_vector(to_unsigned(4,8) ,
39402	 => std_logic_vector(to_unsigned(7,8) ,
39403	 => std_logic_vector(to_unsigned(45,8) ,
39404	 => std_logic_vector(to_unsigned(154,8) ,
39405	 => std_logic_vector(to_unsigned(159,8) ,
39406	 => std_logic_vector(to_unsigned(159,8) ,
39407	 => std_logic_vector(to_unsigned(159,8) ,
39408	 => std_logic_vector(to_unsigned(164,8) ,
39409	 => std_logic_vector(to_unsigned(161,8) ,
39410	 => std_logic_vector(to_unsigned(159,8) ,
39411	 => std_logic_vector(to_unsigned(157,8) ,
39412	 => std_logic_vector(to_unsigned(156,8) ,
39413	 => std_logic_vector(to_unsigned(154,8) ,
39414	 => std_logic_vector(to_unsigned(152,8) ,
39415	 => std_logic_vector(to_unsigned(152,8) ,
39416	 => std_logic_vector(to_unsigned(147,8) ,
39417	 => std_logic_vector(to_unsigned(131,8) ,
39418	 => std_logic_vector(to_unsigned(133,8) ,
39419	 => std_logic_vector(to_unsigned(133,8) ,
39420	 => std_logic_vector(to_unsigned(79,8) ,
39421	 => std_logic_vector(to_unsigned(4,8) ,
39422	 => std_logic_vector(to_unsigned(0,8) ,
39423	 => std_logic_vector(to_unsigned(1,8) ,
39424	 => std_logic_vector(to_unsigned(4,8) ,
39425	 => std_logic_vector(to_unsigned(3,8) ,
39426	 => std_logic_vector(to_unsigned(48,8) ,
39427	 => std_logic_vector(to_unsigned(183,8) ,
39428	 => std_logic_vector(to_unsigned(36,8) ,
39429	 => std_logic_vector(to_unsigned(1,8) ,
39430	 => std_logic_vector(to_unsigned(13,8) ,
39431	 => std_logic_vector(to_unsigned(27,8) ,
39432	 => std_logic_vector(to_unsigned(3,8) ,
39433	 => std_logic_vector(to_unsigned(1,8) ,
39434	 => std_logic_vector(to_unsigned(73,8) ,
39435	 => std_logic_vector(to_unsigned(91,8) ,
39436	 => std_logic_vector(to_unsigned(14,8) ,
39437	 => std_logic_vector(to_unsigned(6,8) ,
39438	 => std_logic_vector(to_unsigned(3,8) ,
39439	 => std_logic_vector(to_unsigned(3,8) ,
39440	 => std_logic_vector(to_unsigned(2,8) ,
39441	 => std_logic_vector(to_unsigned(2,8) ,
39442	 => std_logic_vector(to_unsigned(3,8) ,
39443	 => std_logic_vector(to_unsigned(2,8) ,
39444	 => std_logic_vector(to_unsigned(1,8) ,
39445	 => std_logic_vector(to_unsigned(1,8) ,
39446	 => std_logic_vector(to_unsigned(0,8) ,
39447	 => std_logic_vector(to_unsigned(0,8) ,
39448	 => std_logic_vector(to_unsigned(0,8) ,
39449	 => std_logic_vector(to_unsigned(0,8) ,
39450	 => std_logic_vector(to_unsigned(0,8) ,
39451	 => std_logic_vector(to_unsigned(0,8) ,
39452	 => std_logic_vector(to_unsigned(2,8) ,
39453	 => std_logic_vector(to_unsigned(4,8) ,
39454	 => std_logic_vector(to_unsigned(2,8) ,
39455	 => std_logic_vector(to_unsigned(3,8) ,
39456	 => std_logic_vector(to_unsigned(6,8) ,
39457	 => std_logic_vector(to_unsigned(4,8) ,
39458	 => std_logic_vector(to_unsigned(4,8) ,
39459	 => std_logic_vector(to_unsigned(2,8) ,
39460	 => std_logic_vector(to_unsigned(1,8) ,
39461	 => std_logic_vector(to_unsigned(2,8) ,
39462	 => std_logic_vector(to_unsigned(1,8) ,
39463	 => std_logic_vector(to_unsigned(4,8) ,
39464	 => std_logic_vector(to_unsigned(27,8) ,
39465	 => std_logic_vector(to_unsigned(8,8) ,
39466	 => std_logic_vector(to_unsigned(5,8) ,
39467	 => std_logic_vector(to_unsigned(4,8) ,
39468	 => std_logic_vector(to_unsigned(1,8) ,
39469	 => std_logic_vector(to_unsigned(0,8) ,
39470	 => std_logic_vector(to_unsigned(0,8) ,
39471	 => std_logic_vector(to_unsigned(0,8) ,
39472	 => std_logic_vector(to_unsigned(0,8) ,
39473	 => std_logic_vector(to_unsigned(1,8) ,
39474	 => std_logic_vector(to_unsigned(0,8) ,
39475	 => std_logic_vector(to_unsigned(18,8) ,
39476	 => std_logic_vector(to_unsigned(125,8) ,
39477	 => std_logic_vector(to_unsigned(122,8) ,
39478	 => std_logic_vector(to_unsigned(127,8) ,
39479	 => std_logic_vector(to_unsigned(86,8) ,
39480	 => std_logic_vector(to_unsigned(7,8) ,
39481	 => std_logic_vector(to_unsigned(1,8) ,
39482	 => std_logic_vector(to_unsigned(1,8) ,
39483	 => std_logic_vector(to_unsigned(3,8) ,
39484	 => std_logic_vector(to_unsigned(8,8) ,
39485	 => std_logic_vector(to_unsigned(5,8) ,
39486	 => std_logic_vector(to_unsigned(4,8) ,
39487	 => std_logic_vector(to_unsigned(3,8) ,
39488	 => std_logic_vector(to_unsigned(3,8) ,
39489	 => std_logic_vector(to_unsigned(2,8) ,
39490	 => std_logic_vector(to_unsigned(0,8) ,
39491	 => std_logic_vector(to_unsigned(2,8) ,
39492	 => std_logic_vector(to_unsigned(7,8) ,
39493	 => std_logic_vector(to_unsigned(6,8) ,
39494	 => std_logic_vector(to_unsigned(4,8) ,
39495	 => std_logic_vector(to_unsigned(4,8) ,
39496	 => std_logic_vector(to_unsigned(5,8) ,
39497	 => std_logic_vector(to_unsigned(7,8) ,
39498	 => std_logic_vector(to_unsigned(6,8) ,
39499	 => std_logic_vector(to_unsigned(4,8) ,
39500	 => std_logic_vector(to_unsigned(4,8) ,
39501	 => std_logic_vector(to_unsigned(5,8) ,
39502	 => std_logic_vector(to_unsigned(3,8) ,
39503	 => std_logic_vector(to_unsigned(1,8) ,
39504	 => std_logic_vector(to_unsigned(0,8) ,
39505	 => std_logic_vector(to_unsigned(0,8) ,
39506	 => std_logic_vector(to_unsigned(1,8) ,
39507	 => std_logic_vector(to_unsigned(1,8) ,
39508	 => std_logic_vector(to_unsigned(1,8) ,
39509	 => std_logic_vector(to_unsigned(2,8) ,
39510	 => std_logic_vector(to_unsigned(2,8) ,
39511	 => std_logic_vector(to_unsigned(2,8) ,
39512	 => std_logic_vector(to_unsigned(5,8) ,
39513	 => std_logic_vector(to_unsigned(9,8) ,
39514	 => std_logic_vector(to_unsigned(8,8) ,
39515	 => std_logic_vector(to_unsigned(3,8) ,
39516	 => std_logic_vector(to_unsigned(1,8) ,
39517	 => std_logic_vector(to_unsigned(0,8) ,
39518	 => std_logic_vector(to_unsigned(2,8) ,
39519	 => std_logic_vector(to_unsigned(6,8) ,
39520	 => std_logic_vector(to_unsigned(9,8) ,
39521	 => std_logic_vector(to_unsigned(7,8) ,
39522	 => std_logic_vector(to_unsigned(8,8) ,
39523	 => std_logic_vector(to_unsigned(6,8) ,
39524	 => std_logic_vector(to_unsigned(3,8) ,
39525	 => std_logic_vector(to_unsigned(5,8) ,
39526	 => std_logic_vector(to_unsigned(3,8) ,
39527	 => std_logic_vector(to_unsigned(1,8) ,
39528	 => std_logic_vector(to_unsigned(1,8) ,
39529	 => std_logic_vector(to_unsigned(1,8) ,
39530	 => std_logic_vector(to_unsigned(1,8) ,
39531	 => std_logic_vector(to_unsigned(1,8) ,
39532	 => std_logic_vector(to_unsigned(1,8) ,
39533	 => std_logic_vector(to_unsigned(1,8) ,
39534	 => std_logic_vector(to_unsigned(1,8) ,
39535	 => std_logic_vector(to_unsigned(3,8) ,
39536	 => std_logic_vector(to_unsigned(5,8) ,
39537	 => std_logic_vector(to_unsigned(3,8) ,
39538	 => std_logic_vector(to_unsigned(2,8) ,
39539	 => std_logic_vector(to_unsigned(3,8) ,
39540	 => std_logic_vector(to_unsigned(3,8) ,
39541	 => std_logic_vector(to_unsigned(1,8) ,
39542	 => std_logic_vector(to_unsigned(1,8) ,
39543	 => std_logic_vector(to_unsigned(3,8) ,
39544	 => std_logic_vector(to_unsigned(5,8) ,
39545	 => std_logic_vector(to_unsigned(3,8) ,
39546	 => std_logic_vector(to_unsigned(3,8) ,
39547	 => std_logic_vector(to_unsigned(2,8) ,
39548	 => std_logic_vector(to_unsigned(2,8) ,
39549	 => std_logic_vector(to_unsigned(3,8) ,
39550	 => std_logic_vector(to_unsigned(1,8) ,
39551	 => std_logic_vector(to_unsigned(0,8) ,
39552	 => std_logic_vector(to_unsigned(0,8) ,
39553	 => std_logic_vector(to_unsigned(0,8) ,
39554	 => std_logic_vector(to_unsigned(0,8) ,
39555	 => std_logic_vector(to_unsigned(1,8) ,
39556	 => std_logic_vector(to_unsigned(1,8) ,
39557	 => std_logic_vector(to_unsigned(1,8) ,
39558	 => std_logic_vector(to_unsigned(1,8) ,
39559	 => std_logic_vector(to_unsigned(1,8) ,
39560	 => std_logic_vector(to_unsigned(2,8) ,
39561	 => std_logic_vector(to_unsigned(3,8) ,
39562	 => std_logic_vector(to_unsigned(2,8) ,
39563	 => std_logic_vector(to_unsigned(2,8) ,
39564	 => std_logic_vector(to_unsigned(2,8) ,
39565	 => std_logic_vector(to_unsigned(2,8) ,
39566	 => std_logic_vector(to_unsigned(2,8) ,
39567	 => std_logic_vector(to_unsigned(4,8) ,
39568	 => std_logic_vector(to_unsigned(4,8) ,
39569	 => std_logic_vector(to_unsigned(6,8) ,
39570	 => std_logic_vector(to_unsigned(6,8) ,
39571	 => std_logic_vector(to_unsigned(5,8) ,
39572	 => std_logic_vector(to_unsigned(4,8) ,
39573	 => std_logic_vector(to_unsigned(1,8) ,
39574	 => std_logic_vector(to_unsigned(31,8) ,
39575	 => std_logic_vector(to_unsigned(125,8) ,
39576	 => std_logic_vector(to_unsigned(99,8) ,
39577	 => std_logic_vector(to_unsigned(49,8) ,
39578	 => std_logic_vector(to_unsigned(36,8) ,
39579	 => std_logic_vector(to_unsigned(37,8) ,
39580	 => std_logic_vector(to_unsigned(12,8) ,
39581	 => std_logic_vector(to_unsigned(3,8) ,
39582	 => std_logic_vector(to_unsigned(0,8) ,
39583	 => std_logic_vector(to_unsigned(0,8) ,
39584	 => std_logic_vector(to_unsigned(0,8) ,
39585	 => std_logic_vector(to_unsigned(1,8) ,
39586	 => std_logic_vector(to_unsigned(1,8) ,
39587	 => std_logic_vector(to_unsigned(2,8) ,
39588	 => std_logic_vector(to_unsigned(1,8) ,
39589	 => std_logic_vector(to_unsigned(4,8) ,
39590	 => std_logic_vector(to_unsigned(77,8) ,
39591	 => std_logic_vector(to_unsigned(108,8) ,
39592	 => std_logic_vector(to_unsigned(108,8) ,
39593	 => std_logic_vector(to_unsigned(136,8) ,
39594	 => std_logic_vector(to_unsigned(93,8) ,
39595	 => std_logic_vector(to_unsigned(17,8) ,
39596	 => std_logic_vector(to_unsigned(8,8) ,
39597	 => std_logic_vector(to_unsigned(2,8) ,
39598	 => std_logic_vector(to_unsigned(1,8) ,
39599	 => std_logic_vector(to_unsigned(2,8) ,
39600	 => std_logic_vector(to_unsigned(6,8) ,
39601	 => std_logic_vector(to_unsigned(4,8) ,
39602	 => std_logic_vector(to_unsigned(1,8) ,
39603	 => std_logic_vector(to_unsigned(2,8) ,
39604	 => std_logic_vector(to_unsigned(4,8) ,
39605	 => std_logic_vector(to_unsigned(4,8) ,
39606	 => std_logic_vector(to_unsigned(16,8) ,
39607	 => std_logic_vector(to_unsigned(29,8) ,
39608	 => std_logic_vector(to_unsigned(12,8) ,
39609	 => std_logic_vector(to_unsigned(1,8) ,
39610	 => std_logic_vector(to_unsigned(2,8) ,
39611	 => std_logic_vector(to_unsigned(2,8) ,
39612	 => std_logic_vector(to_unsigned(3,8) ,
39613	 => std_logic_vector(to_unsigned(3,8) ,
39614	 => std_logic_vector(to_unsigned(2,8) ,
39615	 => std_logic_vector(to_unsigned(2,8) ,
39616	 => std_logic_vector(to_unsigned(3,8) ,
39617	 => std_logic_vector(to_unsigned(2,8) ,
39618	 => std_logic_vector(to_unsigned(2,8) ,
39619	 => std_logic_vector(to_unsigned(4,8) ,
39620	 => std_logic_vector(to_unsigned(7,8) ,
39621	 => std_logic_vector(to_unsigned(2,8) ,
39622	 => std_logic_vector(to_unsigned(4,8) ,
39623	 => std_logic_vector(to_unsigned(14,8) ,
39624	 => std_logic_vector(to_unsigned(20,8) ,
39625	 => std_logic_vector(to_unsigned(8,8) ,
39626	 => std_logic_vector(to_unsigned(38,8) ,
39627	 => std_logic_vector(to_unsigned(86,8) ,
39628	 => std_logic_vector(to_unsigned(17,8) ,
39629	 => std_logic_vector(to_unsigned(9,8) ,
39630	 => std_logic_vector(to_unsigned(23,8) ,
39631	 => std_logic_vector(to_unsigned(116,8) ,
39632	 => std_logic_vector(to_unsigned(139,8) ,
39633	 => std_logic_vector(to_unsigned(81,8) ,
39634	 => std_logic_vector(to_unsigned(24,8) ,
39635	 => std_logic_vector(to_unsigned(18,8) ,
39636	 => std_logic_vector(to_unsigned(7,8) ,
39637	 => std_logic_vector(to_unsigned(2,8) ,
39638	 => std_logic_vector(to_unsigned(1,8) ,
39639	 => std_logic_vector(to_unsigned(0,8) ,
39640	 => std_logic_vector(to_unsigned(1,8) ,
39641	 => std_logic_vector(to_unsigned(1,8) ,
39642	 => std_logic_vector(to_unsigned(2,8) ,
39643	 => std_logic_vector(to_unsigned(5,8) ,
39644	 => std_logic_vector(to_unsigned(4,8) ,
39645	 => std_logic_vector(to_unsigned(5,8) ,
39646	 => std_logic_vector(to_unsigned(10,8) ,
39647	 => std_logic_vector(to_unsigned(15,8) ,
39648	 => std_logic_vector(to_unsigned(12,8) ,
39649	 => std_logic_vector(to_unsigned(17,8) ,
39650	 => std_logic_vector(to_unsigned(27,8) ,
39651	 => std_logic_vector(to_unsigned(20,8) ,
39652	 => std_logic_vector(to_unsigned(13,8) ,
39653	 => std_logic_vector(to_unsigned(13,8) ,
39654	 => std_logic_vector(to_unsigned(17,8) ,
39655	 => std_logic_vector(to_unsigned(11,8) ,
39656	 => std_logic_vector(to_unsigned(2,8) ,
39657	 => std_logic_vector(to_unsigned(0,8) ,
39658	 => std_logic_vector(to_unsigned(0,8) ,
39659	 => std_logic_vector(to_unsigned(0,8) ,
39660	 => std_logic_vector(to_unsigned(0,8) ,
39661	 => std_logic_vector(to_unsigned(0,8) ,
39662	 => std_logic_vector(to_unsigned(0,8) ,
39663	 => std_logic_vector(to_unsigned(0,8) ,
39664	 => std_logic_vector(to_unsigned(0,8) ,
39665	 => std_logic_vector(to_unsigned(0,8) ,
39666	 => std_logic_vector(to_unsigned(0,8) ,
39667	 => std_logic_vector(to_unsigned(0,8) ,
39668	 => std_logic_vector(to_unsigned(0,8) ,
39669	 => std_logic_vector(to_unsigned(1,8) ,
39670	 => std_logic_vector(to_unsigned(2,8) ,
39671	 => std_logic_vector(to_unsigned(2,8) ,
39672	 => std_logic_vector(to_unsigned(5,8) ,
39673	 => std_logic_vector(to_unsigned(6,8) ,
39674	 => std_logic_vector(to_unsigned(7,8) ,
39675	 => std_logic_vector(to_unsigned(12,8) ,
39676	 => std_logic_vector(to_unsigned(18,8) ,
39677	 => std_logic_vector(to_unsigned(20,8) ,
39678	 => std_logic_vector(to_unsigned(37,8) ,
39679	 => std_logic_vector(to_unsigned(45,8) ,
39680	 => std_logic_vector(to_unsigned(64,8) ,
39681	 => std_logic_vector(to_unsigned(146,8) ,
39682	 => std_logic_vector(to_unsigned(146,8) ,
39683	 => std_logic_vector(to_unsigned(142,8) ,
39684	 => std_logic_vector(to_unsigned(128,8) ,
39685	 => std_logic_vector(to_unsigned(131,8) ,
39686	 => std_logic_vector(to_unsigned(128,8) ,
39687	 => std_logic_vector(to_unsigned(121,8) ,
39688	 => std_logic_vector(to_unsigned(121,8) ,
39689	 => std_logic_vector(to_unsigned(127,8) ,
39690	 => std_logic_vector(to_unsigned(124,8) ,
39691	 => std_logic_vector(to_unsigned(122,8) ,
39692	 => std_logic_vector(to_unsigned(125,8) ,
39693	 => std_logic_vector(to_unsigned(133,8) ,
39694	 => std_logic_vector(to_unsigned(142,8) ,
39695	 => std_logic_vector(to_unsigned(115,8) ,
39696	 => std_logic_vector(to_unsigned(10,8) ,
39697	 => std_logic_vector(to_unsigned(10,8) ,
39698	 => std_logic_vector(to_unsigned(7,8) ,
39699	 => std_logic_vector(to_unsigned(1,8) ,
39700	 => std_logic_vector(to_unsigned(62,8) ,
39701	 => std_logic_vector(to_unsigned(170,8) ,
39702	 => std_logic_vector(to_unsigned(147,8) ,
39703	 => std_logic_vector(to_unsigned(152,8) ,
39704	 => std_logic_vector(to_unsigned(147,8) ,
39705	 => std_logic_vector(to_unsigned(154,8) ,
39706	 => std_logic_vector(to_unsigned(159,8) ,
39707	 => std_logic_vector(to_unsigned(152,8) ,
39708	 => std_logic_vector(to_unsigned(142,8) ,
39709	 => std_logic_vector(to_unsigned(144,8) ,
39710	 => std_logic_vector(to_unsigned(149,8) ,
39711	 => std_logic_vector(to_unsigned(157,8) ,
39712	 => std_logic_vector(to_unsigned(151,8) ,
39713	 => std_logic_vector(to_unsigned(16,8) ,
39714	 => std_logic_vector(to_unsigned(1,8) ,
39715	 => std_logic_vector(to_unsigned(1,8) ,
39716	 => std_logic_vector(to_unsigned(1,8) ,
39717	 => std_logic_vector(to_unsigned(1,8) ,
39718	 => std_logic_vector(to_unsigned(1,8) ,
39719	 => std_logic_vector(to_unsigned(4,8) ,
39720	 => std_logic_vector(to_unsigned(9,8) ,
39721	 => std_logic_vector(to_unsigned(23,8) ,
39722	 => std_logic_vector(to_unsigned(76,8) ,
39723	 => std_logic_vector(to_unsigned(157,8) ,
39724	 => std_logic_vector(to_unsigned(170,8) ,
39725	 => std_logic_vector(to_unsigned(154,8) ,
39726	 => std_logic_vector(to_unsigned(159,8) ,
39727	 => std_logic_vector(to_unsigned(161,8) ,
39728	 => std_logic_vector(to_unsigned(157,8) ,
39729	 => std_logic_vector(to_unsigned(161,8) ,
39730	 => std_logic_vector(to_unsigned(157,8) ,
39731	 => std_logic_vector(to_unsigned(156,8) ,
39732	 => std_logic_vector(to_unsigned(157,8) ,
39733	 => std_logic_vector(to_unsigned(156,8) ,
39734	 => std_logic_vector(to_unsigned(151,8) ,
39735	 => std_logic_vector(to_unsigned(152,8) ,
39736	 => std_logic_vector(to_unsigned(157,8) ,
39737	 => std_logic_vector(to_unsigned(152,8) ,
39738	 => std_logic_vector(to_unsigned(151,8) ,
39739	 => std_logic_vector(to_unsigned(173,8) ,
39740	 => std_logic_vector(to_unsigned(142,8) ,
39741	 => std_logic_vector(to_unsigned(7,8) ,
39742	 => std_logic_vector(to_unsigned(0,8) ,
39743	 => std_logic_vector(to_unsigned(1,8) ,
39744	 => std_logic_vector(to_unsigned(4,8) ,
39745	 => std_logic_vector(to_unsigned(3,8) ,
39746	 => std_logic_vector(to_unsigned(12,8) ,
39747	 => std_logic_vector(to_unsigned(134,8) ,
39748	 => std_logic_vector(to_unsigned(121,8) ,
39749	 => std_logic_vector(to_unsigned(45,8) ,
39750	 => std_logic_vector(to_unsigned(27,8) ,
39751	 => std_logic_vector(to_unsigned(17,8) ,
39752	 => std_logic_vector(to_unsigned(15,8) ,
39753	 => std_logic_vector(to_unsigned(51,8) ,
39754	 => std_logic_vector(to_unsigned(133,8) ,
39755	 => std_logic_vector(to_unsigned(136,8) ,
39756	 => std_logic_vector(to_unsigned(97,8) ,
39757	 => std_logic_vector(to_unsigned(45,8) ,
39758	 => std_logic_vector(to_unsigned(20,8) ,
39759	 => std_logic_vector(to_unsigned(11,8) ,
39760	 => std_logic_vector(to_unsigned(6,8) ,
39761	 => std_logic_vector(to_unsigned(3,8) ,
39762	 => std_logic_vector(to_unsigned(1,8) ,
39763	 => std_logic_vector(to_unsigned(1,8) ,
39764	 => std_logic_vector(to_unsigned(2,8) ,
39765	 => std_logic_vector(to_unsigned(2,8) ,
39766	 => std_logic_vector(to_unsigned(18,8) ,
39767	 => std_logic_vector(to_unsigned(61,8) ,
39768	 => std_logic_vector(to_unsigned(44,8) ,
39769	 => std_logic_vector(to_unsigned(38,8) ,
39770	 => std_logic_vector(to_unsigned(26,8) ,
39771	 => std_logic_vector(to_unsigned(13,8) ,
39772	 => std_logic_vector(to_unsigned(4,8) ,
39773	 => std_logic_vector(to_unsigned(5,8) ,
39774	 => std_logic_vector(to_unsigned(4,8) ,
39775	 => std_logic_vector(to_unsigned(5,8) ,
39776	 => std_logic_vector(to_unsigned(5,8) ,
39777	 => std_logic_vector(to_unsigned(4,8) ,
39778	 => std_logic_vector(to_unsigned(5,8) ,
39779	 => std_logic_vector(to_unsigned(3,8) ,
39780	 => std_logic_vector(to_unsigned(2,8) ,
39781	 => std_logic_vector(to_unsigned(1,8) ,
39782	 => std_logic_vector(to_unsigned(0,8) ,
39783	 => std_logic_vector(to_unsigned(1,8) ,
39784	 => std_logic_vector(to_unsigned(30,8) ,
39785	 => std_logic_vector(to_unsigned(25,8) ,
39786	 => std_logic_vector(to_unsigned(22,8) ,
39787	 => std_logic_vector(to_unsigned(15,8) ,
39788	 => std_logic_vector(to_unsigned(2,8) ,
39789	 => std_logic_vector(to_unsigned(0,8) ,
39790	 => std_logic_vector(to_unsigned(0,8) ,
39791	 => std_logic_vector(to_unsigned(0,8) ,
39792	 => std_logic_vector(to_unsigned(0,8) ,
39793	 => std_logic_vector(to_unsigned(1,8) ,
39794	 => std_logic_vector(to_unsigned(1,8) ,
39795	 => std_logic_vector(to_unsigned(4,8) ,
39796	 => std_logic_vector(to_unsigned(72,8) ,
39797	 => std_logic_vector(to_unsigned(131,8) ,
39798	 => std_logic_vector(to_unsigned(103,8) ,
39799	 => std_logic_vector(to_unsigned(114,8) ,
39800	 => std_logic_vector(to_unsigned(25,8) ,
39801	 => std_logic_vector(to_unsigned(2,8) ,
39802	 => std_logic_vector(to_unsigned(3,8) ,
39803	 => std_logic_vector(to_unsigned(4,8) ,
39804	 => std_logic_vector(to_unsigned(8,8) ,
39805	 => std_logic_vector(to_unsigned(5,8) ,
39806	 => std_logic_vector(to_unsigned(2,8) ,
39807	 => std_logic_vector(to_unsigned(4,8) ,
39808	 => std_logic_vector(to_unsigned(6,8) ,
39809	 => std_logic_vector(to_unsigned(2,8) ,
39810	 => std_logic_vector(to_unsigned(0,8) ,
39811	 => std_logic_vector(to_unsigned(2,8) ,
39812	 => std_logic_vector(to_unsigned(5,8) ,
39813	 => std_logic_vector(to_unsigned(6,8) ,
39814	 => std_logic_vector(to_unsigned(4,8) ,
39815	 => std_logic_vector(to_unsigned(4,8) ,
39816	 => std_logic_vector(to_unsigned(5,8) ,
39817	 => std_logic_vector(to_unsigned(3,8) ,
39818	 => std_logic_vector(to_unsigned(2,8) ,
39819	 => std_logic_vector(to_unsigned(2,8) ,
39820	 => std_logic_vector(to_unsigned(4,8) ,
39821	 => std_logic_vector(to_unsigned(6,8) ,
39822	 => std_logic_vector(to_unsigned(2,8) ,
39823	 => std_logic_vector(to_unsigned(1,8) ,
39824	 => std_logic_vector(to_unsigned(1,8) ,
39825	 => std_logic_vector(to_unsigned(0,8) ,
39826	 => std_logic_vector(to_unsigned(1,8) ,
39827	 => std_logic_vector(to_unsigned(1,8) ,
39828	 => std_logic_vector(to_unsigned(2,8) ,
39829	 => std_logic_vector(to_unsigned(3,8) ,
39830	 => std_logic_vector(to_unsigned(2,8) ,
39831	 => std_logic_vector(to_unsigned(2,8) ,
39832	 => std_logic_vector(to_unsigned(7,8) ,
39833	 => std_logic_vector(to_unsigned(11,8) ,
39834	 => std_logic_vector(to_unsigned(8,8) ,
39835	 => std_logic_vector(to_unsigned(4,8) ,
39836	 => std_logic_vector(to_unsigned(1,8) ,
39837	 => std_logic_vector(to_unsigned(0,8) ,
39838	 => std_logic_vector(to_unsigned(3,8) ,
39839	 => std_logic_vector(to_unsigned(5,8) ,
39840	 => std_logic_vector(to_unsigned(7,8) ,
39841	 => std_logic_vector(to_unsigned(6,8) ,
39842	 => std_logic_vector(to_unsigned(9,8) ,
39843	 => std_logic_vector(to_unsigned(9,8) ,
39844	 => std_logic_vector(to_unsigned(3,8) ,
39845	 => std_logic_vector(to_unsigned(5,8) ,
39846	 => std_logic_vector(to_unsigned(3,8) ,
39847	 => std_logic_vector(to_unsigned(0,8) ,
39848	 => std_logic_vector(to_unsigned(0,8) ,
39849	 => std_logic_vector(to_unsigned(0,8) ,
39850	 => std_logic_vector(to_unsigned(1,8) ,
39851	 => std_logic_vector(to_unsigned(1,8) ,
39852	 => std_logic_vector(to_unsigned(1,8) ,
39853	 => std_logic_vector(to_unsigned(2,8) ,
39854	 => std_logic_vector(to_unsigned(2,8) ,
39855	 => std_logic_vector(to_unsigned(3,8) ,
39856	 => std_logic_vector(to_unsigned(5,8) ,
39857	 => std_logic_vector(to_unsigned(3,8) ,
39858	 => std_logic_vector(to_unsigned(4,8) ,
39859	 => std_logic_vector(to_unsigned(5,8) ,
39860	 => std_logic_vector(to_unsigned(3,8) ,
39861	 => std_logic_vector(to_unsigned(1,8) ,
39862	 => std_logic_vector(to_unsigned(1,8) ,
39863	 => std_logic_vector(to_unsigned(3,8) ,
39864	 => std_logic_vector(to_unsigned(4,8) ,
39865	 => std_logic_vector(to_unsigned(3,8) ,
39866	 => std_logic_vector(to_unsigned(3,8) ,
39867	 => std_logic_vector(to_unsigned(3,8) ,
39868	 => std_logic_vector(to_unsigned(2,8) ,
39869	 => std_logic_vector(to_unsigned(2,8) ,
39870	 => std_logic_vector(to_unsigned(2,8) ,
39871	 => std_logic_vector(to_unsigned(1,8) ,
39872	 => std_logic_vector(to_unsigned(0,8) ,
39873	 => std_logic_vector(to_unsigned(0,8) ,
39874	 => std_logic_vector(to_unsigned(0,8) ,
39875	 => std_logic_vector(to_unsigned(0,8) ,
39876	 => std_logic_vector(to_unsigned(1,8) ,
39877	 => std_logic_vector(to_unsigned(1,8) ,
39878	 => std_logic_vector(to_unsigned(1,8) ,
39879	 => std_logic_vector(to_unsigned(1,8) ,
39880	 => std_logic_vector(to_unsigned(2,8) ,
39881	 => std_logic_vector(to_unsigned(2,8) ,
39882	 => std_logic_vector(to_unsigned(2,8) ,
39883	 => std_logic_vector(to_unsigned(2,8) ,
39884	 => std_logic_vector(to_unsigned(2,8) ,
39885	 => std_logic_vector(to_unsigned(1,8) ,
39886	 => std_logic_vector(to_unsigned(1,8) ,
39887	 => std_logic_vector(to_unsigned(3,8) ,
39888	 => std_logic_vector(to_unsigned(4,8) ,
39889	 => std_logic_vector(to_unsigned(7,8) ,
39890	 => std_logic_vector(to_unsigned(6,8) ,
39891	 => std_logic_vector(to_unsigned(5,8) ,
39892	 => std_logic_vector(to_unsigned(4,8) ,
39893	 => std_logic_vector(to_unsigned(1,8) ,
39894	 => std_logic_vector(to_unsigned(42,8) ,
39895	 => std_logic_vector(to_unsigned(133,8) ,
39896	 => std_logic_vector(to_unsigned(103,8) ,
39897	 => std_logic_vector(to_unsigned(58,8) ,
39898	 => std_logic_vector(to_unsigned(41,8) ,
39899	 => std_logic_vector(to_unsigned(30,8) ,
39900	 => std_logic_vector(to_unsigned(10,8) ,
39901	 => std_logic_vector(to_unsigned(1,8) ,
39902	 => std_logic_vector(to_unsigned(0,8) ,
39903	 => std_logic_vector(to_unsigned(0,8) ,
39904	 => std_logic_vector(to_unsigned(0,8) ,
39905	 => std_logic_vector(to_unsigned(1,8) ,
39906	 => std_logic_vector(to_unsigned(2,8) ,
39907	 => std_logic_vector(to_unsigned(2,8) ,
39908	 => std_logic_vector(to_unsigned(1,8) ,
39909	 => std_logic_vector(to_unsigned(5,8) ,
39910	 => std_logic_vector(to_unsigned(67,8) ,
39911	 => std_logic_vector(to_unsigned(109,8) ,
39912	 => std_logic_vector(to_unsigned(111,8) ,
39913	 => std_logic_vector(to_unsigned(131,8) ,
39914	 => std_logic_vector(to_unsigned(116,8) ,
39915	 => std_logic_vector(to_unsigned(34,8) ,
39916	 => std_logic_vector(to_unsigned(9,8) ,
39917	 => std_logic_vector(to_unsigned(3,8) ,
39918	 => std_logic_vector(to_unsigned(1,8) ,
39919	 => std_logic_vector(to_unsigned(2,8) ,
39920	 => std_logic_vector(to_unsigned(4,8) ,
39921	 => std_logic_vector(to_unsigned(4,8) ,
39922	 => std_logic_vector(to_unsigned(2,8) ,
39923	 => std_logic_vector(to_unsigned(1,8) ,
39924	 => std_logic_vector(to_unsigned(3,8) ,
39925	 => std_logic_vector(to_unsigned(4,8) ,
39926	 => std_logic_vector(to_unsigned(7,8) ,
39927	 => std_logic_vector(to_unsigned(14,8) ,
39928	 => std_logic_vector(to_unsigned(16,8) ,
39929	 => std_logic_vector(to_unsigned(1,8) ,
39930	 => std_logic_vector(to_unsigned(1,8) ,
39931	 => std_logic_vector(to_unsigned(2,8) ,
39932	 => std_logic_vector(to_unsigned(3,8) ,
39933	 => std_logic_vector(to_unsigned(2,8) ,
39934	 => std_logic_vector(to_unsigned(3,8) ,
39935	 => std_logic_vector(to_unsigned(2,8) ,
39936	 => std_logic_vector(to_unsigned(2,8) ,
39937	 => std_logic_vector(to_unsigned(2,8) ,
39938	 => std_logic_vector(to_unsigned(2,8) ,
39939	 => std_logic_vector(to_unsigned(5,8) ,
39940	 => std_logic_vector(to_unsigned(5,8) ,
39941	 => std_logic_vector(to_unsigned(2,8) ,
39942	 => std_logic_vector(to_unsigned(3,8) ,
39943	 => std_logic_vector(to_unsigned(9,8) ,
39944	 => std_logic_vector(to_unsigned(12,8) ,
39945	 => std_logic_vector(to_unsigned(7,8) ,
39946	 => std_logic_vector(to_unsigned(23,8) ,
39947	 => std_logic_vector(to_unsigned(71,8) ,
39948	 => std_logic_vector(to_unsigned(41,8) ,
39949	 => std_logic_vector(to_unsigned(18,8) ,
39950	 => std_logic_vector(to_unsigned(35,8) ,
39951	 => std_logic_vector(to_unsigned(141,8) ,
39952	 => std_logic_vector(to_unsigned(157,8) ,
39953	 => std_logic_vector(to_unsigned(122,8) ,
39954	 => std_logic_vector(to_unsigned(93,8) ,
39955	 => std_logic_vector(to_unsigned(39,8) ,
39956	 => std_logic_vector(to_unsigned(1,8) ,
39957	 => std_logic_vector(to_unsigned(0,8) ,
39958	 => std_logic_vector(to_unsigned(1,8) ,
39959	 => std_logic_vector(to_unsigned(1,8) ,
39960	 => std_logic_vector(to_unsigned(1,8) ,
39961	 => std_logic_vector(to_unsigned(1,8) ,
39962	 => std_logic_vector(to_unsigned(3,8) ,
39963	 => std_logic_vector(to_unsigned(14,8) ,
39964	 => std_logic_vector(to_unsigned(7,8) ,
39965	 => std_logic_vector(to_unsigned(2,8) ,
39966	 => std_logic_vector(to_unsigned(4,8) ,
39967	 => std_logic_vector(to_unsigned(6,8) ,
39968	 => std_logic_vector(to_unsigned(13,8) ,
39969	 => std_logic_vector(to_unsigned(17,8) ,
39970	 => std_logic_vector(to_unsigned(20,8) ,
39971	 => std_logic_vector(to_unsigned(18,8) ,
39972	 => std_logic_vector(to_unsigned(14,8) ,
39973	 => std_logic_vector(to_unsigned(9,8) ,
39974	 => std_logic_vector(to_unsigned(9,8) ,
39975	 => std_logic_vector(to_unsigned(12,8) ,
39976	 => std_logic_vector(to_unsigned(1,8) ,
39977	 => std_logic_vector(to_unsigned(0,8) ,
39978	 => std_logic_vector(to_unsigned(0,8) ,
39979	 => std_logic_vector(to_unsigned(0,8) ,
39980	 => std_logic_vector(to_unsigned(0,8) ,
39981	 => std_logic_vector(to_unsigned(1,8) ,
39982	 => std_logic_vector(to_unsigned(1,8) ,
39983	 => std_logic_vector(to_unsigned(0,8) ,
39984	 => std_logic_vector(to_unsigned(0,8) ,
39985	 => std_logic_vector(to_unsigned(0,8) ,
39986	 => std_logic_vector(to_unsigned(0,8) ,
39987	 => std_logic_vector(to_unsigned(0,8) ,
39988	 => std_logic_vector(to_unsigned(0,8) ,
39989	 => std_logic_vector(to_unsigned(0,8) ,
39990	 => std_logic_vector(to_unsigned(0,8) ,
39991	 => std_logic_vector(to_unsigned(0,8) ,
39992	 => std_logic_vector(to_unsigned(0,8) ,
39993	 => std_logic_vector(to_unsigned(0,8) ,
39994	 => std_logic_vector(to_unsigned(0,8) ,
39995	 => std_logic_vector(to_unsigned(0,8) ,
39996	 => std_logic_vector(to_unsigned(0,8) ,
39997	 => std_logic_vector(to_unsigned(0,8) ,
39998	 => std_logic_vector(to_unsigned(1,8) ,
39999	 => std_logic_vector(to_unsigned(0,8) ,
40000	 => std_logic_vector(to_unsigned(1,8) ,
40001	 => std_logic_vector(to_unsigned(138,8) ,
40002	 => std_logic_vector(to_unsigned(142,8) ,
40003	 => std_logic_vector(to_unsigned(139,8) ,
40004	 => std_logic_vector(to_unsigned(124,8) ,
40005	 => std_logic_vector(to_unsigned(124,8) ,
40006	 => std_logic_vector(to_unsigned(119,8) ,
40007	 => std_logic_vector(to_unsigned(115,8) ,
40008	 => std_logic_vector(to_unsigned(115,8) ,
40009	 => std_logic_vector(to_unsigned(118,8) ,
40010	 => std_logic_vector(to_unsigned(111,8) ,
40011	 => std_logic_vector(to_unsigned(108,8) ,
40012	 => std_logic_vector(to_unsigned(111,8) ,
40013	 => std_logic_vector(to_unsigned(115,8) ,
40014	 => std_logic_vector(to_unsigned(121,8) ,
40015	 => std_logic_vector(to_unsigned(128,8) ,
40016	 => std_logic_vector(to_unsigned(29,8) ,
40017	 => std_logic_vector(to_unsigned(1,8) ,
40018	 => std_logic_vector(to_unsigned(1,8) ,
40019	 => std_logic_vector(to_unsigned(25,8) ,
40020	 => std_logic_vector(to_unsigned(133,8) ,
40021	 => std_logic_vector(to_unsigned(144,8) ,
40022	 => std_logic_vector(to_unsigned(149,8) ,
40023	 => std_logic_vector(to_unsigned(149,8) ,
40024	 => std_logic_vector(to_unsigned(141,8) ,
40025	 => std_logic_vector(to_unsigned(147,8) ,
40026	 => std_logic_vector(to_unsigned(159,8) ,
40027	 => std_logic_vector(to_unsigned(147,8) ,
40028	 => std_logic_vector(to_unsigned(141,8) ,
40029	 => std_logic_vector(to_unsigned(141,8) ,
40030	 => std_logic_vector(to_unsigned(142,8) ,
40031	 => std_logic_vector(to_unsigned(177,8) ,
40032	 => std_logic_vector(to_unsigned(76,8) ,
40033	 => std_logic_vector(to_unsigned(3,8) ,
40034	 => std_logic_vector(to_unsigned(7,8) ,
40035	 => std_logic_vector(to_unsigned(7,8) ,
40036	 => std_logic_vector(to_unsigned(4,8) ,
40037	 => std_logic_vector(to_unsigned(1,8) ,
40038	 => std_logic_vector(to_unsigned(1,8) ,
40039	 => std_logic_vector(to_unsigned(3,8) ,
40040	 => std_logic_vector(to_unsigned(2,8) ,
40041	 => std_logic_vector(to_unsigned(60,8) ,
40042	 => std_logic_vector(to_unsigned(196,8) ,
40043	 => std_logic_vector(to_unsigned(161,8) ,
40044	 => std_logic_vector(to_unsigned(152,8) ,
40045	 => std_logic_vector(to_unsigned(157,8) ,
40046	 => std_logic_vector(to_unsigned(157,8) ,
40047	 => std_logic_vector(to_unsigned(157,8) ,
40048	 => std_logic_vector(to_unsigned(142,8) ,
40049	 => std_logic_vector(to_unsigned(141,8) ,
40050	 => std_logic_vector(to_unsigned(149,8) ,
40051	 => std_logic_vector(to_unsigned(154,8) ,
40052	 => std_logic_vector(to_unsigned(157,8) ,
40053	 => std_logic_vector(to_unsigned(161,8) ,
40054	 => std_logic_vector(to_unsigned(159,8) ,
40055	 => std_logic_vector(to_unsigned(156,8) ,
40056	 => std_logic_vector(to_unsigned(157,8) ,
40057	 => std_logic_vector(to_unsigned(161,8) ,
40058	 => std_logic_vector(to_unsigned(161,8) ,
40059	 => std_logic_vector(to_unsigned(157,8) ,
40060	 => std_logic_vector(to_unsigned(136,8) ,
40061	 => std_logic_vector(to_unsigned(10,8) ,
40062	 => std_logic_vector(to_unsigned(5,8) ,
40063	 => std_logic_vector(to_unsigned(18,8) ,
40064	 => std_logic_vector(to_unsigned(15,8) ,
40065	 => std_logic_vector(to_unsigned(4,8) ,
40066	 => std_logic_vector(to_unsigned(9,8) ,
40067	 => std_logic_vector(to_unsigned(121,8) ,
40068	 => std_logic_vector(to_unsigned(144,8) ,
40069	 => std_logic_vector(to_unsigned(138,8) ,
40070	 => std_logic_vector(to_unsigned(125,8) ,
40071	 => std_logic_vector(to_unsigned(109,8) ,
40072	 => std_logic_vector(to_unsigned(124,8) ,
40073	 => std_logic_vector(to_unsigned(133,8) ,
40074	 => std_logic_vector(to_unsigned(116,8) ,
40075	 => std_logic_vector(to_unsigned(118,8) ,
40076	 => std_logic_vector(to_unsigned(133,8) ,
40077	 => std_logic_vector(to_unsigned(133,8) ,
40078	 => std_logic_vector(to_unsigned(62,8) ,
40079	 => std_logic_vector(to_unsigned(41,8) ,
40080	 => std_logic_vector(to_unsigned(34,8) ,
40081	 => std_logic_vector(to_unsigned(4,8) ,
40082	 => std_logic_vector(to_unsigned(1,8) ,
40083	 => std_logic_vector(to_unsigned(0,8) ,
40084	 => std_logic_vector(to_unsigned(28,8) ,
40085	 => std_logic_vector(to_unsigned(86,8) ,
40086	 => std_logic_vector(to_unsigned(101,8) ,
40087	 => std_logic_vector(to_unsigned(144,8) ,
40088	 => std_logic_vector(to_unsigned(159,8) ,
40089	 => std_logic_vector(to_unsigned(151,8) ,
40090	 => std_logic_vector(to_unsigned(127,8) ,
40091	 => std_logic_vector(to_unsigned(128,8) ,
40092	 => std_logic_vector(to_unsigned(18,8) ,
40093	 => std_logic_vector(to_unsigned(4,8) ,
40094	 => std_logic_vector(to_unsigned(13,8) ,
40095	 => std_logic_vector(to_unsigned(13,8) ,
40096	 => std_logic_vector(to_unsigned(7,8) ,
40097	 => std_logic_vector(to_unsigned(6,8) ,
40098	 => std_logic_vector(to_unsigned(6,8) ,
40099	 => std_logic_vector(to_unsigned(3,8) ,
40100	 => std_logic_vector(to_unsigned(3,8) ,
40101	 => std_logic_vector(to_unsigned(3,8) ,
40102	 => std_logic_vector(to_unsigned(4,8) ,
40103	 => std_logic_vector(to_unsigned(3,8) ,
40104	 => std_logic_vector(to_unsigned(29,8) ,
40105	 => std_logic_vector(to_unsigned(41,8) ,
40106	 => std_logic_vector(to_unsigned(36,8) ,
40107	 => std_logic_vector(to_unsigned(24,8) ,
40108	 => std_logic_vector(to_unsigned(4,8) ,
40109	 => std_logic_vector(to_unsigned(0,8) ,
40110	 => std_logic_vector(to_unsigned(0,8) ,
40111	 => std_logic_vector(to_unsigned(0,8) ,
40112	 => std_logic_vector(to_unsigned(0,8) ,
40113	 => std_logic_vector(to_unsigned(0,8) ,
40114	 => std_logic_vector(to_unsigned(0,8) ,
40115	 => std_logic_vector(to_unsigned(0,8) ,
40116	 => std_logic_vector(to_unsigned(17,8) ,
40117	 => std_logic_vector(to_unsigned(109,8) ,
40118	 => std_logic_vector(to_unsigned(47,8) ,
40119	 => std_logic_vector(to_unsigned(22,8) ,
40120	 => std_logic_vector(to_unsigned(14,8) ,
40121	 => std_logic_vector(to_unsigned(3,8) ,
40122	 => std_logic_vector(to_unsigned(4,8) ,
40123	 => std_logic_vector(to_unsigned(6,8) ,
40124	 => std_logic_vector(to_unsigned(6,8) ,
40125	 => std_logic_vector(to_unsigned(4,8) ,
40126	 => std_logic_vector(to_unsigned(2,8) ,
40127	 => std_logic_vector(to_unsigned(4,8) ,
40128	 => std_logic_vector(to_unsigned(5,8) ,
40129	 => std_logic_vector(to_unsigned(2,8) ,
40130	 => std_logic_vector(to_unsigned(0,8) ,
40131	 => std_logic_vector(to_unsigned(0,8) ,
40132	 => std_logic_vector(to_unsigned(1,8) ,
40133	 => std_logic_vector(to_unsigned(1,8) ,
40134	 => std_logic_vector(to_unsigned(0,8) ,
40135	 => std_logic_vector(to_unsigned(1,8) ,
40136	 => std_logic_vector(to_unsigned(1,8) ,
40137	 => std_logic_vector(to_unsigned(0,8) ,
40138	 => std_logic_vector(to_unsigned(0,8) ,
40139	 => std_logic_vector(to_unsigned(1,8) ,
40140	 => std_logic_vector(to_unsigned(10,8) ,
40141	 => std_logic_vector(to_unsigned(8,8) ,
40142	 => std_logic_vector(to_unsigned(2,8) ,
40143	 => std_logic_vector(to_unsigned(2,8) ,
40144	 => std_logic_vector(to_unsigned(1,8) ,
40145	 => std_logic_vector(to_unsigned(0,8) ,
40146	 => std_logic_vector(to_unsigned(1,8) ,
40147	 => std_logic_vector(to_unsigned(2,8) ,
40148	 => std_logic_vector(to_unsigned(2,8) ,
40149	 => std_logic_vector(to_unsigned(3,8) ,
40150	 => std_logic_vector(to_unsigned(2,8) ,
40151	 => std_logic_vector(to_unsigned(2,8) ,
40152	 => std_logic_vector(to_unsigned(8,8) ,
40153	 => std_logic_vector(to_unsigned(9,8) ,
40154	 => std_logic_vector(to_unsigned(7,8) ,
40155	 => std_logic_vector(to_unsigned(4,8) ,
40156	 => std_logic_vector(to_unsigned(1,8) ,
40157	 => std_logic_vector(to_unsigned(1,8) ,
40158	 => std_logic_vector(to_unsigned(20,8) ,
40159	 => std_logic_vector(to_unsigned(10,8) ,
40160	 => std_logic_vector(to_unsigned(4,8) ,
40161	 => std_logic_vector(to_unsigned(8,8) ,
40162	 => std_logic_vector(to_unsigned(9,8) ,
40163	 => std_logic_vector(to_unsigned(7,8) ,
40164	 => std_logic_vector(to_unsigned(5,8) ,
40165	 => std_logic_vector(to_unsigned(3,8) ,
40166	 => std_logic_vector(to_unsigned(2,8) ,
40167	 => std_logic_vector(to_unsigned(1,8) ,
40168	 => std_logic_vector(to_unsigned(0,8) ,
40169	 => std_logic_vector(to_unsigned(0,8) ,
40170	 => std_logic_vector(to_unsigned(1,8) ,
40171	 => std_logic_vector(to_unsigned(1,8) ,
40172	 => std_logic_vector(to_unsigned(1,8) ,
40173	 => std_logic_vector(to_unsigned(1,8) ,
40174	 => std_logic_vector(to_unsigned(1,8) ,
40175	 => std_logic_vector(to_unsigned(1,8) ,
40176	 => std_logic_vector(to_unsigned(2,8) ,
40177	 => std_logic_vector(to_unsigned(5,8) ,
40178	 => std_logic_vector(to_unsigned(4,8) ,
40179	 => std_logic_vector(to_unsigned(3,8) ,
40180	 => std_logic_vector(to_unsigned(3,8) ,
40181	 => std_logic_vector(to_unsigned(1,8) ,
40182	 => std_logic_vector(to_unsigned(1,8) ,
40183	 => std_logic_vector(to_unsigned(3,8) ,
40184	 => std_logic_vector(to_unsigned(3,8) ,
40185	 => std_logic_vector(to_unsigned(3,8) ,
40186	 => std_logic_vector(to_unsigned(3,8) ,
40187	 => std_logic_vector(to_unsigned(3,8) ,
40188	 => std_logic_vector(to_unsigned(2,8) ,
40189	 => std_logic_vector(to_unsigned(1,8) ,
40190	 => std_logic_vector(to_unsigned(3,8) ,
40191	 => std_logic_vector(to_unsigned(3,8) ,
40192	 => std_logic_vector(to_unsigned(1,8) ,
40193	 => std_logic_vector(to_unsigned(0,8) ,
40194	 => std_logic_vector(to_unsigned(0,8) ,
40195	 => std_logic_vector(to_unsigned(0,8) ,
40196	 => std_logic_vector(to_unsigned(1,8) ,
40197	 => std_logic_vector(to_unsigned(1,8) ,
40198	 => std_logic_vector(to_unsigned(1,8) ,
40199	 => std_logic_vector(to_unsigned(1,8) ,
40200	 => std_logic_vector(to_unsigned(2,8) ,
40201	 => std_logic_vector(to_unsigned(1,8) ,
40202	 => std_logic_vector(to_unsigned(1,8) ,
40203	 => std_logic_vector(to_unsigned(2,8) ,
40204	 => std_logic_vector(to_unsigned(2,8) ,
40205	 => std_logic_vector(to_unsigned(2,8) ,
40206	 => std_logic_vector(to_unsigned(1,8) ,
40207	 => std_logic_vector(to_unsigned(3,8) ,
40208	 => std_logic_vector(to_unsigned(4,8) ,
40209	 => std_logic_vector(to_unsigned(6,8) ,
40210	 => std_logic_vector(to_unsigned(4,8) ,
40211	 => std_logic_vector(to_unsigned(6,8) ,
40212	 => std_logic_vector(to_unsigned(4,8) ,
40213	 => std_logic_vector(to_unsigned(1,8) ,
40214	 => std_logic_vector(to_unsigned(51,8) ,
40215	 => std_logic_vector(to_unsigned(133,8) ,
40216	 => std_logic_vector(to_unsigned(103,8) ,
40217	 => std_logic_vector(to_unsigned(57,8) ,
40218	 => std_logic_vector(to_unsigned(47,8) ,
40219	 => std_logic_vector(to_unsigned(31,8) ,
40220	 => std_logic_vector(to_unsigned(11,8) ,
40221	 => std_logic_vector(to_unsigned(0,8) ,
40222	 => std_logic_vector(to_unsigned(0,8) ,
40223	 => std_logic_vector(to_unsigned(0,8) ,
40224	 => std_logic_vector(to_unsigned(1,8) ,
40225	 => std_logic_vector(to_unsigned(2,8) ,
40226	 => std_logic_vector(to_unsigned(3,8) ,
40227	 => std_logic_vector(to_unsigned(3,8) ,
40228	 => std_logic_vector(to_unsigned(1,8) ,
40229	 => std_logic_vector(to_unsigned(4,8) ,
40230	 => std_logic_vector(to_unsigned(61,8) ,
40231	 => std_logic_vector(to_unsigned(79,8) ,
40232	 => std_logic_vector(to_unsigned(85,8) ,
40233	 => std_logic_vector(to_unsigned(124,8) ,
40234	 => std_logic_vector(to_unsigned(128,8) ,
40235	 => std_logic_vector(to_unsigned(62,8) ,
40236	 => std_logic_vector(to_unsigned(10,8) ,
40237	 => std_logic_vector(to_unsigned(2,8) ,
40238	 => std_logic_vector(to_unsigned(1,8) ,
40239	 => std_logic_vector(to_unsigned(4,8) ,
40240	 => std_logic_vector(to_unsigned(5,8) ,
40241	 => std_logic_vector(to_unsigned(4,8) ,
40242	 => std_logic_vector(to_unsigned(2,8) ,
40243	 => std_logic_vector(to_unsigned(0,8) ,
40244	 => std_logic_vector(to_unsigned(1,8) ,
40245	 => std_logic_vector(to_unsigned(2,8) ,
40246	 => std_logic_vector(to_unsigned(2,8) ,
40247	 => std_logic_vector(to_unsigned(11,8) ,
40248	 => std_logic_vector(to_unsigned(20,8) ,
40249	 => std_logic_vector(to_unsigned(5,8) ,
40250	 => std_logic_vector(to_unsigned(1,8) ,
40251	 => std_logic_vector(to_unsigned(2,8) ,
40252	 => std_logic_vector(to_unsigned(4,8) ,
40253	 => std_logic_vector(to_unsigned(3,8) ,
40254	 => std_logic_vector(to_unsigned(2,8) ,
40255	 => std_logic_vector(to_unsigned(2,8) ,
40256	 => std_logic_vector(to_unsigned(3,8) ,
40257	 => std_logic_vector(to_unsigned(2,8) ,
40258	 => std_logic_vector(to_unsigned(2,8) ,
40259	 => std_logic_vector(to_unsigned(5,8) ,
40260	 => std_logic_vector(to_unsigned(6,8) ,
40261	 => std_logic_vector(to_unsigned(2,8) ,
40262	 => std_logic_vector(to_unsigned(2,8) ,
40263	 => std_logic_vector(to_unsigned(6,8) ,
40264	 => std_logic_vector(to_unsigned(10,8) ,
40265	 => std_logic_vector(to_unsigned(13,8) ,
40266	 => std_logic_vector(to_unsigned(15,8) ,
40267	 => std_logic_vector(to_unsigned(25,8) ,
40268	 => std_logic_vector(to_unsigned(10,8) ,
40269	 => std_logic_vector(to_unsigned(9,8) ,
40270	 => std_logic_vector(to_unsigned(35,8) ,
40271	 => std_logic_vector(to_unsigned(99,8) ,
40272	 => std_logic_vector(to_unsigned(99,8) ,
40273	 => std_logic_vector(to_unsigned(60,8) ,
40274	 => std_logic_vector(to_unsigned(46,8) ,
40275	 => std_logic_vector(to_unsigned(30,8) ,
40276	 => std_logic_vector(to_unsigned(1,8) ,
40277	 => std_logic_vector(to_unsigned(1,8) ,
40278	 => std_logic_vector(to_unsigned(2,8) ,
40279	 => std_logic_vector(to_unsigned(1,8) ,
40280	 => std_logic_vector(to_unsigned(1,8) ,
40281	 => std_logic_vector(to_unsigned(2,8) ,
40282	 => std_logic_vector(to_unsigned(2,8) ,
40283	 => std_logic_vector(to_unsigned(3,8) ,
40284	 => std_logic_vector(to_unsigned(1,8) ,
40285	 => std_logic_vector(to_unsigned(2,8) ,
40286	 => std_logic_vector(to_unsigned(6,8) ,
40287	 => std_logic_vector(to_unsigned(6,8) ,
40288	 => std_logic_vector(to_unsigned(12,8) ,
40289	 => std_logic_vector(to_unsigned(11,8) ,
40290	 => std_logic_vector(to_unsigned(8,8) ,
40291	 => std_logic_vector(to_unsigned(8,8) ,
40292	 => std_logic_vector(to_unsigned(10,8) ,
40293	 => std_logic_vector(to_unsigned(11,8) ,
40294	 => std_logic_vector(to_unsigned(13,8) ,
40295	 => std_logic_vector(to_unsigned(5,8) ,
40296	 => std_logic_vector(to_unsigned(0,8) ,
40297	 => std_logic_vector(to_unsigned(0,8) ,
40298	 => std_logic_vector(to_unsigned(0,8) ,
40299	 => std_logic_vector(to_unsigned(1,8) ,
40300	 => std_logic_vector(to_unsigned(0,8) ,
40301	 => std_logic_vector(to_unsigned(1,8) ,
40302	 => std_logic_vector(to_unsigned(1,8) ,
40303	 => std_logic_vector(to_unsigned(0,8) ,
40304	 => std_logic_vector(to_unsigned(1,8) ,
40305	 => std_logic_vector(to_unsigned(0,8) ,
40306	 => std_logic_vector(to_unsigned(0,8) ,
40307	 => std_logic_vector(to_unsigned(0,8) ,
40308	 => std_logic_vector(to_unsigned(1,8) ,
40309	 => std_logic_vector(to_unsigned(1,8) ,
40310	 => std_logic_vector(to_unsigned(1,8) ,
40311	 => std_logic_vector(to_unsigned(1,8) ,
40312	 => std_logic_vector(to_unsigned(1,8) ,
40313	 => std_logic_vector(to_unsigned(1,8) ,
40314	 => std_logic_vector(to_unsigned(1,8) ,
40315	 => std_logic_vector(to_unsigned(1,8) ,
40316	 => std_logic_vector(to_unsigned(0,8) ,
40317	 => std_logic_vector(to_unsigned(1,8) ,
40318	 => std_logic_vector(to_unsigned(1,8) ,
40319	 => std_logic_vector(to_unsigned(1,8) ,
40320	 => std_logic_vector(to_unsigned(1,8) ,
40321	 => std_logic_vector(to_unsigned(136,8) ,
40322	 => std_logic_vector(to_unsigned(138,8) ,
40323	 => std_logic_vector(to_unsigned(131,8) ,
40324	 => std_logic_vector(to_unsigned(116,8) ,
40325	 => std_logic_vector(to_unsigned(114,8) ,
40326	 => std_logic_vector(to_unsigned(114,8) ,
40327	 => std_logic_vector(to_unsigned(109,8) ,
40328	 => std_logic_vector(to_unsigned(107,8) ,
40329	 => std_logic_vector(to_unsigned(105,8) ,
40330	 => std_logic_vector(to_unsigned(104,8) ,
40331	 => std_logic_vector(to_unsigned(104,8) ,
40332	 => std_logic_vector(to_unsigned(105,8) ,
40333	 => std_logic_vector(to_unsigned(115,8) ,
40334	 => std_logic_vector(to_unsigned(107,8) ,
40335	 => std_logic_vector(to_unsigned(112,8) ,
40336	 => std_logic_vector(to_unsigned(107,8) ,
40337	 => std_logic_vector(to_unsigned(57,8) ,
40338	 => std_logic_vector(to_unsigned(68,8) ,
40339	 => std_logic_vector(to_unsigned(115,8) ,
40340	 => std_logic_vector(to_unsigned(121,8) ,
40341	 => std_logic_vector(to_unsigned(109,8) ,
40342	 => std_logic_vector(to_unsigned(147,8) ,
40343	 => std_logic_vector(to_unsigned(156,8) ,
40344	 => std_logic_vector(to_unsigned(151,8) ,
40345	 => std_logic_vector(to_unsigned(152,8) ,
40346	 => std_logic_vector(to_unsigned(152,8) ,
40347	 => std_logic_vector(to_unsigned(146,8) ,
40348	 => std_logic_vector(to_unsigned(136,8) ,
40349	 => std_logic_vector(to_unsigned(131,8) ,
40350	 => std_logic_vector(to_unsigned(156,8) ,
40351	 => std_logic_vector(to_unsigned(142,8) ,
40352	 => std_logic_vector(to_unsigned(11,8) ,
40353	 => std_logic_vector(to_unsigned(2,8) ,
40354	 => std_logic_vector(to_unsigned(12,8) ,
40355	 => std_logic_vector(to_unsigned(7,8) ,
40356	 => std_logic_vector(to_unsigned(4,8) ,
40357	 => std_logic_vector(to_unsigned(2,8) ,
40358	 => std_logic_vector(to_unsigned(1,8) ,
40359	 => std_logic_vector(to_unsigned(1,8) ,
40360	 => std_logic_vector(to_unsigned(1,8) ,
40361	 => std_logic_vector(to_unsigned(33,8) ,
40362	 => std_logic_vector(to_unsigned(171,8) ,
40363	 => std_logic_vector(to_unsigned(157,8) ,
40364	 => std_logic_vector(to_unsigned(161,8) ,
40365	 => std_logic_vector(to_unsigned(157,8) ,
40366	 => std_logic_vector(to_unsigned(156,8) ,
40367	 => std_logic_vector(to_unsigned(159,8) ,
40368	 => std_logic_vector(to_unsigned(152,8) ,
40369	 => std_logic_vector(to_unsigned(147,8) ,
40370	 => std_logic_vector(to_unsigned(147,8) ,
40371	 => std_logic_vector(to_unsigned(154,8) ,
40372	 => std_logic_vector(to_unsigned(157,8) ,
40373	 => std_logic_vector(to_unsigned(159,8) ,
40374	 => std_logic_vector(to_unsigned(163,8) ,
40375	 => std_logic_vector(to_unsigned(159,8) ,
40376	 => std_logic_vector(to_unsigned(157,8) ,
40377	 => std_logic_vector(to_unsigned(159,8) ,
40378	 => std_logic_vector(to_unsigned(156,8) ,
40379	 => std_logic_vector(to_unsigned(157,8) ,
40380	 => std_logic_vector(to_unsigned(163,8) ,
40381	 => std_logic_vector(to_unsigned(42,8) ,
40382	 => std_logic_vector(to_unsigned(28,8) ,
40383	 => std_logic_vector(to_unsigned(59,8) ,
40384	 => std_logic_vector(to_unsigned(26,8) ,
40385	 => std_logic_vector(to_unsigned(4,8) ,
40386	 => std_logic_vector(to_unsigned(30,8) ,
40387	 => std_logic_vector(to_unsigned(133,8) ,
40388	 => std_logic_vector(to_unsigned(116,8) ,
40389	 => std_logic_vector(to_unsigned(116,8) ,
40390	 => std_logic_vector(to_unsigned(121,8) ,
40391	 => std_logic_vector(to_unsigned(116,8) ,
40392	 => std_logic_vector(to_unsigned(112,8) ,
40393	 => std_logic_vector(to_unsigned(108,8) ,
40394	 => std_logic_vector(to_unsigned(112,8) ,
40395	 => std_logic_vector(to_unsigned(121,8) ,
40396	 => std_logic_vector(to_unsigned(111,8) ,
40397	 => std_logic_vector(to_unsigned(121,8) ,
40398	 => std_logic_vector(to_unsigned(58,8) ,
40399	 => std_logic_vector(to_unsigned(5,8) ,
40400	 => std_logic_vector(to_unsigned(4,8) ,
40401	 => std_logic_vector(to_unsigned(3,8) ,
40402	 => std_logic_vector(to_unsigned(2,8) ,
40403	 => std_logic_vector(to_unsigned(0,8) ,
40404	 => std_logic_vector(to_unsigned(22,8) ,
40405	 => std_logic_vector(to_unsigned(177,8) ,
40406	 => std_logic_vector(to_unsigned(130,8) ,
40407	 => std_logic_vector(to_unsigned(103,8) ,
40408	 => std_logic_vector(to_unsigned(111,8) ,
40409	 => std_logic_vector(to_unsigned(114,8) ,
40410	 => std_logic_vector(to_unsigned(105,8) ,
40411	 => std_logic_vector(to_unsigned(136,8) ,
40412	 => std_logic_vector(to_unsigned(34,8) ,
40413	 => std_logic_vector(to_unsigned(1,8) ,
40414	 => std_logic_vector(to_unsigned(5,8) ,
40415	 => std_logic_vector(to_unsigned(6,8) ,
40416	 => std_logic_vector(to_unsigned(4,8) ,
40417	 => std_logic_vector(to_unsigned(5,8) ,
40418	 => std_logic_vector(to_unsigned(5,8) ,
40419	 => std_logic_vector(to_unsigned(5,8) ,
40420	 => std_logic_vector(to_unsigned(14,8) ,
40421	 => std_logic_vector(to_unsigned(48,8) ,
40422	 => std_logic_vector(to_unsigned(104,8) ,
40423	 => std_logic_vector(to_unsigned(64,8) ,
40424	 => std_logic_vector(to_unsigned(29,8) ,
40425	 => std_logic_vector(to_unsigned(34,8) ,
40426	 => std_logic_vector(to_unsigned(27,8) ,
40427	 => std_logic_vector(to_unsigned(15,8) ,
40428	 => std_logic_vector(to_unsigned(3,8) ,
40429	 => std_logic_vector(to_unsigned(4,8) ,
40430	 => std_logic_vector(to_unsigned(13,8) ,
40431	 => std_logic_vector(to_unsigned(6,8) ,
40432	 => std_logic_vector(to_unsigned(4,8) ,
40433	 => std_logic_vector(to_unsigned(2,8) ,
40434	 => std_logic_vector(to_unsigned(1,8) ,
40435	 => std_logic_vector(to_unsigned(0,8) ,
40436	 => std_logic_vector(to_unsigned(1,8) ,
40437	 => std_logic_vector(to_unsigned(13,8) ,
40438	 => std_logic_vector(to_unsigned(3,8) ,
40439	 => std_logic_vector(to_unsigned(0,8) ,
40440	 => std_logic_vector(to_unsigned(0,8) ,
40441	 => std_logic_vector(to_unsigned(0,8) ,
40442	 => std_logic_vector(to_unsigned(1,8) ,
40443	 => std_logic_vector(to_unsigned(4,8) ,
40444	 => std_logic_vector(to_unsigned(5,8) ,
40445	 => std_logic_vector(to_unsigned(3,8) ,
40446	 => std_logic_vector(to_unsigned(3,8) ,
40447	 => std_logic_vector(to_unsigned(2,8) ,
40448	 => std_logic_vector(to_unsigned(3,8) ,
40449	 => std_logic_vector(to_unsigned(1,8) ,
40450	 => std_logic_vector(to_unsigned(1,8) ,
40451	 => std_logic_vector(to_unsigned(0,8) ,
40452	 => std_logic_vector(to_unsigned(0,8) ,
40453	 => std_logic_vector(to_unsigned(0,8) ,
40454	 => std_logic_vector(to_unsigned(0,8) ,
40455	 => std_logic_vector(to_unsigned(0,8) ,
40456	 => std_logic_vector(to_unsigned(1,8) ,
40457	 => std_logic_vector(to_unsigned(1,8) ,
40458	 => std_logic_vector(to_unsigned(1,8) ,
40459	 => std_logic_vector(to_unsigned(6,8) ,
40460	 => std_logic_vector(to_unsigned(17,8) ,
40461	 => std_logic_vector(to_unsigned(7,8) ,
40462	 => std_logic_vector(to_unsigned(4,8) ,
40463	 => std_logic_vector(to_unsigned(2,8) ,
40464	 => std_logic_vector(to_unsigned(1,8) ,
40465	 => std_logic_vector(to_unsigned(0,8) ,
40466	 => std_logic_vector(to_unsigned(1,8) ,
40467	 => std_logic_vector(to_unsigned(1,8) ,
40468	 => std_logic_vector(to_unsigned(2,8) ,
40469	 => std_logic_vector(to_unsigned(2,8) ,
40470	 => std_logic_vector(to_unsigned(2,8) ,
40471	 => std_logic_vector(to_unsigned(3,8) ,
40472	 => std_logic_vector(to_unsigned(8,8) ,
40473	 => std_logic_vector(to_unsigned(7,8) ,
40474	 => std_logic_vector(to_unsigned(5,8) ,
40475	 => std_logic_vector(to_unsigned(4,8) ,
40476	 => std_logic_vector(to_unsigned(1,8) ,
40477	 => std_logic_vector(to_unsigned(1,8) ,
40478	 => std_logic_vector(to_unsigned(10,8) ,
40479	 => std_logic_vector(to_unsigned(8,8) ,
40480	 => std_logic_vector(to_unsigned(5,8) ,
40481	 => std_logic_vector(to_unsigned(4,8) ,
40482	 => std_logic_vector(to_unsigned(2,8) ,
40483	 => std_logic_vector(to_unsigned(1,8) ,
40484	 => std_logic_vector(to_unsigned(4,8) ,
40485	 => std_logic_vector(to_unsigned(3,8) ,
40486	 => std_logic_vector(to_unsigned(1,8) ,
40487	 => std_logic_vector(to_unsigned(1,8) ,
40488	 => std_logic_vector(to_unsigned(1,8) ,
40489	 => std_logic_vector(to_unsigned(0,8) ,
40490	 => std_logic_vector(to_unsigned(0,8) ,
40491	 => std_logic_vector(to_unsigned(1,8) ,
40492	 => std_logic_vector(to_unsigned(1,8) ,
40493	 => std_logic_vector(to_unsigned(2,8) ,
40494	 => std_logic_vector(to_unsigned(1,8) ,
40495	 => std_logic_vector(to_unsigned(0,8) ,
40496	 => std_logic_vector(to_unsigned(0,8) ,
40497	 => std_logic_vector(to_unsigned(2,8) ,
40498	 => std_logic_vector(to_unsigned(4,8) ,
40499	 => std_logic_vector(to_unsigned(4,8) ,
40500	 => std_logic_vector(to_unsigned(1,8) ,
40501	 => std_logic_vector(to_unsigned(0,8) ,
40502	 => std_logic_vector(to_unsigned(2,8) ,
40503	 => std_logic_vector(to_unsigned(6,8) ,
40504	 => std_logic_vector(to_unsigned(3,8) ,
40505	 => std_logic_vector(to_unsigned(1,8) ,
40506	 => std_logic_vector(to_unsigned(2,8) ,
40507	 => std_logic_vector(to_unsigned(2,8) ,
40508	 => std_logic_vector(to_unsigned(2,8) ,
40509	 => std_logic_vector(to_unsigned(2,8) ,
40510	 => std_logic_vector(to_unsigned(2,8) ,
40511	 => std_logic_vector(to_unsigned(1,8) ,
40512	 => std_logic_vector(to_unsigned(1,8) ,
40513	 => std_logic_vector(to_unsigned(0,8) ,
40514	 => std_logic_vector(to_unsigned(0,8) ,
40515	 => std_logic_vector(to_unsigned(0,8) ,
40516	 => std_logic_vector(to_unsigned(1,8) ,
40517	 => std_logic_vector(to_unsigned(1,8) ,
40518	 => std_logic_vector(to_unsigned(1,8) ,
40519	 => std_logic_vector(to_unsigned(2,8) ,
40520	 => std_logic_vector(to_unsigned(1,8) ,
40521	 => std_logic_vector(to_unsigned(1,8) ,
40522	 => std_logic_vector(to_unsigned(1,8) ,
40523	 => std_logic_vector(to_unsigned(1,8) ,
40524	 => std_logic_vector(to_unsigned(1,8) ,
40525	 => std_logic_vector(to_unsigned(1,8) ,
40526	 => std_logic_vector(to_unsigned(1,8) ,
40527	 => std_logic_vector(to_unsigned(3,8) ,
40528	 => std_logic_vector(to_unsigned(3,8) ,
40529	 => std_logic_vector(to_unsigned(4,8) ,
40530	 => std_logic_vector(to_unsigned(4,8) ,
40531	 => std_logic_vector(to_unsigned(6,8) ,
40532	 => std_logic_vector(to_unsigned(3,8) ,
40533	 => std_logic_vector(to_unsigned(2,8) ,
40534	 => std_logic_vector(to_unsigned(47,8) ,
40535	 => std_logic_vector(to_unsigned(115,8) ,
40536	 => std_logic_vector(to_unsigned(93,8) ,
40537	 => std_logic_vector(to_unsigned(55,8) ,
40538	 => std_logic_vector(to_unsigned(54,8) ,
40539	 => std_logic_vector(to_unsigned(37,8) ,
40540	 => std_logic_vector(to_unsigned(5,8) ,
40541	 => std_logic_vector(to_unsigned(0,8) ,
40542	 => std_logic_vector(to_unsigned(0,8) ,
40543	 => std_logic_vector(to_unsigned(0,8) ,
40544	 => std_logic_vector(to_unsigned(1,8) ,
40545	 => std_logic_vector(to_unsigned(2,8) ,
40546	 => std_logic_vector(to_unsigned(2,8) ,
40547	 => std_logic_vector(to_unsigned(2,8) ,
40548	 => std_logic_vector(to_unsigned(2,8) ,
40549	 => std_logic_vector(to_unsigned(2,8) ,
40550	 => std_logic_vector(to_unsigned(56,8) ,
40551	 => std_logic_vector(to_unsigned(84,8) ,
40552	 => std_logic_vector(to_unsigned(54,8) ,
40553	 => std_logic_vector(to_unsigned(99,8) ,
40554	 => std_logic_vector(to_unsigned(119,8) ,
40555	 => std_logic_vector(to_unsigned(74,8) ,
40556	 => std_logic_vector(to_unsigned(10,8) ,
40557	 => std_logic_vector(to_unsigned(0,8) ,
40558	 => std_logic_vector(to_unsigned(1,8) ,
40559	 => std_logic_vector(to_unsigned(4,8) ,
40560	 => std_logic_vector(to_unsigned(4,8) ,
40561	 => std_logic_vector(to_unsigned(5,8) ,
40562	 => std_logic_vector(to_unsigned(4,8) ,
40563	 => std_logic_vector(to_unsigned(1,8) ,
40564	 => std_logic_vector(to_unsigned(1,8) ,
40565	 => std_logic_vector(to_unsigned(1,8) ,
40566	 => std_logic_vector(to_unsigned(1,8) ,
40567	 => std_logic_vector(to_unsigned(10,8) ,
40568	 => std_logic_vector(to_unsigned(21,8) ,
40569	 => std_logic_vector(to_unsigned(11,8) ,
40570	 => std_logic_vector(to_unsigned(1,8) ,
40571	 => std_logic_vector(to_unsigned(2,8) ,
40572	 => std_logic_vector(to_unsigned(3,8) ,
40573	 => std_logic_vector(to_unsigned(4,8) ,
40574	 => std_logic_vector(to_unsigned(2,8) ,
40575	 => std_logic_vector(to_unsigned(2,8) ,
40576	 => std_logic_vector(to_unsigned(3,8) ,
40577	 => std_logic_vector(to_unsigned(2,8) ,
40578	 => std_logic_vector(to_unsigned(2,8) ,
40579	 => std_logic_vector(to_unsigned(4,8) ,
40580	 => std_logic_vector(to_unsigned(6,8) ,
40581	 => std_logic_vector(to_unsigned(2,8) ,
40582	 => std_logic_vector(to_unsigned(1,8) ,
40583	 => std_logic_vector(to_unsigned(3,8) ,
40584	 => std_logic_vector(to_unsigned(7,8) ,
40585	 => std_logic_vector(to_unsigned(11,8) ,
40586	 => std_logic_vector(to_unsigned(18,8) ,
40587	 => std_logic_vector(to_unsigned(34,8) ,
40588	 => std_logic_vector(to_unsigned(12,8) ,
40589	 => std_logic_vector(to_unsigned(6,8) ,
40590	 => std_logic_vector(to_unsigned(14,8) ,
40591	 => std_logic_vector(to_unsigned(15,8) ,
40592	 => std_logic_vector(to_unsigned(30,8) ,
40593	 => std_logic_vector(to_unsigned(54,8) ,
40594	 => std_logic_vector(to_unsigned(13,8) ,
40595	 => std_logic_vector(to_unsigned(5,8) ,
40596	 => std_logic_vector(to_unsigned(2,8) ,
40597	 => std_logic_vector(to_unsigned(1,8) ,
40598	 => std_logic_vector(to_unsigned(1,8) ,
40599	 => std_logic_vector(to_unsigned(1,8) ,
40600	 => std_logic_vector(to_unsigned(2,8) ,
40601	 => std_logic_vector(to_unsigned(3,8) ,
40602	 => std_logic_vector(to_unsigned(2,8) ,
40603	 => std_logic_vector(to_unsigned(2,8) ,
40604	 => std_logic_vector(to_unsigned(2,8) ,
40605	 => std_logic_vector(to_unsigned(6,8) ,
40606	 => std_logic_vector(to_unsigned(5,8) ,
40607	 => std_logic_vector(to_unsigned(6,8) ,
40608	 => std_logic_vector(to_unsigned(10,8) ,
40609	 => std_logic_vector(to_unsigned(6,8) ,
40610	 => std_logic_vector(to_unsigned(5,8) ,
40611	 => std_logic_vector(to_unsigned(7,8) ,
40612	 => std_logic_vector(to_unsigned(7,8) ,
40613	 => std_logic_vector(to_unsigned(9,8) ,
40614	 => std_logic_vector(to_unsigned(18,8) ,
40615	 => std_logic_vector(to_unsigned(9,8) ,
40616	 => std_logic_vector(to_unsigned(0,8) ,
40617	 => std_logic_vector(to_unsigned(0,8) ,
40618	 => std_logic_vector(to_unsigned(0,8) ,
40619	 => std_logic_vector(to_unsigned(1,8) ,
40620	 => std_logic_vector(to_unsigned(1,8) ,
40621	 => std_logic_vector(to_unsigned(1,8) ,
40622	 => std_logic_vector(to_unsigned(1,8) ,
40623	 => std_logic_vector(to_unsigned(0,8) ,
40624	 => std_logic_vector(to_unsigned(1,8) ,
40625	 => std_logic_vector(to_unsigned(1,8) ,
40626	 => std_logic_vector(to_unsigned(1,8) ,
40627	 => std_logic_vector(to_unsigned(1,8) ,
40628	 => std_logic_vector(to_unsigned(1,8) ,
40629	 => std_logic_vector(to_unsigned(1,8) ,
40630	 => std_logic_vector(to_unsigned(1,8) ,
40631	 => std_logic_vector(to_unsigned(1,8) ,
40632	 => std_logic_vector(to_unsigned(1,8) ,
40633	 => std_logic_vector(to_unsigned(1,8) ,
40634	 => std_logic_vector(to_unsigned(1,8) ,
40635	 => std_logic_vector(to_unsigned(1,8) ,
40636	 => std_logic_vector(to_unsigned(1,8) ,
40637	 => std_logic_vector(to_unsigned(1,8) ,
40638	 => std_logic_vector(to_unsigned(1,8) ,
40639	 => std_logic_vector(to_unsigned(1,8) ,
40640	 => std_logic_vector(to_unsigned(1,8) ,
40641	 => std_logic_vector(to_unsigned(136,8) ,
40642	 => std_logic_vector(to_unsigned(131,8) ,
40643	 => std_logic_vector(to_unsigned(128,8) ,
40644	 => std_logic_vector(to_unsigned(116,8) ,
40645	 => std_logic_vector(to_unsigned(109,8) ,
40646	 => std_logic_vector(to_unsigned(109,8) ,
40647	 => std_logic_vector(to_unsigned(108,8) ,
40648	 => std_logic_vector(to_unsigned(96,8) ,
40649	 => std_logic_vector(to_unsigned(91,8) ,
40650	 => std_logic_vector(to_unsigned(93,8) ,
40651	 => std_logic_vector(to_unsigned(103,8) ,
40652	 => std_logic_vector(to_unsigned(112,8) ,
40653	 => std_logic_vector(to_unsigned(116,8) ,
40654	 => std_logic_vector(to_unsigned(105,8) ,
40655	 => std_logic_vector(to_unsigned(114,8) ,
40656	 => std_logic_vector(to_unsigned(130,8) ,
40657	 => std_logic_vector(to_unsigned(156,8) ,
40658	 => std_logic_vector(to_unsigned(170,8) ,
40659	 => std_logic_vector(to_unsigned(142,8) ,
40660	 => std_logic_vector(to_unsigned(111,8) ,
40661	 => std_logic_vector(to_unsigned(109,8) ,
40662	 => std_logic_vector(to_unsigned(134,8) ,
40663	 => std_logic_vector(to_unsigned(147,8) ,
40664	 => std_logic_vector(to_unsigned(142,8) ,
40665	 => std_logic_vector(to_unsigned(142,8) ,
40666	 => std_logic_vector(to_unsigned(151,8) ,
40667	 => std_logic_vector(to_unsigned(141,8) ,
40668	 => std_logic_vector(to_unsigned(130,8) ,
40669	 => std_logic_vector(to_unsigned(139,8) ,
40670	 => std_logic_vector(to_unsigned(154,8) ,
40671	 => std_logic_vector(to_unsigned(33,8) ,
40672	 => std_logic_vector(to_unsigned(2,8) ,
40673	 => std_logic_vector(to_unsigned(17,8) ,
40674	 => std_logic_vector(to_unsigned(14,8) ,
40675	 => std_logic_vector(to_unsigned(4,8) ,
40676	 => std_logic_vector(to_unsigned(2,8) ,
40677	 => std_logic_vector(to_unsigned(2,8) ,
40678	 => std_logic_vector(to_unsigned(2,8) ,
40679	 => std_logic_vector(to_unsigned(2,8) ,
40680	 => std_logic_vector(to_unsigned(1,8) ,
40681	 => std_logic_vector(to_unsigned(35,8) ,
40682	 => std_logic_vector(to_unsigned(179,8) ,
40683	 => std_logic_vector(to_unsigned(154,8) ,
40684	 => std_logic_vector(to_unsigned(157,8) ,
40685	 => std_logic_vector(to_unsigned(161,8) ,
40686	 => std_logic_vector(to_unsigned(161,8) ,
40687	 => std_logic_vector(to_unsigned(161,8) ,
40688	 => std_logic_vector(to_unsigned(161,8) ,
40689	 => std_logic_vector(to_unsigned(164,8) ,
40690	 => std_logic_vector(to_unsigned(161,8) ,
40691	 => std_logic_vector(to_unsigned(161,8) ,
40692	 => std_logic_vector(to_unsigned(156,8) ,
40693	 => std_logic_vector(to_unsigned(157,8) ,
40694	 => std_logic_vector(to_unsigned(157,8) ,
40695	 => std_logic_vector(to_unsigned(157,8) ,
40696	 => std_logic_vector(to_unsigned(161,8) ,
40697	 => std_logic_vector(to_unsigned(161,8) ,
40698	 => std_logic_vector(to_unsigned(161,8) ,
40699	 => std_logic_vector(to_unsigned(159,8) ,
40700	 => std_logic_vector(to_unsigned(166,8) ,
40701	 => std_logic_vector(to_unsigned(93,8) ,
40702	 => std_logic_vector(to_unsigned(9,8) ,
40703	 => std_logic_vector(to_unsigned(9,8) ,
40704	 => std_logic_vector(to_unsigned(5,8) ,
40705	 => std_logic_vector(to_unsigned(14,8) ,
40706	 => std_logic_vector(to_unsigned(124,8) ,
40707	 => std_logic_vector(to_unsigned(142,8) ,
40708	 => std_logic_vector(to_unsigned(118,8) ,
40709	 => std_logic_vector(to_unsigned(119,8) ,
40710	 => std_logic_vector(to_unsigned(118,8) ,
40711	 => std_logic_vector(to_unsigned(108,8) ,
40712	 => std_logic_vector(to_unsigned(104,8) ,
40713	 => std_logic_vector(to_unsigned(111,8) ,
40714	 => std_logic_vector(to_unsigned(122,8) ,
40715	 => std_logic_vector(to_unsigned(116,8) ,
40716	 => std_logic_vector(to_unsigned(111,8) ,
40717	 => std_logic_vector(to_unsigned(109,8) ,
40718	 => std_logic_vector(to_unsigned(25,8) ,
40719	 => std_logic_vector(to_unsigned(1,8) ,
40720	 => std_logic_vector(to_unsigned(4,8) ,
40721	 => std_logic_vector(to_unsigned(11,8) ,
40722	 => std_logic_vector(to_unsigned(2,8) ,
40723	 => std_logic_vector(to_unsigned(0,8) ,
40724	 => std_logic_vector(to_unsigned(1,8) ,
40725	 => std_logic_vector(to_unsigned(68,8) ,
40726	 => std_logic_vector(to_unsigned(151,8) ,
40727	 => std_logic_vector(to_unsigned(111,8) ,
40728	 => std_logic_vector(to_unsigned(105,8) ,
40729	 => std_logic_vector(to_unsigned(115,8) ,
40730	 => std_logic_vector(to_unsigned(103,8) ,
40731	 => std_logic_vector(to_unsigned(114,8) ,
40732	 => std_logic_vector(to_unsigned(69,8) ,
40733	 => std_logic_vector(to_unsigned(15,8) ,
40734	 => std_logic_vector(to_unsigned(32,8) ,
40735	 => std_logic_vector(to_unsigned(25,8) ,
40736	 => std_logic_vector(to_unsigned(51,8) ,
40737	 => std_logic_vector(to_unsigned(48,8) ,
40738	 => std_logic_vector(to_unsigned(20,8) ,
40739	 => std_logic_vector(to_unsigned(4,8) ,
40740	 => std_logic_vector(to_unsigned(20,8) ,
40741	 => std_logic_vector(to_unsigned(127,8) ,
40742	 => std_logic_vector(to_unsigned(151,8) ,
40743	 => std_logic_vector(to_unsigned(72,8) ,
40744	 => std_logic_vector(to_unsigned(3,8) ,
40745	 => std_logic_vector(to_unsigned(4,8) ,
40746	 => std_logic_vector(to_unsigned(3,8) ,
40747	 => std_logic_vector(to_unsigned(1,8) ,
40748	 => std_logic_vector(to_unsigned(0,8) ,
40749	 => std_logic_vector(to_unsigned(9,8) ,
40750	 => std_logic_vector(to_unsigned(111,8) ,
40751	 => std_logic_vector(to_unsigned(133,8) ,
40752	 => std_logic_vector(to_unsigned(81,8) ,
40753	 => std_logic_vector(to_unsigned(67,8) ,
40754	 => std_logic_vector(to_unsigned(63,8) ,
40755	 => std_logic_vector(to_unsigned(46,8) ,
40756	 => std_logic_vector(to_unsigned(34,8) ,
40757	 => std_logic_vector(to_unsigned(17,8) ,
40758	 => std_logic_vector(to_unsigned(12,8) ,
40759	 => std_logic_vector(to_unsigned(13,8) ,
40760	 => std_logic_vector(to_unsigned(9,8) ,
40761	 => std_logic_vector(to_unsigned(5,8) ,
40762	 => std_logic_vector(to_unsigned(3,8) ,
40763	 => std_logic_vector(to_unsigned(1,8) ,
40764	 => std_logic_vector(to_unsigned(1,8) ,
40765	 => std_logic_vector(to_unsigned(1,8) ,
40766	 => std_logic_vector(to_unsigned(4,8) ,
40767	 => std_logic_vector(to_unsigned(7,8) ,
40768	 => std_logic_vector(to_unsigned(4,8) ,
40769	 => std_logic_vector(to_unsigned(1,8) ,
40770	 => std_logic_vector(to_unsigned(0,8) ,
40771	 => std_logic_vector(to_unsigned(0,8) ,
40772	 => std_logic_vector(to_unsigned(0,8) ,
40773	 => std_logic_vector(to_unsigned(0,8) ,
40774	 => std_logic_vector(to_unsigned(0,8) ,
40775	 => std_logic_vector(to_unsigned(0,8) ,
40776	 => std_logic_vector(to_unsigned(1,8) ,
40777	 => std_logic_vector(to_unsigned(1,8) ,
40778	 => std_logic_vector(to_unsigned(2,8) ,
40779	 => std_logic_vector(to_unsigned(21,8) ,
40780	 => std_logic_vector(to_unsigned(20,8) ,
40781	 => std_logic_vector(to_unsigned(7,8) ,
40782	 => std_logic_vector(to_unsigned(3,8) ,
40783	 => std_logic_vector(to_unsigned(2,8) ,
40784	 => std_logic_vector(to_unsigned(1,8) ,
40785	 => std_logic_vector(to_unsigned(1,8) ,
40786	 => std_logic_vector(to_unsigned(1,8) ,
40787	 => std_logic_vector(to_unsigned(1,8) ,
40788	 => std_logic_vector(to_unsigned(3,8) ,
40789	 => std_logic_vector(to_unsigned(3,8) ,
40790	 => std_logic_vector(to_unsigned(3,8) ,
40791	 => std_logic_vector(to_unsigned(4,8) ,
40792	 => std_logic_vector(to_unsigned(4,8) ,
40793	 => std_logic_vector(to_unsigned(4,8) ,
40794	 => std_logic_vector(to_unsigned(3,8) ,
40795	 => std_logic_vector(to_unsigned(3,8) ,
40796	 => std_logic_vector(to_unsigned(1,8) ,
40797	 => std_logic_vector(to_unsigned(0,8) ,
40798	 => std_logic_vector(to_unsigned(0,8) ,
40799	 => std_logic_vector(to_unsigned(1,8) ,
40800	 => std_logic_vector(to_unsigned(1,8) ,
40801	 => std_logic_vector(to_unsigned(0,8) ,
40802	 => std_logic_vector(to_unsigned(0,8) ,
40803	 => std_logic_vector(to_unsigned(2,8) ,
40804	 => std_logic_vector(to_unsigned(9,8) ,
40805	 => std_logic_vector(to_unsigned(6,8) ,
40806	 => std_logic_vector(to_unsigned(2,8) ,
40807	 => std_logic_vector(to_unsigned(1,8) ,
40808	 => std_logic_vector(to_unsigned(2,8) ,
40809	 => std_logic_vector(to_unsigned(1,8) ,
40810	 => std_logic_vector(to_unsigned(1,8) ,
40811	 => std_logic_vector(to_unsigned(1,8) ,
40812	 => std_logic_vector(to_unsigned(1,8) ,
40813	 => std_logic_vector(to_unsigned(1,8) ,
40814	 => std_logic_vector(to_unsigned(1,8) ,
40815	 => std_logic_vector(to_unsigned(1,8) ,
40816	 => std_logic_vector(to_unsigned(1,8) ,
40817	 => std_logic_vector(to_unsigned(0,8) ,
40818	 => std_logic_vector(to_unsigned(1,8) ,
40819	 => std_logic_vector(to_unsigned(3,8) ,
40820	 => std_logic_vector(to_unsigned(0,8) ,
40821	 => std_logic_vector(to_unsigned(0,8) ,
40822	 => std_logic_vector(to_unsigned(3,8) ,
40823	 => std_logic_vector(to_unsigned(10,8) ,
40824	 => std_logic_vector(to_unsigned(6,8) ,
40825	 => std_logic_vector(to_unsigned(3,8) ,
40826	 => std_logic_vector(to_unsigned(2,8) ,
40827	 => std_logic_vector(to_unsigned(1,8) ,
40828	 => std_logic_vector(to_unsigned(2,8) ,
40829	 => std_logic_vector(to_unsigned(2,8) ,
40830	 => std_logic_vector(to_unsigned(1,8) ,
40831	 => std_logic_vector(to_unsigned(1,8) ,
40832	 => std_logic_vector(to_unsigned(0,8) ,
40833	 => std_logic_vector(to_unsigned(0,8) ,
40834	 => std_logic_vector(to_unsigned(0,8) ,
40835	 => std_logic_vector(to_unsigned(1,8) ,
40836	 => std_logic_vector(to_unsigned(1,8) ,
40837	 => std_logic_vector(to_unsigned(1,8) ,
40838	 => std_logic_vector(to_unsigned(1,8) ,
40839	 => std_logic_vector(to_unsigned(1,8) ,
40840	 => std_logic_vector(to_unsigned(1,8) ,
40841	 => std_logic_vector(to_unsigned(1,8) ,
40842	 => std_logic_vector(to_unsigned(1,8) ,
40843	 => std_logic_vector(to_unsigned(1,8) ,
40844	 => std_logic_vector(to_unsigned(2,8) ,
40845	 => std_logic_vector(to_unsigned(1,8) ,
40846	 => std_logic_vector(to_unsigned(2,8) ,
40847	 => std_logic_vector(to_unsigned(2,8) ,
40848	 => std_logic_vector(to_unsigned(2,8) ,
40849	 => std_logic_vector(to_unsigned(5,8) ,
40850	 => std_logic_vector(to_unsigned(6,8) ,
40851	 => std_logic_vector(to_unsigned(7,8) ,
40852	 => std_logic_vector(to_unsigned(2,8) ,
40853	 => std_logic_vector(to_unsigned(4,8) ,
40854	 => std_logic_vector(to_unsigned(57,8) ,
40855	 => std_logic_vector(to_unsigned(86,8) ,
40856	 => std_logic_vector(to_unsigned(86,8) ,
40857	 => std_logic_vector(to_unsigned(61,8) ,
40858	 => std_logic_vector(to_unsigned(62,8) ,
40859	 => std_logic_vector(to_unsigned(41,8) ,
40860	 => std_logic_vector(to_unsigned(6,8) ,
40861	 => std_logic_vector(to_unsigned(0,8) ,
40862	 => std_logic_vector(to_unsigned(0,8) ,
40863	 => std_logic_vector(to_unsigned(1,8) ,
40864	 => std_logic_vector(to_unsigned(1,8) ,
40865	 => std_logic_vector(to_unsigned(2,8) ,
40866	 => std_logic_vector(to_unsigned(2,8) ,
40867	 => std_logic_vector(to_unsigned(2,8) ,
40868	 => std_logic_vector(to_unsigned(2,8) ,
40869	 => std_logic_vector(to_unsigned(3,8) ,
40870	 => std_logic_vector(to_unsigned(54,8) ,
40871	 => std_logic_vector(to_unsigned(144,8) ,
40872	 => std_logic_vector(to_unsigned(114,8) ,
40873	 => std_logic_vector(to_unsigned(93,8) ,
40874	 => std_logic_vector(to_unsigned(112,8) ,
40875	 => std_logic_vector(to_unsigned(77,8) ,
40876	 => std_logic_vector(to_unsigned(12,8) ,
40877	 => std_logic_vector(to_unsigned(0,8) ,
40878	 => std_logic_vector(to_unsigned(1,8) ,
40879	 => std_logic_vector(to_unsigned(7,8) ,
40880	 => std_logic_vector(to_unsigned(6,8) ,
40881	 => std_logic_vector(to_unsigned(4,8) ,
40882	 => std_logic_vector(to_unsigned(5,8) ,
40883	 => std_logic_vector(to_unsigned(2,8) ,
40884	 => std_logic_vector(to_unsigned(1,8) ,
40885	 => std_logic_vector(to_unsigned(1,8) ,
40886	 => std_logic_vector(to_unsigned(1,8) ,
40887	 => std_logic_vector(to_unsigned(7,8) ,
40888	 => std_logic_vector(to_unsigned(13,8) ,
40889	 => std_logic_vector(to_unsigned(12,8) ,
40890	 => std_logic_vector(to_unsigned(2,8) ,
40891	 => std_logic_vector(to_unsigned(2,8) ,
40892	 => std_logic_vector(to_unsigned(3,8) ,
40893	 => std_logic_vector(to_unsigned(3,8) ,
40894	 => std_logic_vector(to_unsigned(2,8) ,
40895	 => std_logic_vector(to_unsigned(2,8) ,
40896	 => std_logic_vector(to_unsigned(2,8) ,
40897	 => std_logic_vector(to_unsigned(1,8) ,
40898	 => std_logic_vector(to_unsigned(2,8) ,
40899	 => std_logic_vector(to_unsigned(5,8) ,
40900	 => std_logic_vector(to_unsigned(6,8) ,
40901	 => std_logic_vector(to_unsigned(2,8) ,
40902	 => std_logic_vector(to_unsigned(1,8) ,
40903	 => std_logic_vector(to_unsigned(2,8) ,
40904	 => std_logic_vector(to_unsigned(5,8) ,
40905	 => std_logic_vector(to_unsigned(6,8) ,
40906	 => std_logic_vector(to_unsigned(19,8) ,
40907	 => std_logic_vector(to_unsigned(44,8) ,
40908	 => std_logic_vector(to_unsigned(25,8) ,
40909	 => std_logic_vector(to_unsigned(13,8) ,
40910	 => std_logic_vector(to_unsigned(8,8) ,
40911	 => std_logic_vector(to_unsigned(4,8) ,
40912	 => std_logic_vector(to_unsigned(15,8) ,
40913	 => std_logic_vector(to_unsigned(35,8) ,
40914	 => std_logic_vector(to_unsigned(12,8) ,
40915	 => std_logic_vector(to_unsigned(5,8) ,
40916	 => std_logic_vector(to_unsigned(1,8) ,
40917	 => std_logic_vector(to_unsigned(1,8) ,
40918	 => std_logic_vector(to_unsigned(2,8) ,
40919	 => std_logic_vector(to_unsigned(2,8) ,
40920	 => std_logic_vector(to_unsigned(3,8) ,
40921	 => std_logic_vector(to_unsigned(3,8) ,
40922	 => std_logic_vector(to_unsigned(2,8) ,
40923	 => std_logic_vector(to_unsigned(3,8) ,
40924	 => std_logic_vector(to_unsigned(7,8) ,
40925	 => std_logic_vector(to_unsigned(6,8) ,
40926	 => std_logic_vector(to_unsigned(5,8) ,
40927	 => std_logic_vector(to_unsigned(8,8) ,
40928	 => std_logic_vector(to_unsigned(8,8) ,
40929	 => std_logic_vector(to_unsigned(7,8) ,
40930	 => std_logic_vector(to_unsigned(5,8) ,
40931	 => std_logic_vector(to_unsigned(6,8) ,
40932	 => std_logic_vector(to_unsigned(3,8) ,
40933	 => std_logic_vector(to_unsigned(2,8) ,
40934	 => std_logic_vector(to_unsigned(7,8) ,
40935	 => std_logic_vector(to_unsigned(11,8) ,
40936	 => std_logic_vector(to_unsigned(1,8) ,
40937	 => std_logic_vector(to_unsigned(0,8) ,
40938	 => std_logic_vector(to_unsigned(1,8) ,
40939	 => std_logic_vector(to_unsigned(1,8) ,
40940	 => std_logic_vector(to_unsigned(1,8) ,
40941	 => std_logic_vector(to_unsigned(1,8) ,
40942	 => std_logic_vector(to_unsigned(1,8) ,
40943	 => std_logic_vector(to_unsigned(1,8) ,
40944	 => std_logic_vector(to_unsigned(1,8) ,
40945	 => std_logic_vector(to_unsigned(1,8) ,
40946	 => std_logic_vector(to_unsigned(1,8) ,
40947	 => std_logic_vector(to_unsigned(1,8) ,
40948	 => std_logic_vector(to_unsigned(1,8) ,
40949	 => std_logic_vector(to_unsigned(1,8) ,
40950	 => std_logic_vector(to_unsigned(1,8) ,
40951	 => std_logic_vector(to_unsigned(1,8) ,
40952	 => std_logic_vector(to_unsigned(1,8) ,
40953	 => std_logic_vector(to_unsigned(1,8) ,
40954	 => std_logic_vector(to_unsigned(1,8) ,
40955	 => std_logic_vector(to_unsigned(1,8) ,
40956	 => std_logic_vector(to_unsigned(1,8) ,
40957	 => std_logic_vector(to_unsigned(1,8) ,
40958	 => std_logic_vector(to_unsigned(1,8) ,
40959	 => std_logic_vector(to_unsigned(1,8) ,
40960	 => std_logic_vector(to_unsigned(1,8) ,
40961	 => std_logic_vector(to_unsigned(124,8) ,
40962	 => std_logic_vector(to_unsigned(119,8) ,
40963	 => std_logic_vector(to_unsigned(122,8) ,
40964	 => std_logic_vector(to_unsigned(121,8) ,
40965	 => std_logic_vector(to_unsigned(111,8) ,
40966	 => std_logic_vector(to_unsigned(103,8) ,
40967	 => std_logic_vector(to_unsigned(101,8) ,
40968	 => std_logic_vector(to_unsigned(93,8) ,
40969	 => std_logic_vector(to_unsigned(92,8) ,
40970	 => std_logic_vector(to_unsigned(92,8) ,
40971	 => std_logic_vector(to_unsigned(95,8) ,
40972	 => std_logic_vector(to_unsigned(93,8) ,
40973	 => std_logic_vector(to_unsigned(99,8) ,
40974	 => std_logic_vector(to_unsigned(99,8) ,
40975	 => std_logic_vector(to_unsigned(103,8) ,
40976	 => std_logic_vector(to_unsigned(109,8) ,
40977	 => std_logic_vector(to_unsigned(114,8) ,
40978	 => std_logic_vector(to_unsigned(119,8) ,
40979	 => std_logic_vector(to_unsigned(138,8) ,
40980	 => std_logic_vector(to_unsigned(147,8) ,
40981	 => std_logic_vector(to_unsigned(146,8) ,
40982	 => std_logic_vector(to_unsigned(136,8) ,
40983	 => std_logic_vector(to_unsigned(133,8) ,
40984	 => std_logic_vector(to_unsigned(146,8) ,
40985	 => std_logic_vector(to_unsigned(151,8) ,
40986	 => std_logic_vector(to_unsigned(151,8) ,
40987	 => std_logic_vector(to_unsigned(138,8) ,
40988	 => std_logic_vector(to_unsigned(139,8) ,
40989	 => std_logic_vector(to_unsigned(166,8) ,
40990	 => std_logic_vector(to_unsigned(72,8) ,
40991	 => std_logic_vector(to_unsigned(11,8) ,
40992	 => std_logic_vector(to_unsigned(16,8) ,
40993	 => std_logic_vector(to_unsigned(23,8) ,
40994	 => std_logic_vector(to_unsigned(11,8) ,
40995	 => std_logic_vector(to_unsigned(6,8) ,
40996	 => std_logic_vector(to_unsigned(3,8) ,
40997	 => std_logic_vector(to_unsigned(2,8) ,
40998	 => std_logic_vector(to_unsigned(1,8) ,
40999	 => std_logic_vector(to_unsigned(3,8) ,
41000	 => std_logic_vector(to_unsigned(13,8) ,
41001	 => std_logic_vector(to_unsigned(114,8) ,
41002	 => std_logic_vector(to_unsigned(170,8) ,
41003	 => std_logic_vector(to_unsigned(152,8) ,
41004	 => std_logic_vector(to_unsigned(159,8) ,
41005	 => std_logic_vector(to_unsigned(152,8) ,
41006	 => std_logic_vector(to_unsigned(156,8) ,
41007	 => std_logic_vector(to_unsigned(157,8) ,
41008	 => std_logic_vector(to_unsigned(163,8) ,
41009	 => std_logic_vector(to_unsigned(163,8) ,
41010	 => std_logic_vector(to_unsigned(157,8) ,
41011	 => std_logic_vector(to_unsigned(161,8) ,
41012	 => std_logic_vector(to_unsigned(161,8) ,
41013	 => std_logic_vector(to_unsigned(163,8) ,
41014	 => std_logic_vector(to_unsigned(161,8) ,
41015	 => std_logic_vector(to_unsigned(163,8) ,
41016	 => std_logic_vector(to_unsigned(163,8) ,
41017	 => std_logic_vector(to_unsigned(157,8) ,
41018	 => std_logic_vector(to_unsigned(163,8) ,
41019	 => std_logic_vector(to_unsigned(149,8) ,
41020	 => std_logic_vector(to_unsigned(142,8) ,
41021	 => std_logic_vector(to_unsigned(149,8) ,
41022	 => std_logic_vector(to_unsigned(61,8) ,
41023	 => std_logic_vector(to_unsigned(26,8) ,
41024	 => std_logic_vector(to_unsigned(48,8) ,
41025	 => std_logic_vector(to_unsigned(114,8) ,
41026	 => std_logic_vector(to_unsigned(156,8) ,
41027	 => std_logic_vector(to_unsigned(130,8) ,
41028	 => std_logic_vector(to_unsigned(130,8) ,
41029	 => std_logic_vector(to_unsigned(141,8) ,
41030	 => std_logic_vector(to_unsigned(141,8) ,
41031	 => std_logic_vector(to_unsigned(128,8) ,
41032	 => std_logic_vector(to_unsigned(121,8) ,
41033	 => std_logic_vector(to_unsigned(124,8) ,
41034	 => std_logic_vector(to_unsigned(122,8) ,
41035	 => std_logic_vector(to_unsigned(111,8) ,
41036	 => std_logic_vector(to_unsigned(125,8) ,
41037	 => std_logic_vector(to_unsigned(144,8) ,
41038	 => std_logic_vector(to_unsigned(23,8) ,
41039	 => std_logic_vector(to_unsigned(2,8) ,
41040	 => std_logic_vector(to_unsigned(11,8) ,
41041	 => std_logic_vector(to_unsigned(3,8) ,
41042	 => std_logic_vector(to_unsigned(0,8) ,
41043	 => std_logic_vector(to_unsigned(1,8) ,
41044	 => std_logic_vector(to_unsigned(0,8) ,
41045	 => std_logic_vector(to_unsigned(5,8) ,
41046	 => std_logic_vector(to_unsigned(99,8) ,
41047	 => std_logic_vector(to_unsigned(127,8) ,
41048	 => std_logic_vector(to_unsigned(101,8) ,
41049	 => std_logic_vector(to_unsigned(107,8) ,
41050	 => std_logic_vector(to_unsigned(109,8) ,
41051	 => std_logic_vector(to_unsigned(105,8) ,
41052	 => std_logic_vector(to_unsigned(111,8) ,
41053	 => std_logic_vector(to_unsigned(131,8) ,
41054	 => std_logic_vector(to_unsigned(116,8) ,
41055	 => std_logic_vector(to_unsigned(65,8) ,
41056	 => std_logic_vector(to_unsigned(99,8) ,
41057	 => std_logic_vector(to_unsigned(14,8) ,
41058	 => std_logic_vector(to_unsigned(2,8) ,
41059	 => std_logic_vector(to_unsigned(0,8) ,
41060	 => std_logic_vector(to_unsigned(3,8) ,
41061	 => std_logic_vector(to_unsigned(87,8) ,
41062	 => std_logic_vector(to_unsigned(138,8) ,
41063	 => std_logic_vector(to_unsigned(66,8) ,
41064	 => std_logic_vector(to_unsigned(3,8) ,
41065	 => std_logic_vector(to_unsigned(0,8) ,
41066	 => std_logic_vector(to_unsigned(0,8) ,
41067	 => std_logic_vector(to_unsigned(0,8) ,
41068	 => std_logic_vector(to_unsigned(0,8) ,
41069	 => std_logic_vector(to_unsigned(0,8) ,
41070	 => std_logic_vector(to_unsigned(27,8) ,
41071	 => std_logic_vector(to_unsigned(151,8) ,
41072	 => std_logic_vector(to_unsigned(133,8) ,
41073	 => std_logic_vector(to_unsigned(125,8) ,
41074	 => std_logic_vector(to_unsigned(136,8) ,
41075	 => std_logic_vector(to_unsigned(133,8) ,
41076	 => std_logic_vector(to_unsigned(134,8) ,
41077	 => std_logic_vector(to_unsigned(136,8) ,
41078	 => std_logic_vector(to_unsigned(125,8) ,
41079	 => std_logic_vector(to_unsigned(118,8) ,
41080	 => std_logic_vector(to_unsigned(109,8) ,
41081	 => std_logic_vector(to_unsigned(93,8) ,
41082	 => std_logic_vector(to_unsigned(70,8) ,
41083	 => std_logic_vector(to_unsigned(60,8) ,
41084	 => std_logic_vector(to_unsigned(39,8) ,
41085	 => std_logic_vector(to_unsigned(9,8) ,
41086	 => std_logic_vector(to_unsigned(13,8) ,
41087	 => std_logic_vector(to_unsigned(17,8) ,
41088	 => std_logic_vector(to_unsigned(6,8) ,
41089	 => std_logic_vector(to_unsigned(3,8) ,
41090	 => std_logic_vector(to_unsigned(3,8) ,
41091	 => std_logic_vector(to_unsigned(2,8) ,
41092	 => std_logic_vector(to_unsigned(2,8) ,
41093	 => std_logic_vector(to_unsigned(1,8) ,
41094	 => std_logic_vector(to_unsigned(1,8) ,
41095	 => std_logic_vector(to_unsigned(0,8) ,
41096	 => std_logic_vector(to_unsigned(0,8) ,
41097	 => std_logic_vector(to_unsigned(0,8) ,
41098	 => std_logic_vector(to_unsigned(2,8) ,
41099	 => std_logic_vector(to_unsigned(23,8) ,
41100	 => std_logic_vector(to_unsigned(17,8) ,
41101	 => std_logic_vector(to_unsigned(5,8) ,
41102	 => std_logic_vector(to_unsigned(1,8) ,
41103	 => std_logic_vector(to_unsigned(2,8) ,
41104	 => std_logic_vector(to_unsigned(1,8) ,
41105	 => std_logic_vector(to_unsigned(0,8) ,
41106	 => std_logic_vector(to_unsigned(1,8) ,
41107	 => std_logic_vector(to_unsigned(2,8) ,
41108	 => std_logic_vector(to_unsigned(2,8) ,
41109	 => std_logic_vector(to_unsigned(4,8) ,
41110	 => std_logic_vector(to_unsigned(6,8) ,
41111	 => std_logic_vector(to_unsigned(7,8) ,
41112	 => std_logic_vector(to_unsigned(5,8) ,
41113	 => std_logic_vector(to_unsigned(1,8) ,
41114	 => std_logic_vector(to_unsigned(1,8) ,
41115	 => std_logic_vector(to_unsigned(2,8) ,
41116	 => std_logic_vector(to_unsigned(0,8) ,
41117	 => std_logic_vector(to_unsigned(0,8) ,
41118	 => std_logic_vector(to_unsigned(0,8) ,
41119	 => std_logic_vector(to_unsigned(0,8) ,
41120	 => std_logic_vector(to_unsigned(0,8) ,
41121	 => std_logic_vector(to_unsigned(0,8) ,
41122	 => std_logic_vector(to_unsigned(0,8) ,
41123	 => std_logic_vector(to_unsigned(4,8) ,
41124	 => std_logic_vector(to_unsigned(10,8) ,
41125	 => std_logic_vector(to_unsigned(4,8) ,
41126	 => std_logic_vector(to_unsigned(2,8) ,
41127	 => std_logic_vector(to_unsigned(3,8) ,
41128	 => std_logic_vector(to_unsigned(4,8) ,
41129	 => std_logic_vector(to_unsigned(1,8) ,
41130	 => std_logic_vector(to_unsigned(1,8) ,
41131	 => std_logic_vector(to_unsigned(1,8) ,
41132	 => std_logic_vector(to_unsigned(1,8) ,
41133	 => std_logic_vector(to_unsigned(2,8) ,
41134	 => std_logic_vector(to_unsigned(2,8) ,
41135	 => std_logic_vector(to_unsigned(2,8) ,
41136	 => std_logic_vector(to_unsigned(1,8) ,
41137	 => std_logic_vector(to_unsigned(1,8) ,
41138	 => std_logic_vector(to_unsigned(0,8) ,
41139	 => std_logic_vector(to_unsigned(0,8) ,
41140	 => std_logic_vector(to_unsigned(0,8) ,
41141	 => std_logic_vector(to_unsigned(0,8) ,
41142	 => std_logic_vector(to_unsigned(3,8) ,
41143	 => std_logic_vector(to_unsigned(7,8) ,
41144	 => std_logic_vector(to_unsigned(5,8) ,
41145	 => std_logic_vector(to_unsigned(4,8) ,
41146	 => std_logic_vector(to_unsigned(2,8) ,
41147	 => std_logic_vector(to_unsigned(1,8) ,
41148	 => std_logic_vector(to_unsigned(1,8) ,
41149	 => std_logic_vector(to_unsigned(1,8) ,
41150	 => std_logic_vector(to_unsigned(1,8) ,
41151	 => std_logic_vector(to_unsigned(1,8) ,
41152	 => std_logic_vector(to_unsigned(7,8) ,
41153	 => std_logic_vector(to_unsigned(3,8) ,
41154	 => std_logic_vector(to_unsigned(0,8) ,
41155	 => std_logic_vector(to_unsigned(0,8) ,
41156	 => std_logic_vector(to_unsigned(0,8) ,
41157	 => std_logic_vector(to_unsigned(1,8) ,
41158	 => std_logic_vector(to_unsigned(1,8) ,
41159	 => std_logic_vector(to_unsigned(1,8) ,
41160	 => std_logic_vector(to_unsigned(1,8) ,
41161	 => std_logic_vector(to_unsigned(1,8) ,
41162	 => std_logic_vector(to_unsigned(1,8) ,
41163	 => std_logic_vector(to_unsigned(1,8) ,
41164	 => std_logic_vector(to_unsigned(1,8) ,
41165	 => std_logic_vector(to_unsigned(2,8) ,
41166	 => std_logic_vector(to_unsigned(3,8) ,
41167	 => std_logic_vector(to_unsigned(1,8) ,
41168	 => std_logic_vector(to_unsigned(4,8) ,
41169	 => std_logic_vector(to_unsigned(8,8) ,
41170	 => std_logic_vector(to_unsigned(10,8) ,
41171	 => std_logic_vector(to_unsigned(10,8) ,
41172	 => std_logic_vector(to_unsigned(3,8) ,
41173	 => std_logic_vector(to_unsigned(5,8) ,
41174	 => std_logic_vector(to_unsigned(81,8) ,
41175	 => std_logic_vector(to_unsigned(72,8) ,
41176	 => std_logic_vector(to_unsigned(79,8) ,
41177	 => std_logic_vector(to_unsigned(63,8) ,
41178	 => std_logic_vector(to_unsigned(58,8) ,
41179	 => std_logic_vector(to_unsigned(53,8) ,
41180	 => std_logic_vector(to_unsigned(20,8) ,
41181	 => std_logic_vector(to_unsigned(1,8) ,
41182	 => std_logic_vector(to_unsigned(0,8) ,
41183	 => std_logic_vector(to_unsigned(0,8) ,
41184	 => std_logic_vector(to_unsigned(1,8) ,
41185	 => std_logic_vector(to_unsigned(1,8) ,
41186	 => std_logic_vector(to_unsigned(2,8) ,
41187	 => std_logic_vector(to_unsigned(2,8) ,
41188	 => std_logic_vector(to_unsigned(1,8) ,
41189	 => std_logic_vector(to_unsigned(4,8) ,
41190	 => std_logic_vector(to_unsigned(76,8) ,
41191	 => std_logic_vector(to_unsigned(131,8) ,
41192	 => std_logic_vector(to_unsigned(138,8) ,
41193	 => std_logic_vector(to_unsigned(111,8) ,
41194	 => std_logic_vector(to_unsigned(99,8) ,
41195	 => std_logic_vector(to_unsigned(76,8) ,
41196	 => std_logic_vector(to_unsigned(15,8) ,
41197	 => std_logic_vector(to_unsigned(1,8) ,
41198	 => std_logic_vector(to_unsigned(1,8) ,
41199	 => std_logic_vector(to_unsigned(7,8) ,
41200	 => std_logic_vector(to_unsigned(7,8) ,
41201	 => std_logic_vector(to_unsigned(6,8) ,
41202	 => std_logic_vector(to_unsigned(6,8) ,
41203	 => std_logic_vector(to_unsigned(4,8) ,
41204	 => std_logic_vector(to_unsigned(2,8) ,
41205	 => std_logic_vector(to_unsigned(2,8) ,
41206	 => std_logic_vector(to_unsigned(1,8) ,
41207	 => std_logic_vector(to_unsigned(5,8) ,
41208	 => std_logic_vector(to_unsigned(18,8) ,
41209	 => std_logic_vector(to_unsigned(14,8) ,
41210	 => std_logic_vector(to_unsigned(3,8) ,
41211	 => std_logic_vector(to_unsigned(1,8) ,
41212	 => std_logic_vector(to_unsigned(2,8) ,
41213	 => std_logic_vector(to_unsigned(2,8) ,
41214	 => std_logic_vector(to_unsigned(2,8) ,
41215	 => std_logic_vector(to_unsigned(2,8) ,
41216	 => std_logic_vector(to_unsigned(3,8) ,
41217	 => std_logic_vector(to_unsigned(3,8) ,
41218	 => std_logic_vector(to_unsigned(3,8) ,
41219	 => std_logic_vector(to_unsigned(6,8) ,
41220	 => std_logic_vector(to_unsigned(5,8) ,
41221	 => std_logic_vector(to_unsigned(3,8) ,
41222	 => std_logic_vector(to_unsigned(2,8) ,
41223	 => std_logic_vector(to_unsigned(2,8) ,
41224	 => std_logic_vector(to_unsigned(3,8) ,
41225	 => std_logic_vector(to_unsigned(6,8) ,
41226	 => std_logic_vector(to_unsigned(30,8) ,
41227	 => std_logic_vector(to_unsigned(72,8) ,
41228	 => std_logic_vector(to_unsigned(36,8) ,
41229	 => std_logic_vector(to_unsigned(14,8) ,
41230	 => std_logic_vector(to_unsigned(5,8) ,
41231	 => std_logic_vector(to_unsigned(7,8) ,
41232	 => std_logic_vector(to_unsigned(13,8) ,
41233	 => std_logic_vector(to_unsigned(37,8) ,
41234	 => std_logic_vector(to_unsigned(30,8) ,
41235	 => std_logic_vector(to_unsigned(6,8) ,
41236	 => std_logic_vector(to_unsigned(1,8) ,
41237	 => std_logic_vector(to_unsigned(1,8) ,
41238	 => std_logic_vector(to_unsigned(2,8) ,
41239	 => std_logic_vector(to_unsigned(3,8) ,
41240	 => std_logic_vector(to_unsigned(3,8) ,
41241	 => std_logic_vector(to_unsigned(3,8) ,
41242	 => std_logic_vector(to_unsigned(2,8) ,
41243	 => std_logic_vector(to_unsigned(5,8) ,
41244	 => std_logic_vector(to_unsigned(6,8) ,
41245	 => std_logic_vector(to_unsigned(4,8) ,
41246	 => std_logic_vector(to_unsigned(8,8) ,
41247	 => std_logic_vector(to_unsigned(11,8) ,
41248	 => std_logic_vector(to_unsigned(7,8) ,
41249	 => std_logic_vector(to_unsigned(8,8) ,
41250	 => std_logic_vector(to_unsigned(5,8) ,
41251	 => std_logic_vector(to_unsigned(4,8) ,
41252	 => std_logic_vector(to_unsigned(3,8) ,
41253	 => std_logic_vector(to_unsigned(0,8) ,
41254	 => std_logic_vector(to_unsigned(1,8) ,
41255	 => std_logic_vector(to_unsigned(1,8) ,
41256	 => std_logic_vector(to_unsigned(0,8) ,
41257	 => std_logic_vector(to_unsigned(1,8) ,
41258	 => std_logic_vector(to_unsigned(1,8) ,
41259	 => std_logic_vector(to_unsigned(1,8) ,
41260	 => std_logic_vector(to_unsigned(1,8) ,
41261	 => std_logic_vector(to_unsigned(1,8) ,
41262	 => std_logic_vector(to_unsigned(2,8) ,
41263	 => std_logic_vector(to_unsigned(1,8) ,
41264	 => std_logic_vector(to_unsigned(1,8) ,
41265	 => std_logic_vector(to_unsigned(1,8) ,
41266	 => std_logic_vector(to_unsigned(1,8) ,
41267	 => std_logic_vector(to_unsigned(2,8) ,
41268	 => std_logic_vector(to_unsigned(1,8) ,
41269	 => std_logic_vector(to_unsigned(1,8) ,
41270	 => std_logic_vector(to_unsigned(1,8) ,
41271	 => std_logic_vector(to_unsigned(1,8) ,
41272	 => std_logic_vector(to_unsigned(1,8) ,
41273	 => std_logic_vector(to_unsigned(1,8) ,
41274	 => std_logic_vector(to_unsigned(2,8) ,
41275	 => std_logic_vector(to_unsigned(1,8) ,
41276	 => std_logic_vector(to_unsigned(1,8) ,
41277	 => std_logic_vector(to_unsigned(1,8) ,
41278	 => std_logic_vector(to_unsigned(1,8) ,
41279	 => std_logic_vector(to_unsigned(2,8) ,
41280	 => std_logic_vector(to_unsigned(1,8) ,
41281	 => std_logic_vector(to_unsigned(119,8) ,
41282	 => std_logic_vector(to_unsigned(121,8) ,
41283	 => std_logic_vector(to_unsigned(118,8) ,
41284	 => std_logic_vector(to_unsigned(122,8) ,
41285	 => std_logic_vector(to_unsigned(116,8) ,
41286	 => std_logic_vector(to_unsigned(99,8) ,
41287	 => std_logic_vector(to_unsigned(87,8) ,
41288	 => std_logic_vector(to_unsigned(84,8) ,
41289	 => std_logic_vector(to_unsigned(87,8) ,
41290	 => std_logic_vector(to_unsigned(88,8) ,
41291	 => std_logic_vector(to_unsigned(86,8) ,
41292	 => std_logic_vector(to_unsigned(88,8) ,
41293	 => std_logic_vector(to_unsigned(93,8) ,
41294	 => std_logic_vector(to_unsigned(93,8) ,
41295	 => std_logic_vector(to_unsigned(91,8) ,
41296	 => std_logic_vector(to_unsigned(103,8) ,
41297	 => std_logic_vector(to_unsigned(111,8) ,
41298	 => std_logic_vector(to_unsigned(116,8) ,
41299	 => std_logic_vector(to_unsigned(128,8) ,
41300	 => std_logic_vector(to_unsigned(149,8) ,
41301	 => std_logic_vector(to_unsigned(147,8) ,
41302	 => std_logic_vector(to_unsigned(121,8) ,
41303	 => std_logic_vector(to_unsigned(112,8) ,
41304	 => std_logic_vector(to_unsigned(136,8) ,
41305	 => std_logic_vector(to_unsigned(152,8) ,
41306	 => std_logic_vector(to_unsigned(149,8) ,
41307	 => std_logic_vector(to_unsigned(156,8) ,
41308	 => std_logic_vector(to_unsigned(163,8) ,
41309	 => std_logic_vector(to_unsigned(84,8) ,
41310	 => std_logic_vector(to_unsigned(14,8) ,
41311	 => std_logic_vector(to_unsigned(13,8) ,
41312	 => std_logic_vector(to_unsigned(22,8) ,
41313	 => std_logic_vector(to_unsigned(18,8) ,
41314	 => std_logic_vector(to_unsigned(12,8) ,
41315	 => std_logic_vector(to_unsigned(6,8) ,
41316	 => std_logic_vector(to_unsigned(3,8) ,
41317	 => std_logic_vector(to_unsigned(6,8) ,
41318	 => std_logic_vector(to_unsigned(46,8) ,
41319	 => std_logic_vector(to_unsigned(79,8) ,
41320	 => std_logic_vector(to_unsigned(124,8) ,
41321	 => std_logic_vector(to_unsigned(151,8) ,
41322	 => std_logic_vector(to_unsigned(146,8) ,
41323	 => std_logic_vector(to_unsigned(151,8) ,
41324	 => std_logic_vector(to_unsigned(156,8) ,
41325	 => std_logic_vector(to_unsigned(138,8) ,
41326	 => std_logic_vector(to_unsigned(138,8) ,
41327	 => std_logic_vector(to_unsigned(149,8) ,
41328	 => std_logic_vector(to_unsigned(163,8) ,
41329	 => std_logic_vector(to_unsigned(159,8) ,
41330	 => std_logic_vector(to_unsigned(154,8) ,
41331	 => std_logic_vector(to_unsigned(161,8) ,
41332	 => std_logic_vector(to_unsigned(164,8) ,
41333	 => std_logic_vector(to_unsigned(161,8) ,
41334	 => std_logic_vector(to_unsigned(164,8) ,
41335	 => std_logic_vector(to_unsigned(163,8) ,
41336	 => std_logic_vector(to_unsigned(161,8) ,
41337	 => std_logic_vector(to_unsigned(156,8) ,
41338	 => std_logic_vector(to_unsigned(156,8) ,
41339	 => std_logic_vector(to_unsigned(154,8) ,
41340	 => std_logic_vector(to_unsigned(142,8) ,
41341	 => std_logic_vector(to_unsigned(152,8) ,
41342	 => std_logic_vector(to_unsigned(152,8) ,
41343	 => std_logic_vector(to_unsigned(122,8) ,
41344	 => std_logic_vector(to_unsigned(125,8) ,
41345	 => std_logic_vector(to_unsigned(115,8) ,
41346	 => std_logic_vector(to_unsigned(104,8) ,
41347	 => std_logic_vector(to_unsigned(107,8) ,
41348	 => std_logic_vector(to_unsigned(134,8) ,
41349	 => std_logic_vector(to_unsigned(157,8) ,
41350	 => std_logic_vector(to_unsigned(154,8) ,
41351	 => std_logic_vector(to_unsigned(149,8) ,
41352	 => std_logic_vector(to_unsigned(144,8) ,
41353	 => std_logic_vector(to_unsigned(142,8) ,
41354	 => std_logic_vector(to_unsigned(141,8) ,
41355	 => std_logic_vector(to_unsigned(111,8) ,
41356	 => std_logic_vector(to_unsigned(114,8) ,
41357	 => std_logic_vector(to_unsigned(151,8) ,
41358	 => std_logic_vector(to_unsigned(30,8) ,
41359	 => std_logic_vector(to_unsigned(8,8) ,
41360	 => std_logic_vector(to_unsigned(12,8) ,
41361	 => std_logic_vector(to_unsigned(2,8) ,
41362	 => std_logic_vector(to_unsigned(1,8) ,
41363	 => std_logic_vector(to_unsigned(2,8) ,
41364	 => std_logic_vector(to_unsigned(2,8) ,
41365	 => std_logic_vector(to_unsigned(1,8) ,
41366	 => std_logic_vector(to_unsigned(51,8) ,
41367	 => std_logic_vector(to_unsigned(138,8) ,
41368	 => std_logic_vector(to_unsigned(103,8) ,
41369	 => std_logic_vector(to_unsigned(105,8) ,
41370	 => std_logic_vector(to_unsigned(101,8) ,
41371	 => std_logic_vector(to_unsigned(105,8) ,
41372	 => std_logic_vector(to_unsigned(111,8) ,
41373	 => std_logic_vector(to_unsigned(116,8) ,
41374	 => std_logic_vector(to_unsigned(105,8) ,
41375	 => std_logic_vector(to_unsigned(24,8) ,
41376	 => std_logic_vector(to_unsigned(8,8) ,
41377	 => std_logic_vector(to_unsigned(2,8) ,
41378	 => std_logic_vector(to_unsigned(2,8) ,
41379	 => std_logic_vector(to_unsigned(2,8) ,
41380	 => std_logic_vector(to_unsigned(3,8) ,
41381	 => std_logic_vector(to_unsigned(18,8) ,
41382	 => std_logic_vector(to_unsigned(130,8) ,
41383	 => std_logic_vector(to_unsigned(86,8) ,
41384	 => std_logic_vector(to_unsigned(3,8) ,
41385	 => std_logic_vector(to_unsigned(1,8) ,
41386	 => std_logic_vector(to_unsigned(1,8) ,
41387	 => std_logic_vector(to_unsigned(0,8) ,
41388	 => std_logic_vector(to_unsigned(1,8) ,
41389	 => std_logic_vector(to_unsigned(2,8) ,
41390	 => std_logic_vector(to_unsigned(1,8) ,
41391	 => std_logic_vector(to_unsigned(50,8) ,
41392	 => std_logic_vector(to_unsigned(142,8) ,
41393	 => std_logic_vector(to_unsigned(104,8) ,
41394	 => std_logic_vector(to_unsigned(109,8) ,
41395	 => std_logic_vector(to_unsigned(119,8) ,
41396	 => std_logic_vector(to_unsigned(128,8) ,
41397	 => std_logic_vector(to_unsigned(128,8) ,
41398	 => std_logic_vector(to_unsigned(130,8) ,
41399	 => std_logic_vector(to_unsigned(128,8) ,
41400	 => std_logic_vector(to_unsigned(128,8) ,
41401	 => std_logic_vector(to_unsigned(125,8) ,
41402	 => std_logic_vector(to_unsigned(128,8) ,
41403	 => std_logic_vector(to_unsigned(146,8) ,
41404	 => std_logic_vector(to_unsigned(45,8) ,
41405	 => std_logic_vector(to_unsigned(6,8) ,
41406	 => std_logic_vector(to_unsigned(34,8) ,
41407	 => std_logic_vector(to_unsigned(27,8) ,
41408	 => std_logic_vector(to_unsigned(3,8) ,
41409	 => std_logic_vector(to_unsigned(12,8) ,
41410	 => std_logic_vector(to_unsigned(80,8) ,
41411	 => std_logic_vector(to_unsigned(81,8) ,
41412	 => std_logic_vector(to_unsigned(76,8) ,
41413	 => std_logic_vector(to_unsigned(70,8) ,
41414	 => std_logic_vector(to_unsigned(51,8) ,
41415	 => std_logic_vector(to_unsigned(37,8) ,
41416	 => std_logic_vector(to_unsigned(22,8) ,
41417	 => std_logic_vector(to_unsigned(4,8) ,
41418	 => std_logic_vector(to_unsigned(4,8) ,
41419	 => std_logic_vector(to_unsigned(16,8) ,
41420	 => std_logic_vector(to_unsigned(10,8) ,
41421	 => std_logic_vector(to_unsigned(4,8) ,
41422	 => std_logic_vector(to_unsigned(1,8) ,
41423	 => std_logic_vector(to_unsigned(0,8) ,
41424	 => std_logic_vector(to_unsigned(1,8) ,
41425	 => std_logic_vector(to_unsigned(0,8) ,
41426	 => std_logic_vector(to_unsigned(1,8) ,
41427	 => std_logic_vector(to_unsigned(2,8) ,
41428	 => std_logic_vector(to_unsigned(1,8) ,
41429	 => std_logic_vector(to_unsigned(1,8) ,
41430	 => std_logic_vector(to_unsigned(2,8) ,
41431	 => std_logic_vector(to_unsigned(2,8) ,
41432	 => std_logic_vector(to_unsigned(4,8) ,
41433	 => std_logic_vector(to_unsigned(1,8) ,
41434	 => std_logic_vector(to_unsigned(3,8) ,
41435	 => std_logic_vector(to_unsigned(2,8) ,
41436	 => std_logic_vector(to_unsigned(0,8) ,
41437	 => std_logic_vector(to_unsigned(0,8) ,
41438	 => std_logic_vector(to_unsigned(0,8) ,
41439	 => std_logic_vector(to_unsigned(1,8) ,
41440	 => std_logic_vector(to_unsigned(1,8) ,
41441	 => std_logic_vector(to_unsigned(0,8) ,
41442	 => std_logic_vector(to_unsigned(1,8) ,
41443	 => std_logic_vector(to_unsigned(4,8) ,
41444	 => std_logic_vector(to_unsigned(8,8) ,
41445	 => std_logic_vector(to_unsigned(4,8) ,
41446	 => std_logic_vector(to_unsigned(2,8) ,
41447	 => std_logic_vector(to_unsigned(3,8) ,
41448	 => std_logic_vector(to_unsigned(1,8) ,
41449	 => std_logic_vector(to_unsigned(0,8) ,
41450	 => std_logic_vector(to_unsigned(1,8) ,
41451	 => std_logic_vector(to_unsigned(1,8) ,
41452	 => std_logic_vector(to_unsigned(1,8) ,
41453	 => std_logic_vector(to_unsigned(2,8) ,
41454	 => std_logic_vector(to_unsigned(1,8) ,
41455	 => std_logic_vector(to_unsigned(2,8) ,
41456	 => std_logic_vector(to_unsigned(1,8) ,
41457	 => std_logic_vector(to_unsigned(0,8) ,
41458	 => std_logic_vector(to_unsigned(0,8) ,
41459	 => std_logic_vector(to_unsigned(1,8) ,
41460	 => std_logic_vector(to_unsigned(1,8) ,
41461	 => std_logic_vector(to_unsigned(0,8) ,
41462	 => std_logic_vector(to_unsigned(0,8) ,
41463	 => std_logic_vector(to_unsigned(1,8) ,
41464	 => std_logic_vector(to_unsigned(1,8) ,
41465	 => std_logic_vector(to_unsigned(0,8) ,
41466	 => std_logic_vector(to_unsigned(0,8) ,
41467	 => std_logic_vector(to_unsigned(0,8) ,
41468	 => std_logic_vector(to_unsigned(11,8) ,
41469	 => std_logic_vector(to_unsigned(27,8) ,
41470	 => std_logic_vector(to_unsigned(12,8) ,
41471	 => std_logic_vector(to_unsigned(3,8) ,
41472	 => std_logic_vector(to_unsigned(10,8) ,
41473	 => std_logic_vector(to_unsigned(8,8) ,
41474	 => std_logic_vector(to_unsigned(0,8) ,
41475	 => std_logic_vector(to_unsigned(0,8) ,
41476	 => std_logic_vector(to_unsigned(0,8) ,
41477	 => std_logic_vector(to_unsigned(1,8) ,
41478	 => std_logic_vector(to_unsigned(1,8) ,
41479	 => std_logic_vector(to_unsigned(1,8) ,
41480	 => std_logic_vector(to_unsigned(1,8) ,
41481	 => std_logic_vector(to_unsigned(1,8) ,
41482	 => std_logic_vector(to_unsigned(1,8) ,
41483	 => std_logic_vector(to_unsigned(1,8) ,
41484	 => std_logic_vector(to_unsigned(1,8) ,
41485	 => std_logic_vector(to_unsigned(1,8) ,
41486	 => std_logic_vector(to_unsigned(3,8) ,
41487	 => std_logic_vector(to_unsigned(2,8) ,
41488	 => std_logic_vector(to_unsigned(4,8) ,
41489	 => std_logic_vector(to_unsigned(9,8) ,
41490	 => std_logic_vector(to_unsigned(9,8) ,
41491	 => std_logic_vector(to_unsigned(6,8) ,
41492	 => std_logic_vector(to_unsigned(3,8) ,
41493	 => std_logic_vector(to_unsigned(13,8) ,
41494	 => std_logic_vector(to_unsigned(112,8) ,
41495	 => std_logic_vector(to_unsigned(82,8) ,
41496	 => std_logic_vector(to_unsigned(61,8) ,
41497	 => std_logic_vector(to_unsigned(65,8) ,
41498	 => std_logic_vector(to_unsigned(67,8) ,
41499	 => std_logic_vector(to_unsigned(48,8) ,
41500	 => std_logic_vector(to_unsigned(23,8) ,
41501	 => std_logic_vector(to_unsigned(1,8) ,
41502	 => std_logic_vector(to_unsigned(0,8) ,
41503	 => std_logic_vector(to_unsigned(1,8) ,
41504	 => std_logic_vector(to_unsigned(1,8) ,
41505	 => std_logic_vector(to_unsigned(1,8) ,
41506	 => std_logic_vector(to_unsigned(2,8) ,
41507	 => std_logic_vector(to_unsigned(1,8) ,
41508	 => std_logic_vector(to_unsigned(1,8) ,
41509	 => std_logic_vector(to_unsigned(7,8) ,
41510	 => std_logic_vector(to_unsigned(104,8) ,
41511	 => std_logic_vector(to_unsigned(128,8) ,
41512	 => std_logic_vector(to_unsigned(128,8) ,
41513	 => std_logic_vector(to_unsigned(114,8) ,
41514	 => std_logic_vector(to_unsigned(80,8) ,
41515	 => std_logic_vector(to_unsigned(88,8) ,
41516	 => std_logic_vector(to_unsigned(26,8) ,
41517	 => std_logic_vector(to_unsigned(1,8) ,
41518	 => std_logic_vector(to_unsigned(2,8) ,
41519	 => std_logic_vector(to_unsigned(8,8) ,
41520	 => std_logic_vector(to_unsigned(9,8) ,
41521	 => std_logic_vector(to_unsigned(8,8) ,
41522	 => std_logic_vector(to_unsigned(8,8) ,
41523	 => std_logic_vector(to_unsigned(4,8) ,
41524	 => std_logic_vector(to_unsigned(2,8) ,
41525	 => std_logic_vector(to_unsigned(2,8) ,
41526	 => std_logic_vector(to_unsigned(1,8) ,
41527	 => std_logic_vector(to_unsigned(2,8) ,
41528	 => std_logic_vector(to_unsigned(13,8) ,
41529	 => std_logic_vector(to_unsigned(11,8) ,
41530	 => std_logic_vector(to_unsigned(3,8) ,
41531	 => std_logic_vector(to_unsigned(1,8) ,
41532	 => std_logic_vector(to_unsigned(2,8) ,
41533	 => std_logic_vector(to_unsigned(2,8) ,
41534	 => std_logic_vector(to_unsigned(2,8) ,
41535	 => std_logic_vector(to_unsigned(3,8) ,
41536	 => std_logic_vector(to_unsigned(2,8) ,
41537	 => std_logic_vector(to_unsigned(2,8) ,
41538	 => std_logic_vector(to_unsigned(4,8) ,
41539	 => std_logic_vector(to_unsigned(5,8) ,
41540	 => std_logic_vector(to_unsigned(4,8) ,
41541	 => std_logic_vector(to_unsigned(3,8) ,
41542	 => std_logic_vector(to_unsigned(1,8) ,
41543	 => std_logic_vector(to_unsigned(1,8) ,
41544	 => std_logic_vector(to_unsigned(0,8) ,
41545	 => std_logic_vector(to_unsigned(3,8) ,
41546	 => std_logic_vector(to_unsigned(46,8) ,
41547	 => std_logic_vector(to_unsigned(77,8) ,
41548	 => std_logic_vector(to_unsigned(49,8) ,
41549	 => std_logic_vector(to_unsigned(21,8) ,
41550	 => std_logic_vector(to_unsigned(8,8) ,
41551	 => std_logic_vector(to_unsigned(4,8) ,
41552	 => std_logic_vector(to_unsigned(13,8) ,
41553	 => std_logic_vector(to_unsigned(49,8) ,
41554	 => std_logic_vector(to_unsigned(33,8) ,
41555	 => std_logic_vector(to_unsigned(3,8) ,
41556	 => std_logic_vector(to_unsigned(1,8) ,
41557	 => std_logic_vector(to_unsigned(2,8) ,
41558	 => std_logic_vector(to_unsigned(2,8) ,
41559	 => std_logic_vector(to_unsigned(2,8) ,
41560	 => std_logic_vector(to_unsigned(3,8) ,
41561	 => std_logic_vector(to_unsigned(3,8) ,
41562	 => std_logic_vector(to_unsigned(2,8) ,
41563	 => std_logic_vector(to_unsigned(7,8) ,
41564	 => std_logic_vector(to_unsigned(6,8) ,
41565	 => std_logic_vector(to_unsigned(6,8) ,
41566	 => std_logic_vector(to_unsigned(10,8) ,
41567	 => std_logic_vector(to_unsigned(12,8) ,
41568	 => std_logic_vector(to_unsigned(8,8) ,
41569	 => std_logic_vector(to_unsigned(8,8) ,
41570	 => std_logic_vector(to_unsigned(7,8) ,
41571	 => std_logic_vector(to_unsigned(4,8) ,
41572	 => std_logic_vector(to_unsigned(5,8) ,
41573	 => std_logic_vector(to_unsigned(3,8) ,
41574	 => std_logic_vector(to_unsigned(1,8) ,
41575	 => std_logic_vector(to_unsigned(0,8) ,
41576	 => std_logic_vector(to_unsigned(1,8) ,
41577	 => std_logic_vector(to_unsigned(1,8) ,
41578	 => std_logic_vector(to_unsigned(1,8) ,
41579	 => std_logic_vector(to_unsigned(1,8) ,
41580	 => std_logic_vector(to_unsigned(1,8) ,
41581	 => std_logic_vector(to_unsigned(1,8) ,
41582	 => std_logic_vector(to_unsigned(1,8) ,
41583	 => std_logic_vector(to_unsigned(1,8) ,
41584	 => std_logic_vector(to_unsigned(1,8) ,
41585	 => std_logic_vector(to_unsigned(1,8) ,
41586	 => std_logic_vector(to_unsigned(1,8) ,
41587	 => std_logic_vector(to_unsigned(1,8) ,
41588	 => std_logic_vector(to_unsigned(1,8) ,
41589	 => std_logic_vector(to_unsigned(1,8) ,
41590	 => std_logic_vector(to_unsigned(1,8) ,
41591	 => std_logic_vector(to_unsigned(1,8) ,
41592	 => std_logic_vector(to_unsigned(1,8) ,
41593	 => std_logic_vector(to_unsigned(2,8) ,
41594	 => std_logic_vector(to_unsigned(2,8) ,
41595	 => std_logic_vector(to_unsigned(2,8) ,
41596	 => std_logic_vector(to_unsigned(2,8) ,
41597	 => std_logic_vector(to_unsigned(1,8) ,
41598	 => std_logic_vector(to_unsigned(2,8) ,
41599	 => std_logic_vector(to_unsigned(2,8) ,
41600	 => std_logic_vector(to_unsigned(2,8) ,
41601	 => std_logic_vector(to_unsigned(119,8) ,
41602	 => std_logic_vector(to_unsigned(122,8) ,
41603	 => std_logic_vector(to_unsigned(114,8) ,
41604	 => std_logic_vector(to_unsigned(107,8) ,
41605	 => std_logic_vector(to_unsigned(96,8) ,
41606	 => std_logic_vector(to_unsigned(82,8) ,
41607	 => std_logic_vector(to_unsigned(84,8) ,
41608	 => std_logic_vector(to_unsigned(84,8) ,
41609	 => std_logic_vector(to_unsigned(85,8) ,
41610	 => std_logic_vector(to_unsigned(78,8) ,
41611	 => std_logic_vector(to_unsigned(78,8) ,
41612	 => std_logic_vector(to_unsigned(77,8) ,
41613	 => std_logic_vector(to_unsigned(79,8) ,
41614	 => std_logic_vector(to_unsigned(86,8) ,
41615	 => std_logic_vector(to_unsigned(81,8) ,
41616	 => std_logic_vector(to_unsigned(119,8) ,
41617	 => std_logic_vector(to_unsigned(144,8) ,
41618	 => std_logic_vector(to_unsigned(133,8) ,
41619	 => std_logic_vector(to_unsigned(138,8) ,
41620	 => std_logic_vector(to_unsigned(131,8) ,
41621	 => std_logic_vector(to_unsigned(127,8) ,
41622	 => std_logic_vector(to_unsigned(111,8) ,
41623	 => std_logic_vector(to_unsigned(95,8) ,
41624	 => std_logic_vector(to_unsigned(122,8) ,
41625	 => std_logic_vector(to_unsigned(146,8) ,
41626	 => std_logic_vector(to_unsigned(154,8) ,
41627	 => std_logic_vector(to_unsigned(139,8) ,
41628	 => std_logic_vector(to_unsigned(54,8) ,
41629	 => std_logic_vector(to_unsigned(17,8) ,
41630	 => std_logic_vector(to_unsigned(19,8) ,
41631	 => std_logic_vector(to_unsigned(15,8) ,
41632	 => std_logic_vector(to_unsigned(10,8) ,
41633	 => std_logic_vector(to_unsigned(14,8) ,
41634	 => std_logic_vector(to_unsigned(7,8) ,
41635	 => std_logic_vector(to_unsigned(2,8) ,
41636	 => std_logic_vector(to_unsigned(9,8) ,
41637	 => std_logic_vector(to_unsigned(73,8) ,
41638	 => std_logic_vector(to_unsigned(179,8) ,
41639	 => std_logic_vector(to_unsigned(186,8) ,
41640	 => std_logic_vector(to_unsigned(146,8) ,
41641	 => std_logic_vector(to_unsigned(131,8) ,
41642	 => std_logic_vector(to_unsigned(144,8) ,
41643	 => std_logic_vector(to_unsigned(136,8) ,
41644	 => std_logic_vector(to_unsigned(152,8) ,
41645	 => std_logic_vector(to_unsigned(130,8) ,
41646	 => std_logic_vector(to_unsigned(136,8) ,
41647	 => std_logic_vector(to_unsigned(147,8) ,
41648	 => std_logic_vector(to_unsigned(159,8) ,
41649	 => std_logic_vector(to_unsigned(159,8) ,
41650	 => std_logic_vector(to_unsigned(147,8) ,
41651	 => std_logic_vector(to_unsigned(161,8) ,
41652	 => std_logic_vector(to_unsigned(159,8) ,
41653	 => std_logic_vector(to_unsigned(152,8) ,
41654	 => std_logic_vector(to_unsigned(142,8) ,
41655	 => std_logic_vector(to_unsigned(142,8) ,
41656	 => std_logic_vector(to_unsigned(149,8) ,
41657	 => std_logic_vector(to_unsigned(156,8) ,
41658	 => std_logic_vector(to_unsigned(157,8) ,
41659	 => std_logic_vector(to_unsigned(161,8) ,
41660	 => std_logic_vector(to_unsigned(164,8) ,
41661	 => std_logic_vector(to_unsigned(152,8) ,
41662	 => std_logic_vector(to_unsigned(141,8) ,
41663	 => std_logic_vector(to_unsigned(131,8) ,
41664	 => std_logic_vector(to_unsigned(136,8) ,
41665	 => std_logic_vector(to_unsigned(119,8) ,
41666	 => std_logic_vector(to_unsigned(118,8) ,
41667	 => std_logic_vector(to_unsigned(131,8) ,
41668	 => std_logic_vector(to_unsigned(149,8) ,
41669	 => std_logic_vector(to_unsigned(142,8) ,
41670	 => std_logic_vector(to_unsigned(149,8) ,
41671	 => std_logic_vector(to_unsigned(144,8) ,
41672	 => std_logic_vector(to_unsigned(141,8) ,
41673	 => std_logic_vector(to_unsigned(149,8) ,
41674	 => std_logic_vector(to_unsigned(154,8) ,
41675	 => std_logic_vector(to_unsigned(112,8) ,
41676	 => std_logic_vector(to_unsigned(127,8) ,
41677	 => std_logic_vector(to_unsigned(67,8) ,
41678	 => std_logic_vector(to_unsigned(14,8) ,
41679	 => std_logic_vector(to_unsigned(23,8) ,
41680	 => std_logic_vector(to_unsigned(6,8) ,
41681	 => std_logic_vector(to_unsigned(2,8) ,
41682	 => std_logic_vector(to_unsigned(2,8) ,
41683	 => std_logic_vector(to_unsigned(1,8) ,
41684	 => std_logic_vector(to_unsigned(2,8) ,
41685	 => std_logic_vector(to_unsigned(1,8) ,
41686	 => std_logic_vector(to_unsigned(38,8) ,
41687	 => std_logic_vector(to_unsigned(144,8) ,
41688	 => std_logic_vector(to_unsigned(111,8) ,
41689	 => std_logic_vector(to_unsigned(112,8) ,
41690	 => std_logic_vector(to_unsigned(107,8) ,
41691	 => std_logic_vector(to_unsigned(109,8) ,
41692	 => std_logic_vector(to_unsigned(111,8) ,
41693	 => std_logic_vector(to_unsigned(119,8) ,
41694	 => std_logic_vector(to_unsigned(104,8) ,
41695	 => std_logic_vector(to_unsigned(8,8) ,
41696	 => std_logic_vector(to_unsigned(0,8) ,
41697	 => std_logic_vector(to_unsigned(3,8) ,
41698	 => std_logic_vector(to_unsigned(4,8) ,
41699	 => std_logic_vector(to_unsigned(3,8) ,
41700	 => std_logic_vector(to_unsigned(5,8) ,
41701	 => std_logic_vector(to_unsigned(11,8) ,
41702	 => std_logic_vector(to_unsigned(46,8) ,
41703	 => std_logic_vector(to_unsigned(16,8) ,
41704	 => std_logic_vector(to_unsigned(0,8) ,
41705	 => std_logic_vector(to_unsigned(0,8) ,
41706	 => std_logic_vector(to_unsigned(0,8) ,
41707	 => std_logic_vector(to_unsigned(0,8) ,
41708	 => std_logic_vector(to_unsigned(4,8) ,
41709	 => std_logic_vector(to_unsigned(7,8) ,
41710	 => std_logic_vector(to_unsigned(0,8) ,
41711	 => std_logic_vector(to_unsigned(9,8) ,
41712	 => std_logic_vector(to_unsigned(124,8) ,
41713	 => std_logic_vector(to_unsigned(116,8) ,
41714	 => std_logic_vector(to_unsigned(111,8) ,
41715	 => std_logic_vector(to_unsigned(121,8) ,
41716	 => std_logic_vector(to_unsigned(127,8) ,
41717	 => std_logic_vector(to_unsigned(122,8) ,
41718	 => std_logic_vector(to_unsigned(131,8) ,
41719	 => std_logic_vector(to_unsigned(136,8) ,
41720	 => std_logic_vector(to_unsigned(128,8) ,
41721	 => std_logic_vector(to_unsigned(119,8) ,
41722	 => std_logic_vector(to_unsigned(119,8) ,
41723	 => std_logic_vector(to_unsigned(122,8) ,
41724	 => std_logic_vector(to_unsigned(13,8) ,
41725	 => std_logic_vector(to_unsigned(0,8) ,
41726	 => std_logic_vector(to_unsigned(10,8) ,
41727	 => std_logic_vector(to_unsigned(8,8) ,
41728	 => std_logic_vector(to_unsigned(0,8) ,
41729	 => std_logic_vector(to_unsigned(5,8) ,
41730	 => std_logic_vector(to_unsigned(107,8) ,
41731	 => std_logic_vector(to_unsigned(156,8) ,
41732	 => std_logic_vector(to_unsigned(157,8) ,
41733	 => std_logic_vector(to_unsigned(173,8) ,
41734	 => std_logic_vector(to_unsigned(163,8) ,
41735	 => std_logic_vector(to_unsigned(173,8) ,
41736	 => std_logic_vector(to_unsigned(101,8) ,
41737	 => std_logic_vector(to_unsigned(7,8) ,
41738	 => std_logic_vector(to_unsigned(4,8) ,
41739	 => std_logic_vector(to_unsigned(8,8) ,
41740	 => std_logic_vector(to_unsigned(4,8) ,
41741	 => std_logic_vector(to_unsigned(9,8) ,
41742	 => std_logic_vector(to_unsigned(54,8) ,
41743	 => std_logic_vector(to_unsigned(51,8) ,
41744	 => std_logic_vector(to_unsigned(43,8) ,
41745	 => std_logic_vector(to_unsigned(34,8) ,
41746	 => std_logic_vector(to_unsigned(25,8) ,
41747	 => std_logic_vector(to_unsigned(15,8) ,
41748	 => std_logic_vector(to_unsigned(9,8) ,
41749	 => std_logic_vector(to_unsigned(5,8) ,
41750	 => std_logic_vector(to_unsigned(2,8) ,
41751	 => std_logic_vector(to_unsigned(1,8) ,
41752	 => std_logic_vector(to_unsigned(4,8) ,
41753	 => std_logic_vector(to_unsigned(2,8) ,
41754	 => std_logic_vector(to_unsigned(4,8) ,
41755	 => std_logic_vector(to_unsigned(3,8) ,
41756	 => std_logic_vector(to_unsigned(1,8) ,
41757	 => std_logic_vector(to_unsigned(0,8) ,
41758	 => std_logic_vector(to_unsigned(0,8) ,
41759	 => std_logic_vector(to_unsigned(0,8) ,
41760	 => std_logic_vector(to_unsigned(0,8) ,
41761	 => std_logic_vector(to_unsigned(0,8) ,
41762	 => std_logic_vector(to_unsigned(4,8) ,
41763	 => std_logic_vector(to_unsigned(14,8) ,
41764	 => std_logic_vector(to_unsigned(6,8) ,
41765	 => std_logic_vector(to_unsigned(4,8) ,
41766	 => std_logic_vector(to_unsigned(3,8) ,
41767	 => std_logic_vector(to_unsigned(1,8) ,
41768	 => std_logic_vector(to_unsigned(1,8) ,
41769	 => std_logic_vector(to_unsigned(1,8) ,
41770	 => std_logic_vector(to_unsigned(1,8) ,
41771	 => std_logic_vector(to_unsigned(2,8) ,
41772	 => std_logic_vector(to_unsigned(2,8) ,
41773	 => std_logic_vector(to_unsigned(3,8) ,
41774	 => std_logic_vector(to_unsigned(3,8) ,
41775	 => std_logic_vector(to_unsigned(3,8) ,
41776	 => std_logic_vector(to_unsigned(3,8) ,
41777	 => std_logic_vector(to_unsigned(1,8) ,
41778	 => std_logic_vector(to_unsigned(0,8) ,
41779	 => std_logic_vector(to_unsigned(1,8) ,
41780	 => std_logic_vector(to_unsigned(1,8) ,
41781	 => std_logic_vector(to_unsigned(0,8) ,
41782	 => std_logic_vector(to_unsigned(0,8) ,
41783	 => std_logic_vector(to_unsigned(0,8) ,
41784	 => std_logic_vector(to_unsigned(0,8) ,
41785	 => std_logic_vector(to_unsigned(0,8) ,
41786	 => std_logic_vector(to_unsigned(0,8) ,
41787	 => std_logic_vector(to_unsigned(1,8) ,
41788	 => std_logic_vector(to_unsigned(13,8) ,
41789	 => std_logic_vector(to_unsigned(51,8) ,
41790	 => std_logic_vector(to_unsigned(42,8) ,
41791	 => std_logic_vector(to_unsigned(8,8) ,
41792	 => std_logic_vector(to_unsigned(17,8) ,
41793	 => std_logic_vector(to_unsigned(16,8) ,
41794	 => std_logic_vector(to_unsigned(1,8) ,
41795	 => std_logic_vector(to_unsigned(0,8) ,
41796	 => std_logic_vector(to_unsigned(1,8) ,
41797	 => std_logic_vector(to_unsigned(1,8) ,
41798	 => std_logic_vector(to_unsigned(1,8) ,
41799	 => std_logic_vector(to_unsigned(1,8) ,
41800	 => std_logic_vector(to_unsigned(1,8) ,
41801	 => std_logic_vector(to_unsigned(2,8) ,
41802	 => std_logic_vector(to_unsigned(1,8) ,
41803	 => std_logic_vector(to_unsigned(2,8) ,
41804	 => std_logic_vector(to_unsigned(2,8) ,
41805	 => std_logic_vector(to_unsigned(1,8) ,
41806	 => std_logic_vector(to_unsigned(2,8) ,
41807	 => std_logic_vector(to_unsigned(2,8) ,
41808	 => std_logic_vector(to_unsigned(2,8) ,
41809	 => std_logic_vector(to_unsigned(3,8) ,
41810	 => std_logic_vector(to_unsigned(4,8) ,
41811	 => std_logic_vector(to_unsigned(2,8) ,
41812	 => std_logic_vector(to_unsigned(2,8) ,
41813	 => std_logic_vector(to_unsigned(63,8) ,
41814	 => std_logic_vector(to_unsigned(119,8) ,
41815	 => std_logic_vector(to_unsigned(79,8) ,
41816	 => std_logic_vector(to_unsigned(65,8) ,
41817	 => std_logic_vector(to_unsigned(64,8) ,
41818	 => std_logic_vector(to_unsigned(51,8) ,
41819	 => std_logic_vector(to_unsigned(30,8) ,
41820	 => std_logic_vector(to_unsigned(8,8) ,
41821	 => std_logic_vector(to_unsigned(0,8) ,
41822	 => std_logic_vector(to_unsigned(0,8) ,
41823	 => std_logic_vector(to_unsigned(0,8) ,
41824	 => std_logic_vector(to_unsigned(1,8) ,
41825	 => std_logic_vector(to_unsigned(1,8) ,
41826	 => std_logic_vector(to_unsigned(1,8) ,
41827	 => std_logic_vector(to_unsigned(2,8) ,
41828	 => std_logic_vector(to_unsigned(0,8) ,
41829	 => std_logic_vector(to_unsigned(8,8) ,
41830	 => std_logic_vector(to_unsigned(111,8) ,
41831	 => std_logic_vector(to_unsigned(116,8) ,
41832	 => std_logic_vector(to_unsigned(61,8) ,
41833	 => std_logic_vector(to_unsigned(88,8) ,
41834	 => std_logic_vector(to_unsigned(107,8) ,
41835	 => std_logic_vector(to_unsigned(116,8) ,
41836	 => std_logic_vector(to_unsigned(37,8) ,
41837	 => std_logic_vector(to_unsigned(1,8) ,
41838	 => std_logic_vector(to_unsigned(2,8) ,
41839	 => std_logic_vector(to_unsigned(10,8) ,
41840	 => std_logic_vector(to_unsigned(8,8) ,
41841	 => std_logic_vector(to_unsigned(4,8) ,
41842	 => std_logic_vector(to_unsigned(6,8) ,
41843	 => std_logic_vector(to_unsigned(5,8) ,
41844	 => std_logic_vector(to_unsigned(3,8) ,
41845	 => std_logic_vector(to_unsigned(2,8) ,
41846	 => std_logic_vector(to_unsigned(0,8) ,
41847	 => std_logic_vector(to_unsigned(1,8) ,
41848	 => std_logic_vector(to_unsigned(11,8) ,
41849	 => std_logic_vector(to_unsigned(10,8) ,
41850	 => std_logic_vector(to_unsigned(2,8) ,
41851	 => std_logic_vector(to_unsigned(1,8) ,
41852	 => std_logic_vector(to_unsigned(2,8) ,
41853	 => std_logic_vector(to_unsigned(1,8) ,
41854	 => std_logic_vector(to_unsigned(1,8) ,
41855	 => std_logic_vector(to_unsigned(1,8) ,
41856	 => std_logic_vector(to_unsigned(1,8) ,
41857	 => std_logic_vector(to_unsigned(2,8) ,
41858	 => std_logic_vector(to_unsigned(5,8) ,
41859	 => std_logic_vector(to_unsigned(6,8) ,
41860	 => std_logic_vector(to_unsigned(5,8) ,
41861	 => std_logic_vector(to_unsigned(3,8) ,
41862	 => std_logic_vector(to_unsigned(1,8) ,
41863	 => std_logic_vector(to_unsigned(1,8) ,
41864	 => std_logic_vector(to_unsigned(0,8) ,
41865	 => std_logic_vector(to_unsigned(2,8) ,
41866	 => std_logic_vector(to_unsigned(50,8) ,
41867	 => std_logic_vector(to_unsigned(81,8) ,
41868	 => std_logic_vector(to_unsigned(64,8) ,
41869	 => std_logic_vector(to_unsigned(29,8) ,
41870	 => std_logic_vector(to_unsigned(13,8) ,
41871	 => std_logic_vector(to_unsigned(5,8) ,
41872	 => std_logic_vector(to_unsigned(13,8) ,
41873	 => std_logic_vector(to_unsigned(41,8) ,
41874	 => std_logic_vector(to_unsigned(41,8) ,
41875	 => std_logic_vector(to_unsigned(4,8) ,
41876	 => std_logic_vector(to_unsigned(1,8) ,
41877	 => std_logic_vector(to_unsigned(2,8) ,
41878	 => std_logic_vector(to_unsigned(1,8) ,
41879	 => std_logic_vector(to_unsigned(1,8) ,
41880	 => std_logic_vector(to_unsigned(2,8) ,
41881	 => std_logic_vector(to_unsigned(2,8) ,
41882	 => std_logic_vector(to_unsigned(2,8) ,
41883	 => std_logic_vector(to_unsigned(7,8) ,
41884	 => std_logic_vector(to_unsigned(7,8) ,
41885	 => std_logic_vector(to_unsigned(9,8) ,
41886	 => std_logic_vector(to_unsigned(18,8) ,
41887	 => std_logic_vector(to_unsigned(11,8) ,
41888	 => std_logic_vector(to_unsigned(8,8) ,
41889	 => std_logic_vector(to_unsigned(8,8) ,
41890	 => std_logic_vector(to_unsigned(7,8) ,
41891	 => std_logic_vector(to_unsigned(3,8) ,
41892	 => std_logic_vector(to_unsigned(6,8) ,
41893	 => std_logic_vector(to_unsigned(4,8) ,
41894	 => std_logic_vector(to_unsigned(1,8) ,
41895	 => std_logic_vector(to_unsigned(1,8) ,
41896	 => std_logic_vector(to_unsigned(1,8) ,
41897	 => std_logic_vector(to_unsigned(1,8) ,
41898	 => std_logic_vector(to_unsigned(1,8) ,
41899	 => std_logic_vector(to_unsigned(2,8) ,
41900	 => std_logic_vector(to_unsigned(1,8) ,
41901	 => std_logic_vector(to_unsigned(1,8) ,
41902	 => std_logic_vector(to_unsigned(1,8) ,
41903	 => std_logic_vector(to_unsigned(1,8) ,
41904	 => std_logic_vector(to_unsigned(1,8) ,
41905	 => std_logic_vector(to_unsigned(2,8) ,
41906	 => std_logic_vector(to_unsigned(2,8) ,
41907	 => std_logic_vector(to_unsigned(1,8) ,
41908	 => std_logic_vector(to_unsigned(2,8) ,
41909	 => std_logic_vector(to_unsigned(2,8) ,
41910	 => std_logic_vector(to_unsigned(1,8) ,
41911	 => std_logic_vector(to_unsigned(1,8) ,
41912	 => std_logic_vector(to_unsigned(1,8) ,
41913	 => std_logic_vector(to_unsigned(2,8) ,
41914	 => std_logic_vector(to_unsigned(1,8) ,
41915	 => std_logic_vector(to_unsigned(1,8) ,
41916	 => std_logic_vector(to_unsigned(3,8) ,
41917	 => std_logic_vector(to_unsigned(3,8) ,
41918	 => std_logic_vector(to_unsigned(3,8) ,
41919	 => std_logic_vector(to_unsigned(2,8) ,
41920	 => std_logic_vector(to_unsigned(3,8) ,
41921	 => std_logic_vector(to_unsigned(96,8) ,
41922	 => std_logic_vector(to_unsigned(91,8) ,
41923	 => std_logic_vector(to_unsigned(87,8) ,
41924	 => std_logic_vector(to_unsigned(86,8) ,
41925	 => std_logic_vector(to_unsigned(81,8) ,
41926	 => std_logic_vector(to_unsigned(71,8) ,
41927	 => std_logic_vector(to_unsigned(76,8) ,
41928	 => std_logic_vector(to_unsigned(78,8) ,
41929	 => std_logic_vector(to_unsigned(72,8) ,
41930	 => std_logic_vector(to_unsigned(77,8) ,
41931	 => std_logic_vector(to_unsigned(72,8) ,
41932	 => std_logic_vector(to_unsigned(38,8) ,
41933	 => std_logic_vector(to_unsigned(33,8) ,
41934	 => std_logic_vector(to_unsigned(69,8) ,
41935	 => std_logic_vector(to_unsigned(93,8) ,
41936	 => std_logic_vector(to_unsigned(112,8) ,
41937	 => std_logic_vector(to_unsigned(138,8) ,
41938	 => std_logic_vector(to_unsigned(131,8) ,
41939	 => std_logic_vector(to_unsigned(139,8) ,
41940	 => std_logic_vector(to_unsigned(138,8) ,
41941	 => std_logic_vector(to_unsigned(142,8) ,
41942	 => std_logic_vector(to_unsigned(138,8) ,
41943	 => std_logic_vector(to_unsigned(128,8) ,
41944	 => std_logic_vector(to_unsigned(134,8) ,
41945	 => std_logic_vector(to_unsigned(159,8) ,
41946	 => std_logic_vector(to_unsigned(152,8) ,
41947	 => std_logic_vector(to_unsigned(35,8) ,
41948	 => std_logic_vector(to_unsigned(8,8) ,
41949	 => std_logic_vector(to_unsigned(27,8) ,
41950	 => std_logic_vector(to_unsigned(19,8) ,
41951	 => std_logic_vector(to_unsigned(7,8) ,
41952	 => std_logic_vector(to_unsigned(6,8) ,
41953	 => std_logic_vector(to_unsigned(4,8) ,
41954	 => std_logic_vector(to_unsigned(2,8) ,
41955	 => std_logic_vector(to_unsigned(12,8) ,
41956	 => std_logic_vector(to_unsigned(80,8) ,
41957	 => std_logic_vector(to_unsigned(171,8) ,
41958	 => std_logic_vector(to_unsigned(151,8) ,
41959	 => std_logic_vector(to_unsigned(152,8) ,
41960	 => std_logic_vector(to_unsigned(136,8) ,
41961	 => std_logic_vector(to_unsigned(125,8) ,
41962	 => std_logic_vector(to_unsigned(144,8) ,
41963	 => std_logic_vector(to_unsigned(133,8) ,
41964	 => std_logic_vector(to_unsigned(141,8) ,
41965	 => std_logic_vector(to_unsigned(127,8) ,
41966	 => std_logic_vector(to_unsigned(131,8) ,
41967	 => std_logic_vector(to_unsigned(139,8) ,
41968	 => std_logic_vector(to_unsigned(152,8) ,
41969	 => std_logic_vector(to_unsigned(156,8) ,
41970	 => std_logic_vector(to_unsigned(146,8) ,
41971	 => std_logic_vector(to_unsigned(159,8) ,
41972	 => std_logic_vector(to_unsigned(161,8) ,
41973	 => std_logic_vector(to_unsigned(149,8) ,
41974	 => std_logic_vector(to_unsigned(125,8) ,
41975	 => std_logic_vector(to_unsigned(114,8) ,
41976	 => std_logic_vector(to_unsigned(121,8) ,
41977	 => std_logic_vector(to_unsigned(121,8) ,
41978	 => std_logic_vector(to_unsigned(133,8) ,
41979	 => std_logic_vector(to_unsigned(139,8) ,
41980	 => std_logic_vector(to_unsigned(136,8) ,
41981	 => std_logic_vector(to_unsigned(138,8) ,
41982	 => std_logic_vector(to_unsigned(141,8) ,
41983	 => std_logic_vector(to_unsigned(136,8) ,
41984	 => std_logic_vector(to_unsigned(138,8) ,
41985	 => std_logic_vector(to_unsigned(133,8) ,
41986	 => std_logic_vector(to_unsigned(136,8) ,
41987	 => std_logic_vector(to_unsigned(154,8) ,
41988	 => std_logic_vector(to_unsigned(157,8) ,
41989	 => std_logic_vector(to_unsigned(156,8) ,
41990	 => std_logic_vector(to_unsigned(154,8) ,
41991	 => std_logic_vector(to_unsigned(128,8) ,
41992	 => std_logic_vector(to_unsigned(124,8) ,
41993	 => std_logic_vector(to_unsigned(142,8) ,
41994	 => std_logic_vector(to_unsigned(144,8) ,
41995	 => std_logic_vector(to_unsigned(152,8) ,
41996	 => std_logic_vector(to_unsigned(130,8) ,
41997	 => std_logic_vector(to_unsigned(18,8) ,
41998	 => std_logic_vector(to_unsigned(19,8) ,
41999	 => std_logic_vector(to_unsigned(16,8) ,
42000	 => std_logic_vector(to_unsigned(3,8) ,
42001	 => std_logic_vector(to_unsigned(2,8) ,
42002	 => std_logic_vector(to_unsigned(1,8) ,
42003	 => std_logic_vector(to_unsigned(1,8) ,
42004	 => std_logic_vector(to_unsigned(2,8) ,
42005	 => std_logic_vector(to_unsigned(0,8) ,
42006	 => std_logic_vector(to_unsigned(25,8) ,
42007	 => std_logic_vector(to_unsigned(138,8) ,
42008	 => std_logic_vector(to_unsigned(108,8) ,
42009	 => std_logic_vector(to_unsigned(109,8) ,
42010	 => std_logic_vector(to_unsigned(109,8) ,
42011	 => std_logic_vector(to_unsigned(103,8) ,
42012	 => std_logic_vector(to_unsigned(112,8) ,
42013	 => std_logic_vector(to_unsigned(130,8) ,
42014	 => std_logic_vector(to_unsigned(69,8) ,
42015	 => std_logic_vector(to_unsigned(5,8) ,
42016	 => std_logic_vector(to_unsigned(10,8) ,
42017	 => std_logic_vector(to_unsigned(19,8) ,
42018	 => std_logic_vector(to_unsigned(24,8) ,
42019	 => std_logic_vector(to_unsigned(14,8) ,
42020	 => std_logic_vector(to_unsigned(18,8) ,
42021	 => std_logic_vector(to_unsigned(23,8) ,
42022	 => std_logic_vector(to_unsigned(6,8) ,
42023	 => std_logic_vector(to_unsigned(2,8) ,
42024	 => std_logic_vector(to_unsigned(5,8) ,
42025	 => std_logic_vector(to_unsigned(6,8) ,
42026	 => std_logic_vector(to_unsigned(3,8) ,
42027	 => std_logic_vector(to_unsigned(2,8) ,
42028	 => std_logic_vector(to_unsigned(7,8) ,
42029	 => std_logic_vector(to_unsigned(4,8) ,
42030	 => std_logic_vector(to_unsigned(2,8) ,
42031	 => std_logic_vector(to_unsigned(1,8) ,
42032	 => std_logic_vector(to_unsigned(31,8) ,
42033	 => std_logic_vector(to_unsigned(125,8) ,
42034	 => std_logic_vector(to_unsigned(115,8) ,
42035	 => std_logic_vector(to_unsigned(114,8) ,
42036	 => std_logic_vector(to_unsigned(114,8) ,
42037	 => std_logic_vector(to_unsigned(112,8) ,
42038	 => std_logic_vector(to_unsigned(109,8) ,
42039	 => std_logic_vector(to_unsigned(115,8) ,
42040	 => std_logic_vector(to_unsigned(115,8) ,
42041	 => std_logic_vector(to_unsigned(118,8) ,
42042	 => std_logic_vector(to_unsigned(115,8) ,
42043	 => std_logic_vector(to_unsigned(131,8) ,
42044	 => std_logic_vector(to_unsigned(37,8) ,
42045	 => std_logic_vector(to_unsigned(0,8) ,
42046	 => std_logic_vector(to_unsigned(1,8) ,
42047	 => std_logic_vector(to_unsigned(0,8) ,
42048	 => std_logic_vector(to_unsigned(0,8) ,
42049	 => std_logic_vector(to_unsigned(10,8) ,
42050	 => std_logic_vector(to_unsigned(104,8) ,
42051	 => std_logic_vector(to_unsigned(130,8) ,
42052	 => std_logic_vector(to_unsigned(134,8) ,
42053	 => std_logic_vector(to_unsigned(141,8) ,
42054	 => std_logic_vector(to_unsigned(131,8) ,
42055	 => std_logic_vector(to_unsigned(141,8) ,
42056	 => std_logic_vector(to_unsigned(28,8) ,
42057	 => std_logic_vector(to_unsigned(2,8) ,
42058	 => std_logic_vector(to_unsigned(7,8) ,
42059	 => std_logic_vector(to_unsigned(8,8) ,
42060	 => std_logic_vector(to_unsigned(2,8) ,
42061	 => std_logic_vector(to_unsigned(19,8) ,
42062	 => std_logic_vector(to_unsigned(166,8) ,
42063	 => std_logic_vector(to_unsigned(159,8) ,
42064	 => std_logic_vector(to_unsigned(146,8) ,
42065	 => std_logic_vector(to_unsigned(151,8) ,
42066	 => std_logic_vector(to_unsigned(141,8) ,
42067	 => std_logic_vector(to_unsigned(122,8) ,
42068	 => std_logic_vector(to_unsigned(114,8) ,
42069	 => std_logic_vector(to_unsigned(84,8) ,
42070	 => std_logic_vector(to_unsigned(78,8) ,
42071	 => std_logic_vector(to_unsigned(41,8) ,
42072	 => std_logic_vector(to_unsigned(7,8) ,
42073	 => std_logic_vector(to_unsigned(4,8) ,
42074	 => std_logic_vector(to_unsigned(6,8) ,
42075	 => std_logic_vector(to_unsigned(5,8) ,
42076	 => std_logic_vector(to_unsigned(2,8) ,
42077	 => std_logic_vector(to_unsigned(2,8) ,
42078	 => std_logic_vector(to_unsigned(2,8) ,
42079	 => std_logic_vector(to_unsigned(2,8) ,
42080	 => std_logic_vector(to_unsigned(2,8) ,
42081	 => std_logic_vector(to_unsigned(1,8) ,
42082	 => std_logic_vector(to_unsigned(9,8) ,
42083	 => std_logic_vector(to_unsigned(18,8) ,
42084	 => std_logic_vector(to_unsigned(5,8) ,
42085	 => std_logic_vector(to_unsigned(3,8) ,
42086	 => std_logic_vector(to_unsigned(1,8) ,
42087	 => std_logic_vector(to_unsigned(0,8) ,
42088	 => std_logic_vector(to_unsigned(0,8) ,
42089	 => std_logic_vector(to_unsigned(1,8) ,
42090	 => std_logic_vector(to_unsigned(1,8) ,
42091	 => std_logic_vector(to_unsigned(1,8) ,
42092	 => std_logic_vector(to_unsigned(2,8) ,
42093	 => std_logic_vector(to_unsigned(2,8) ,
42094	 => std_logic_vector(to_unsigned(2,8) ,
42095	 => std_logic_vector(to_unsigned(3,8) ,
42096	 => std_logic_vector(to_unsigned(2,8) ,
42097	 => std_logic_vector(to_unsigned(1,8) ,
42098	 => std_logic_vector(to_unsigned(1,8) ,
42099	 => std_logic_vector(to_unsigned(1,8) ,
42100	 => std_logic_vector(to_unsigned(2,8) ,
42101	 => std_logic_vector(to_unsigned(0,8) ,
42102	 => std_logic_vector(to_unsigned(0,8) ,
42103	 => std_logic_vector(to_unsigned(0,8) ,
42104	 => std_logic_vector(to_unsigned(0,8) ,
42105	 => std_logic_vector(to_unsigned(0,8) ,
42106	 => std_logic_vector(to_unsigned(1,8) ,
42107	 => std_logic_vector(to_unsigned(6,8) ,
42108	 => std_logic_vector(to_unsigned(14,8) ,
42109	 => std_logic_vector(to_unsigned(35,8) ,
42110	 => std_logic_vector(to_unsigned(39,8) ,
42111	 => std_logic_vector(to_unsigned(15,8) ,
42112	 => std_logic_vector(to_unsigned(33,8) ,
42113	 => std_logic_vector(to_unsigned(15,8) ,
42114	 => std_logic_vector(to_unsigned(1,8) ,
42115	 => std_logic_vector(to_unsigned(1,8) ,
42116	 => std_logic_vector(to_unsigned(1,8) ,
42117	 => std_logic_vector(to_unsigned(1,8) ,
42118	 => std_logic_vector(to_unsigned(1,8) ,
42119	 => std_logic_vector(to_unsigned(1,8) ,
42120	 => std_logic_vector(to_unsigned(1,8) ,
42121	 => std_logic_vector(to_unsigned(2,8) ,
42122	 => std_logic_vector(to_unsigned(1,8) ,
42123	 => std_logic_vector(to_unsigned(2,8) ,
42124	 => std_logic_vector(to_unsigned(3,8) ,
42125	 => std_logic_vector(to_unsigned(2,8) ,
42126	 => std_logic_vector(to_unsigned(0,8) ,
42127	 => std_logic_vector(to_unsigned(3,8) ,
42128	 => std_logic_vector(to_unsigned(44,8) ,
42129	 => std_logic_vector(to_unsigned(38,8) ,
42130	 => std_logic_vector(to_unsigned(23,8) ,
42131	 => std_logic_vector(to_unsigned(3,8) ,
42132	 => std_logic_vector(to_unsigned(5,8) ,
42133	 => std_logic_vector(to_unsigned(99,8) ,
42134	 => std_logic_vector(to_unsigned(99,8) ,
42135	 => std_logic_vector(to_unsigned(81,8) ,
42136	 => std_logic_vector(to_unsigned(73,8) ,
42137	 => std_logic_vector(to_unsigned(52,8) ,
42138	 => std_logic_vector(to_unsigned(35,8) ,
42139	 => std_logic_vector(to_unsigned(25,8) ,
42140	 => std_logic_vector(to_unsigned(4,8) ,
42141	 => std_logic_vector(to_unsigned(0,8) ,
42142	 => std_logic_vector(to_unsigned(0,8) ,
42143	 => std_logic_vector(to_unsigned(0,8) ,
42144	 => std_logic_vector(to_unsigned(1,8) ,
42145	 => std_logic_vector(to_unsigned(1,8) ,
42146	 => std_logic_vector(to_unsigned(1,8) ,
42147	 => std_logic_vector(to_unsigned(1,8) ,
42148	 => std_logic_vector(to_unsigned(1,8) ,
42149	 => std_logic_vector(to_unsigned(2,8) ,
42150	 => std_logic_vector(to_unsigned(10,8) ,
42151	 => std_logic_vector(to_unsigned(26,8) ,
42152	 => std_logic_vector(to_unsigned(35,8) ,
42153	 => std_logic_vector(to_unsigned(25,8) ,
42154	 => std_logic_vector(to_unsigned(33,8) ,
42155	 => std_logic_vector(to_unsigned(54,8) ,
42156	 => std_logic_vector(to_unsigned(10,8) ,
42157	 => std_logic_vector(to_unsigned(0,8) ,
42158	 => std_logic_vector(to_unsigned(1,8) ,
42159	 => std_logic_vector(to_unsigned(7,8) ,
42160	 => std_logic_vector(to_unsigned(6,8) ,
42161	 => std_logic_vector(to_unsigned(4,8) ,
42162	 => std_logic_vector(to_unsigned(3,8) ,
42163	 => std_logic_vector(to_unsigned(4,8) ,
42164	 => std_logic_vector(to_unsigned(4,8) ,
42165	 => std_logic_vector(to_unsigned(3,8) ,
42166	 => std_logic_vector(to_unsigned(1,8) ,
42167	 => std_logic_vector(to_unsigned(0,8) ,
42168	 => std_logic_vector(to_unsigned(8,8) ,
42169	 => std_logic_vector(to_unsigned(9,8) ,
42170	 => std_logic_vector(to_unsigned(3,8) ,
42171	 => std_logic_vector(to_unsigned(1,8) ,
42172	 => std_logic_vector(to_unsigned(1,8) ,
42173	 => std_logic_vector(to_unsigned(1,8) ,
42174	 => std_logic_vector(to_unsigned(2,8) ,
42175	 => std_logic_vector(to_unsigned(1,8) ,
42176	 => std_logic_vector(to_unsigned(1,8) ,
42177	 => std_logic_vector(to_unsigned(2,8) ,
42178	 => std_logic_vector(to_unsigned(4,8) ,
42179	 => std_logic_vector(to_unsigned(4,8) ,
42180	 => std_logic_vector(to_unsigned(4,8) ,
42181	 => std_logic_vector(to_unsigned(3,8) ,
42182	 => std_logic_vector(to_unsigned(1,8) ,
42183	 => std_logic_vector(to_unsigned(1,8) ,
42184	 => std_logic_vector(to_unsigned(0,8) ,
42185	 => std_logic_vector(to_unsigned(2,8) ,
42186	 => std_logic_vector(to_unsigned(50,8) ,
42187	 => std_logic_vector(to_unsigned(85,8) ,
42188	 => std_logic_vector(to_unsigned(64,8) ,
42189	 => std_logic_vector(to_unsigned(37,8) ,
42190	 => std_logic_vector(to_unsigned(20,8) ,
42191	 => std_logic_vector(to_unsigned(7,8) ,
42192	 => std_logic_vector(to_unsigned(8,8) ,
42193	 => std_logic_vector(to_unsigned(19,8) ,
42194	 => std_logic_vector(to_unsigned(40,8) ,
42195	 => std_logic_vector(to_unsigned(5,8) ,
42196	 => std_logic_vector(to_unsigned(0,8) ,
42197	 => std_logic_vector(to_unsigned(1,8) ,
42198	 => std_logic_vector(to_unsigned(1,8) ,
42199	 => std_logic_vector(to_unsigned(1,8) ,
42200	 => std_logic_vector(to_unsigned(2,8) ,
42201	 => std_logic_vector(to_unsigned(2,8) ,
42202	 => std_logic_vector(to_unsigned(2,8) ,
42203	 => std_logic_vector(to_unsigned(4,8) ,
42204	 => std_logic_vector(to_unsigned(3,8) ,
42205	 => std_logic_vector(to_unsigned(2,8) ,
42206	 => std_logic_vector(to_unsigned(11,8) ,
42207	 => std_logic_vector(to_unsigned(10,8) ,
42208	 => std_logic_vector(to_unsigned(7,8) ,
42209	 => std_logic_vector(to_unsigned(4,8) ,
42210	 => std_logic_vector(to_unsigned(4,8) ,
42211	 => std_logic_vector(to_unsigned(3,8) ,
42212	 => std_logic_vector(to_unsigned(8,8) ,
42213	 => std_logic_vector(to_unsigned(5,8) ,
42214	 => std_logic_vector(to_unsigned(1,8) ,
42215	 => std_logic_vector(to_unsigned(1,8) ,
42216	 => std_logic_vector(to_unsigned(1,8) ,
42217	 => std_logic_vector(to_unsigned(1,8) ,
42218	 => std_logic_vector(to_unsigned(1,8) ,
42219	 => std_logic_vector(to_unsigned(1,8) ,
42220	 => std_logic_vector(to_unsigned(1,8) ,
42221	 => std_logic_vector(to_unsigned(2,8) ,
42222	 => std_logic_vector(to_unsigned(1,8) ,
42223	 => std_logic_vector(to_unsigned(1,8) ,
42224	 => std_logic_vector(to_unsigned(1,8) ,
42225	 => std_logic_vector(to_unsigned(2,8) ,
42226	 => std_logic_vector(to_unsigned(2,8) ,
42227	 => std_logic_vector(to_unsigned(2,8) ,
42228	 => std_logic_vector(to_unsigned(2,8) ,
42229	 => std_logic_vector(to_unsigned(1,8) ,
42230	 => std_logic_vector(to_unsigned(2,8) ,
42231	 => std_logic_vector(to_unsigned(2,8) ,
42232	 => std_logic_vector(to_unsigned(2,8) ,
42233	 => std_logic_vector(to_unsigned(2,8) ,
42234	 => std_logic_vector(to_unsigned(2,8) ,
42235	 => std_logic_vector(to_unsigned(2,8) ,
42236	 => std_logic_vector(to_unsigned(2,8) ,
42237	 => std_logic_vector(to_unsigned(3,8) ,
42238	 => std_logic_vector(to_unsigned(2,8) ,
42239	 => std_logic_vector(to_unsigned(2,8) ,
42240	 => std_logic_vector(to_unsigned(3,8) ,
42241	 => std_logic_vector(to_unsigned(70,8) ,
42242	 => std_logic_vector(to_unsigned(71,8) ,
42243	 => std_logic_vector(to_unsigned(82,8) ,
42244	 => std_logic_vector(to_unsigned(95,8) ,
42245	 => std_logic_vector(to_unsigned(76,8) ,
42246	 => std_logic_vector(to_unsigned(55,8) ,
42247	 => std_logic_vector(to_unsigned(67,8) ,
42248	 => std_logic_vector(to_unsigned(71,8) ,
42249	 => std_logic_vector(to_unsigned(67,8) ,
42250	 => std_logic_vector(to_unsigned(68,8) ,
42251	 => std_logic_vector(to_unsigned(66,8) ,
42252	 => std_logic_vector(to_unsigned(44,8) ,
42253	 => std_logic_vector(to_unsigned(38,8) ,
42254	 => std_logic_vector(to_unsigned(68,8) ,
42255	 => std_logic_vector(to_unsigned(91,8) ,
42256	 => std_logic_vector(to_unsigned(109,8) ,
42257	 => std_logic_vector(to_unsigned(134,8) ,
42258	 => std_logic_vector(to_unsigned(130,8) ,
42259	 => std_logic_vector(to_unsigned(133,8) ,
42260	 => std_logic_vector(to_unsigned(133,8) ,
42261	 => std_logic_vector(to_unsigned(136,8) ,
42262	 => std_logic_vector(to_unsigned(141,8) ,
42263	 => std_logic_vector(to_unsigned(144,8) ,
42264	 => std_logic_vector(to_unsigned(131,8) ,
42265	 => std_logic_vector(to_unsigned(154,8) ,
42266	 => std_logic_vector(to_unsigned(134,8) ,
42267	 => std_logic_vector(to_unsigned(16,8) ,
42268	 => std_logic_vector(to_unsigned(2,8) ,
42269	 => std_logic_vector(to_unsigned(4,8) ,
42270	 => std_logic_vector(to_unsigned(3,8) ,
42271	 => std_logic_vector(to_unsigned(2,8) ,
42272	 => std_logic_vector(to_unsigned(3,8) ,
42273	 => std_logic_vector(to_unsigned(7,8) ,
42274	 => std_logic_vector(to_unsigned(28,8) ,
42275	 => std_logic_vector(to_unsigned(122,8) ,
42276	 => std_logic_vector(to_unsigned(173,8) ,
42277	 => std_logic_vector(to_unsigned(152,8) ,
42278	 => std_logic_vector(to_unsigned(149,8) ,
42279	 => std_logic_vector(to_unsigned(161,8) ,
42280	 => std_logic_vector(to_unsigned(134,8) ,
42281	 => std_logic_vector(to_unsigned(114,8) ,
42282	 => std_logic_vector(to_unsigned(134,8) ,
42283	 => std_logic_vector(to_unsigned(121,8) ,
42284	 => std_logic_vector(to_unsigned(138,8) ,
42285	 => std_logic_vector(to_unsigned(136,8) ,
42286	 => std_logic_vector(to_unsigned(128,8) ,
42287	 => std_logic_vector(to_unsigned(133,8) ,
42288	 => std_logic_vector(to_unsigned(152,8) ,
42289	 => std_logic_vector(to_unsigned(159,8) ,
42290	 => std_logic_vector(to_unsigned(156,8) ,
42291	 => std_logic_vector(to_unsigned(157,8) ,
42292	 => std_logic_vector(to_unsigned(157,8) ,
42293	 => std_logic_vector(to_unsigned(154,8) ,
42294	 => std_logic_vector(to_unsigned(128,8) ,
42295	 => std_logic_vector(to_unsigned(111,8) ,
42296	 => std_logic_vector(to_unsigned(111,8) ,
42297	 => std_logic_vector(to_unsigned(86,8) ,
42298	 => std_logic_vector(to_unsigned(105,8) ,
42299	 => std_logic_vector(to_unsigned(131,8) ,
42300	 => std_logic_vector(to_unsigned(119,8) ,
42301	 => std_logic_vector(to_unsigned(124,8) ,
42302	 => std_logic_vector(to_unsigned(118,8) ,
42303	 => std_logic_vector(to_unsigned(114,8) ,
42304	 => std_logic_vector(to_unsigned(112,8) ,
42305	 => std_logic_vector(to_unsigned(111,8) ,
42306	 => std_logic_vector(to_unsigned(114,8) ,
42307	 => std_logic_vector(to_unsigned(116,8) ,
42308	 => std_logic_vector(to_unsigned(116,8) ,
42309	 => std_logic_vector(to_unsigned(127,8) ,
42310	 => std_logic_vector(to_unsigned(127,8) ,
42311	 => std_logic_vector(to_unsigned(121,8) ,
42312	 => std_logic_vector(to_unsigned(116,8) ,
42313	 => std_logic_vector(to_unsigned(125,8) ,
42314	 => std_logic_vector(to_unsigned(146,8) ,
42315	 => std_logic_vector(to_unsigned(142,8) ,
42316	 => std_logic_vector(to_unsigned(45,8) ,
42317	 => std_logic_vector(to_unsigned(8,8) ,
42318	 => std_logic_vector(to_unsigned(16,8) ,
42319	 => std_logic_vector(to_unsigned(5,8) ,
42320	 => std_logic_vector(to_unsigned(4,8) ,
42321	 => std_logic_vector(to_unsigned(1,8) ,
42322	 => std_logic_vector(to_unsigned(3,8) ,
42323	 => std_logic_vector(to_unsigned(1,8) ,
42324	 => std_logic_vector(to_unsigned(1,8) ,
42325	 => std_logic_vector(to_unsigned(12,8) ,
42326	 => std_logic_vector(to_unsigned(80,8) ,
42327	 => std_logic_vector(to_unsigned(124,8) ,
42328	 => std_logic_vector(to_unsigned(105,8) ,
42329	 => std_logic_vector(to_unsigned(108,8) ,
42330	 => std_logic_vector(to_unsigned(100,8) ,
42331	 => std_logic_vector(to_unsigned(99,8) ,
42332	 => std_logic_vector(to_unsigned(114,8) ,
42333	 => std_logic_vector(to_unsigned(103,8) ,
42334	 => std_logic_vector(to_unsigned(12,8) ,
42335	 => std_logic_vector(to_unsigned(9,8) ,
42336	 => std_logic_vector(to_unsigned(63,8) ,
42337	 => std_logic_vector(to_unsigned(77,8) ,
42338	 => std_logic_vector(to_unsigned(62,8) ,
42339	 => std_logic_vector(to_unsigned(34,8) ,
42340	 => std_logic_vector(to_unsigned(35,8) ,
42341	 => std_logic_vector(to_unsigned(12,8) ,
42342	 => std_logic_vector(to_unsigned(4,8) ,
42343	 => std_logic_vector(to_unsigned(9,8) ,
42344	 => std_logic_vector(to_unsigned(15,8) ,
42345	 => std_logic_vector(to_unsigned(9,8) ,
42346	 => std_logic_vector(to_unsigned(3,8) ,
42347	 => std_logic_vector(to_unsigned(2,8) ,
42348	 => std_logic_vector(to_unsigned(1,8) ,
42349	 => std_logic_vector(to_unsigned(3,8) ,
42350	 => std_logic_vector(to_unsigned(4,8) ,
42351	 => std_logic_vector(to_unsigned(1,8) ,
42352	 => std_logic_vector(to_unsigned(34,8) ,
42353	 => std_logic_vector(to_unsigned(127,8) ,
42354	 => std_logic_vector(to_unsigned(116,8) ,
42355	 => std_logic_vector(to_unsigned(115,8) ,
42356	 => std_logic_vector(to_unsigned(112,8) ,
42357	 => std_logic_vector(to_unsigned(115,8) ,
42358	 => std_logic_vector(to_unsigned(114,8) ,
42359	 => std_logic_vector(to_unsigned(105,8) ,
42360	 => std_logic_vector(to_unsigned(111,8) ,
42361	 => std_logic_vector(to_unsigned(116,8) ,
42362	 => std_logic_vector(to_unsigned(105,8) ,
42363	 => std_logic_vector(to_unsigned(125,8) ,
42364	 => std_logic_vector(to_unsigned(52,8) ,
42365	 => std_logic_vector(to_unsigned(1,8) ,
42366	 => std_logic_vector(to_unsigned(1,8) ,
42367	 => std_logic_vector(to_unsigned(1,8) ,
42368	 => std_logic_vector(to_unsigned(0,8) ,
42369	 => std_logic_vector(to_unsigned(30,8) ,
42370	 => std_logic_vector(to_unsigned(136,8) ,
42371	 => std_logic_vector(to_unsigned(124,8) ,
42372	 => std_logic_vector(to_unsigned(127,8) ,
42373	 => std_logic_vector(to_unsigned(130,8) ,
42374	 => std_logic_vector(to_unsigned(136,8) ,
42375	 => std_logic_vector(to_unsigned(73,8) ,
42376	 => std_logic_vector(to_unsigned(4,8) ,
42377	 => std_logic_vector(to_unsigned(6,8) ,
42378	 => std_logic_vector(to_unsigned(8,8) ,
42379	 => std_logic_vector(to_unsigned(7,8) ,
42380	 => std_logic_vector(to_unsigned(2,8) ,
42381	 => std_logic_vector(to_unsigned(27,8) ,
42382	 => std_logic_vector(to_unsigned(156,8) ,
42383	 => std_logic_vector(to_unsigned(134,8) ,
42384	 => std_logic_vector(to_unsigned(127,8) ,
42385	 => std_logic_vector(to_unsigned(134,8) ,
42386	 => std_logic_vector(to_unsigned(139,8) ,
42387	 => std_logic_vector(to_unsigned(128,8) ,
42388	 => std_logic_vector(to_unsigned(142,8) ,
42389	 => std_logic_vector(to_unsigned(131,8) ,
42390	 => std_logic_vector(to_unsigned(154,8) ,
42391	 => std_logic_vector(to_unsigned(59,8) ,
42392	 => std_logic_vector(to_unsigned(2,8) ,
42393	 => std_logic_vector(to_unsigned(8,8) ,
42394	 => std_logic_vector(to_unsigned(7,8) ,
42395	 => std_logic_vector(to_unsigned(4,8) ,
42396	 => std_logic_vector(to_unsigned(1,8) ,
42397	 => std_logic_vector(to_unsigned(16,8) ,
42398	 => std_logic_vector(to_unsigned(93,8) ,
42399	 => std_logic_vector(to_unsigned(67,8) ,
42400	 => std_logic_vector(to_unsigned(8,8) ,
42401	 => std_logic_vector(to_unsigned(1,8) ,
42402	 => std_logic_vector(to_unsigned(17,8) ,
42403	 => std_logic_vector(to_unsigned(13,8) ,
42404	 => std_logic_vector(to_unsigned(2,8) ,
42405	 => std_logic_vector(to_unsigned(4,8) ,
42406	 => std_logic_vector(to_unsigned(5,8) ,
42407	 => std_logic_vector(to_unsigned(4,8) ,
42408	 => std_logic_vector(to_unsigned(2,8) ,
42409	 => std_logic_vector(to_unsigned(1,8) ,
42410	 => std_logic_vector(to_unsigned(2,8) ,
42411	 => std_logic_vector(to_unsigned(2,8) ,
42412	 => std_logic_vector(to_unsigned(1,8) ,
42413	 => std_logic_vector(to_unsigned(0,8) ,
42414	 => std_logic_vector(to_unsigned(0,8) ,
42415	 => std_logic_vector(to_unsigned(0,8) ,
42416	 => std_logic_vector(to_unsigned(0,8) ,
42417	 => std_logic_vector(to_unsigned(1,8) ,
42418	 => std_logic_vector(to_unsigned(1,8) ,
42419	 => std_logic_vector(to_unsigned(2,8) ,
42420	 => std_logic_vector(to_unsigned(3,8) ,
42421	 => std_logic_vector(to_unsigned(1,8) ,
42422	 => std_logic_vector(to_unsigned(0,8) ,
42423	 => std_logic_vector(to_unsigned(0,8) ,
42424	 => std_logic_vector(to_unsigned(0,8) ,
42425	 => std_logic_vector(to_unsigned(0,8) ,
42426	 => std_logic_vector(to_unsigned(0,8) ,
42427	 => std_logic_vector(to_unsigned(8,8) ,
42428	 => std_logic_vector(to_unsigned(42,8) ,
42429	 => std_logic_vector(to_unsigned(43,8) ,
42430	 => std_logic_vector(to_unsigned(22,8) ,
42431	 => std_logic_vector(to_unsigned(16,8) ,
42432	 => std_logic_vector(to_unsigned(15,8) ,
42433	 => std_logic_vector(to_unsigned(5,8) ,
42434	 => std_logic_vector(to_unsigned(1,8) ,
42435	 => std_logic_vector(to_unsigned(1,8) ,
42436	 => std_logic_vector(to_unsigned(1,8) ,
42437	 => std_logic_vector(to_unsigned(1,8) ,
42438	 => std_logic_vector(to_unsigned(2,8) ,
42439	 => std_logic_vector(to_unsigned(2,8) ,
42440	 => std_logic_vector(to_unsigned(2,8) ,
42441	 => std_logic_vector(to_unsigned(2,8) ,
42442	 => std_logic_vector(to_unsigned(1,8) ,
42443	 => std_logic_vector(to_unsigned(1,8) ,
42444	 => std_logic_vector(to_unsigned(2,8) ,
42445	 => std_logic_vector(to_unsigned(2,8) ,
42446	 => std_logic_vector(to_unsigned(0,8) ,
42447	 => std_logic_vector(to_unsigned(5,8) ,
42448	 => std_logic_vector(to_unsigned(79,8) ,
42449	 => std_logic_vector(to_unsigned(124,8) ,
42450	 => std_logic_vector(to_unsigned(21,8) ,
42451	 => std_logic_vector(to_unsigned(0,8) ,
42452	 => std_logic_vector(to_unsigned(15,8) ,
42453	 => std_logic_vector(to_unsigned(107,8) ,
42454	 => std_logic_vector(to_unsigned(72,8) ,
42455	 => std_logic_vector(to_unsigned(88,8) ,
42456	 => std_logic_vector(to_unsigned(68,8) ,
42457	 => std_logic_vector(to_unsigned(45,8) ,
42458	 => std_logic_vector(to_unsigned(37,8) ,
42459	 => std_logic_vector(to_unsigned(14,8) ,
42460	 => std_logic_vector(to_unsigned(1,8) ,
42461	 => std_logic_vector(to_unsigned(0,8) ,
42462	 => std_logic_vector(to_unsigned(0,8) ,
42463	 => std_logic_vector(to_unsigned(1,8) ,
42464	 => std_logic_vector(to_unsigned(1,8) ,
42465	 => std_logic_vector(to_unsigned(1,8) ,
42466	 => std_logic_vector(to_unsigned(1,8) ,
42467	 => std_logic_vector(to_unsigned(1,8) ,
42468	 => std_logic_vector(to_unsigned(1,8) ,
42469	 => std_logic_vector(to_unsigned(2,8) ,
42470	 => std_logic_vector(to_unsigned(0,8) ,
42471	 => std_logic_vector(to_unsigned(1,8) ,
42472	 => std_logic_vector(to_unsigned(63,8) ,
42473	 => std_logic_vector(to_unsigned(112,8) ,
42474	 => std_logic_vector(to_unsigned(51,8) ,
42475	 => std_logic_vector(to_unsigned(7,8) ,
42476	 => std_logic_vector(to_unsigned(0,8) ,
42477	 => std_logic_vector(to_unsigned(0,8) ,
42478	 => std_logic_vector(to_unsigned(1,8) ,
42479	 => std_logic_vector(to_unsigned(5,8) ,
42480	 => std_logic_vector(to_unsigned(8,8) ,
42481	 => std_logic_vector(to_unsigned(7,8) ,
42482	 => std_logic_vector(to_unsigned(3,8) ,
42483	 => std_logic_vector(to_unsigned(3,8) ,
42484	 => std_logic_vector(to_unsigned(3,8) ,
42485	 => std_logic_vector(to_unsigned(3,8) ,
42486	 => std_logic_vector(to_unsigned(1,8) ,
42487	 => std_logic_vector(to_unsigned(1,8) ,
42488	 => std_logic_vector(to_unsigned(6,8) ,
42489	 => std_logic_vector(to_unsigned(6,8) ,
42490	 => std_logic_vector(to_unsigned(3,8) ,
42491	 => std_logic_vector(to_unsigned(1,8) ,
42492	 => std_logic_vector(to_unsigned(1,8) ,
42493	 => std_logic_vector(to_unsigned(1,8) ,
42494	 => std_logic_vector(to_unsigned(1,8) ,
42495	 => std_logic_vector(to_unsigned(1,8) ,
42496	 => std_logic_vector(to_unsigned(1,8) ,
42497	 => std_logic_vector(to_unsigned(2,8) ,
42498	 => std_logic_vector(to_unsigned(3,8) ,
42499	 => std_logic_vector(to_unsigned(2,8) ,
42500	 => std_logic_vector(to_unsigned(3,8) ,
42501	 => std_logic_vector(to_unsigned(3,8) ,
42502	 => std_logic_vector(to_unsigned(0,8) ,
42503	 => std_logic_vector(to_unsigned(1,8) ,
42504	 => std_logic_vector(to_unsigned(0,8) ,
42505	 => std_logic_vector(to_unsigned(4,8) ,
42506	 => std_logic_vector(to_unsigned(52,8) ,
42507	 => std_logic_vector(to_unsigned(59,8) ,
42508	 => std_logic_vector(to_unsigned(49,8) ,
42509	 => std_logic_vector(to_unsigned(29,8) ,
42510	 => std_logic_vector(to_unsigned(15,8) ,
42511	 => std_logic_vector(to_unsigned(6,8) ,
42512	 => std_logic_vector(to_unsigned(5,8) ,
42513	 => std_logic_vector(to_unsigned(12,8) ,
42514	 => std_logic_vector(to_unsigned(35,8) ,
42515	 => std_logic_vector(to_unsigned(8,8) ,
42516	 => std_logic_vector(to_unsigned(0,8) ,
42517	 => std_logic_vector(to_unsigned(1,8) ,
42518	 => std_logic_vector(to_unsigned(1,8) ,
42519	 => std_logic_vector(to_unsigned(1,8) ,
42520	 => std_logic_vector(to_unsigned(1,8) ,
42521	 => std_logic_vector(to_unsigned(1,8) ,
42522	 => std_logic_vector(to_unsigned(2,8) ,
42523	 => std_logic_vector(to_unsigned(2,8) ,
42524	 => std_logic_vector(to_unsigned(1,8) ,
42525	 => std_logic_vector(to_unsigned(1,8) ,
42526	 => std_logic_vector(to_unsigned(3,8) ,
42527	 => std_logic_vector(to_unsigned(4,8) ,
42528	 => std_logic_vector(to_unsigned(5,8) ,
42529	 => std_logic_vector(to_unsigned(3,8) ,
42530	 => std_logic_vector(to_unsigned(2,8) ,
42531	 => std_logic_vector(to_unsigned(1,8) ,
42532	 => std_logic_vector(to_unsigned(2,8) ,
42533	 => std_logic_vector(to_unsigned(2,8) ,
42534	 => std_logic_vector(to_unsigned(1,8) ,
42535	 => std_logic_vector(to_unsigned(1,8) ,
42536	 => std_logic_vector(to_unsigned(1,8) ,
42537	 => std_logic_vector(to_unsigned(1,8) ,
42538	 => std_logic_vector(to_unsigned(1,8) ,
42539	 => std_logic_vector(to_unsigned(1,8) ,
42540	 => std_logic_vector(to_unsigned(1,8) ,
42541	 => std_logic_vector(to_unsigned(1,8) ,
42542	 => std_logic_vector(to_unsigned(2,8) ,
42543	 => std_logic_vector(to_unsigned(1,8) ,
42544	 => std_logic_vector(to_unsigned(1,8) ,
42545	 => std_logic_vector(to_unsigned(1,8) ,
42546	 => std_logic_vector(to_unsigned(2,8) ,
42547	 => std_logic_vector(to_unsigned(2,8) ,
42548	 => std_logic_vector(to_unsigned(1,8) ,
42549	 => std_logic_vector(to_unsigned(1,8) ,
42550	 => std_logic_vector(to_unsigned(2,8) ,
42551	 => std_logic_vector(to_unsigned(1,8) ,
42552	 => std_logic_vector(to_unsigned(2,8) ,
42553	 => std_logic_vector(to_unsigned(2,8) ,
42554	 => std_logic_vector(to_unsigned(2,8) ,
42555	 => std_logic_vector(to_unsigned(2,8) ,
42556	 => std_logic_vector(to_unsigned(1,8) ,
42557	 => std_logic_vector(to_unsigned(1,8) ,
42558	 => std_logic_vector(to_unsigned(2,8) ,
42559	 => std_logic_vector(to_unsigned(2,8) ,
42560	 => std_logic_vector(to_unsigned(2,8) ,
42561	 => std_logic_vector(to_unsigned(80,8) ,
42562	 => std_logic_vector(to_unsigned(82,8) ,
42563	 => std_logic_vector(to_unsigned(99,8) ,
42564	 => std_logic_vector(to_unsigned(93,8) ,
42565	 => std_logic_vector(to_unsigned(84,8) ,
42566	 => std_logic_vector(to_unsigned(80,8) ,
42567	 => std_logic_vector(to_unsigned(91,8) ,
42568	 => std_logic_vector(to_unsigned(69,8) ,
42569	 => std_logic_vector(to_unsigned(62,8) ,
42570	 => std_logic_vector(to_unsigned(65,8) ,
42571	 => std_logic_vector(to_unsigned(61,8) ,
42572	 => std_logic_vector(to_unsigned(68,8) ,
42573	 => std_logic_vector(to_unsigned(66,8) ,
42574	 => std_logic_vector(to_unsigned(62,8) ,
42575	 => std_logic_vector(to_unsigned(77,8) ,
42576	 => std_logic_vector(to_unsigned(109,8) ,
42577	 => std_logic_vector(to_unsigned(109,8) ,
42578	 => std_logic_vector(to_unsigned(108,8) ,
42579	 => std_logic_vector(to_unsigned(131,8) ,
42580	 => std_logic_vector(to_unsigned(128,8) ,
42581	 => std_logic_vector(to_unsigned(127,8) ,
42582	 => std_logic_vector(to_unsigned(139,8) ,
42583	 => std_logic_vector(to_unsigned(131,8) ,
42584	 => std_logic_vector(to_unsigned(130,8) ,
42585	 => std_logic_vector(to_unsigned(141,8) ,
42586	 => std_logic_vector(to_unsigned(138,8) ,
42587	 => std_logic_vector(to_unsigned(92,8) ,
42588	 => std_logic_vector(to_unsigned(30,8) ,
42589	 => std_logic_vector(to_unsigned(14,8) ,
42590	 => std_logic_vector(to_unsigned(22,8) ,
42591	 => std_logic_vector(to_unsigned(32,8) ,
42592	 => std_logic_vector(to_unsigned(63,8) ,
42593	 => std_logic_vector(to_unsigned(111,8) ,
42594	 => std_logic_vector(to_unsigned(151,8) ,
42595	 => std_logic_vector(to_unsigned(161,8) ,
42596	 => std_logic_vector(to_unsigned(152,8) ,
42597	 => std_logic_vector(to_unsigned(152,8) ,
42598	 => std_logic_vector(to_unsigned(156,8) ,
42599	 => std_logic_vector(to_unsigned(157,8) ,
42600	 => std_logic_vector(to_unsigned(136,8) ,
42601	 => std_logic_vector(to_unsigned(112,8) ,
42602	 => std_logic_vector(to_unsigned(122,8) ,
42603	 => std_logic_vector(to_unsigned(104,8) ,
42604	 => std_logic_vector(to_unsigned(128,8) ,
42605	 => std_logic_vector(to_unsigned(128,8) ,
42606	 => std_logic_vector(to_unsigned(114,8) ,
42607	 => std_logic_vector(to_unsigned(124,8) ,
42608	 => std_logic_vector(to_unsigned(141,8) ,
42609	 => std_logic_vector(to_unsigned(157,8) ,
42610	 => std_logic_vector(to_unsigned(147,8) ,
42611	 => std_logic_vector(to_unsigned(157,8) ,
42612	 => std_logic_vector(to_unsigned(157,8) ,
42613	 => std_logic_vector(to_unsigned(151,8) ,
42614	 => std_logic_vector(to_unsigned(131,8) ,
42615	 => std_logic_vector(to_unsigned(118,8) ,
42616	 => std_logic_vector(to_unsigned(115,8) ,
42617	 => std_logic_vector(to_unsigned(115,8) ,
42618	 => std_logic_vector(to_unsigned(116,8) ,
42619	 => std_logic_vector(to_unsigned(122,8) ,
42620	 => std_logic_vector(to_unsigned(118,8) ,
42621	 => std_logic_vector(to_unsigned(127,8) ,
42622	 => std_logic_vector(to_unsigned(114,8) ,
42623	 => std_logic_vector(to_unsigned(103,8) ,
42624	 => std_logic_vector(to_unsigned(112,8) ,
42625	 => std_logic_vector(to_unsigned(111,8) ,
42626	 => std_logic_vector(to_unsigned(103,8) ,
42627	 => std_logic_vector(to_unsigned(104,8) ,
42628	 => std_logic_vector(to_unsigned(95,8) ,
42629	 => std_logic_vector(to_unsigned(91,8) ,
42630	 => std_logic_vector(to_unsigned(93,8) ,
42631	 => std_logic_vector(to_unsigned(95,8) ,
42632	 => std_logic_vector(to_unsigned(88,8) ,
42633	 => std_logic_vector(to_unsigned(103,8) ,
42634	 => std_logic_vector(to_unsigned(101,8) ,
42635	 => std_logic_vector(to_unsigned(33,8) ,
42636	 => std_logic_vector(to_unsigned(6,8) ,
42637	 => std_logic_vector(to_unsigned(10,8) ,
42638	 => std_logic_vector(to_unsigned(6,8) ,
42639	 => std_logic_vector(to_unsigned(4,8) ,
42640	 => std_logic_vector(to_unsigned(2,8) ,
42641	 => std_logic_vector(to_unsigned(3,8) ,
42642	 => std_logic_vector(to_unsigned(29,8) ,
42643	 => std_logic_vector(to_unsigned(32,8) ,
42644	 => std_logic_vector(to_unsigned(45,8) ,
42645	 => std_logic_vector(to_unsigned(119,8) ,
42646	 => std_logic_vector(to_unsigned(118,8) ,
42647	 => std_logic_vector(to_unsigned(95,8) ,
42648	 => std_logic_vector(to_unsigned(97,8) ,
42649	 => std_logic_vector(to_unsigned(92,8) ,
42650	 => std_logic_vector(to_unsigned(93,8) ,
42651	 => std_logic_vector(to_unsigned(96,8) ,
42652	 => std_logic_vector(to_unsigned(107,8) ,
42653	 => std_logic_vector(to_unsigned(26,8) ,
42654	 => std_logic_vector(to_unsigned(2,8) ,
42655	 => std_logic_vector(to_unsigned(49,8) ,
42656	 => std_logic_vector(to_unsigned(79,8) ,
42657	 => std_logic_vector(to_unsigned(47,8) ,
42658	 => std_logic_vector(to_unsigned(51,8) ,
42659	 => std_logic_vector(to_unsigned(37,8) ,
42660	 => std_logic_vector(to_unsigned(10,8) ,
42661	 => std_logic_vector(to_unsigned(2,8) ,
42662	 => std_logic_vector(to_unsigned(5,8) ,
42663	 => std_logic_vector(to_unsigned(14,8) ,
42664	 => std_logic_vector(to_unsigned(8,8) ,
42665	 => std_logic_vector(to_unsigned(1,8) ,
42666	 => std_logic_vector(to_unsigned(1,8) ,
42667	 => std_logic_vector(to_unsigned(1,8) ,
42668	 => std_logic_vector(to_unsigned(2,8) ,
42669	 => std_logic_vector(to_unsigned(3,8) ,
42670	 => std_logic_vector(to_unsigned(2,8) ,
42671	 => std_logic_vector(to_unsigned(35,8) ,
42672	 => std_logic_vector(to_unsigned(130,8) ,
42673	 => std_logic_vector(to_unsigned(111,8) ,
42674	 => std_logic_vector(to_unsigned(112,8) ,
42675	 => std_logic_vector(to_unsigned(119,8) ,
42676	 => std_logic_vector(to_unsigned(121,8) ,
42677	 => std_logic_vector(to_unsigned(115,8) ,
42678	 => std_logic_vector(to_unsigned(115,8) ,
42679	 => std_logic_vector(to_unsigned(105,8) ,
42680	 => std_logic_vector(to_unsigned(112,8) ,
42681	 => std_logic_vector(to_unsigned(109,8) ,
42682	 => std_logic_vector(to_unsigned(108,8) ,
42683	 => std_logic_vector(to_unsigned(125,8) ,
42684	 => std_logic_vector(to_unsigned(43,8) ,
42685	 => std_logic_vector(to_unsigned(2,8) ,
42686	 => std_logic_vector(to_unsigned(1,8) ,
42687	 => std_logic_vector(to_unsigned(1,8) ,
42688	 => std_logic_vector(to_unsigned(1,8) ,
42689	 => std_logic_vector(to_unsigned(35,8) ,
42690	 => std_logic_vector(to_unsigned(136,8) ,
42691	 => std_logic_vector(to_unsigned(116,8) ,
42692	 => std_logic_vector(to_unsigned(103,8) ,
42693	 => std_logic_vector(to_unsigned(116,8) ,
42694	 => std_logic_vector(to_unsigned(133,8) ,
42695	 => std_logic_vector(to_unsigned(35,8) ,
42696	 => std_logic_vector(to_unsigned(3,8) ,
42697	 => std_logic_vector(to_unsigned(6,8) ,
42698	 => std_logic_vector(to_unsigned(6,8) ,
42699	 => std_logic_vector(to_unsigned(3,8) ,
42700	 => std_logic_vector(to_unsigned(3,8) ,
42701	 => std_logic_vector(to_unsigned(58,8) ,
42702	 => std_logic_vector(to_unsigned(157,8) ,
42703	 => std_logic_vector(to_unsigned(128,8) ,
42704	 => std_logic_vector(to_unsigned(128,8) ,
42705	 => std_logic_vector(to_unsigned(131,8) ,
42706	 => std_logic_vector(to_unsigned(139,8) ,
42707	 => std_logic_vector(to_unsigned(130,8) ,
42708	 => std_logic_vector(to_unsigned(127,8) ,
42709	 => std_logic_vector(to_unsigned(133,8) ,
42710	 => std_logic_vector(to_unsigned(128,8) ,
42711	 => std_logic_vector(to_unsigned(22,8) ,
42712	 => std_logic_vector(to_unsigned(2,8) ,
42713	 => std_logic_vector(to_unsigned(6,8) ,
42714	 => std_logic_vector(to_unsigned(5,8) ,
42715	 => std_logic_vector(to_unsigned(3,8) ,
42716	 => std_logic_vector(to_unsigned(0,8) ,
42717	 => std_logic_vector(to_unsigned(17,8) ,
42718	 => std_logic_vector(to_unsigned(159,8) ,
42719	 => std_logic_vector(to_unsigned(60,8) ,
42720	 => std_logic_vector(to_unsigned(3,8) ,
42721	 => std_logic_vector(to_unsigned(3,8) ,
42722	 => std_logic_vector(to_unsigned(15,8) ,
42723	 => std_logic_vector(to_unsigned(9,8) ,
42724	 => std_logic_vector(to_unsigned(2,8) ,
42725	 => std_logic_vector(to_unsigned(38,8) ,
42726	 => std_logic_vector(to_unsigned(109,8) ,
42727	 => std_logic_vector(to_unsigned(96,8) ,
42728	 => std_logic_vector(to_unsigned(79,8) ,
42729	 => std_logic_vector(to_unsigned(67,8) ,
42730	 => std_logic_vector(to_unsigned(47,8) ,
42731	 => std_logic_vector(to_unsigned(37,8) ,
42732	 => std_logic_vector(to_unsigned(25,8) ,
42733	 => std_logic_vector(to_unsigned(16,8) ,
42734	 => std_logic_vector(to_unsigned(14,8) ,
42735	 => std_logic_vector(to_unsigned(4,8) ,
42736	 => std_logic_vector(to_unsigned(1,8) ,
42737	 => std_logic_vector(to_unsigned(2,8) ,
42738	 => std_logic_vector(to_unsigned(2,8) ,
42739	 => std_logic_vector(to_unsigned(3,8) ,
42740	 => std_logic_vector(to_unsigned(4,8) ,
42741	 => std_logic_vector(to_unsigned(1,8) ,
42742	 => std_logic_vector(to_unsigned(1,8) ,
42743	 => std_logic_vector(to_unsigned(0,8) ,
42744	 => std_logic_vector(to_unsigned(0,8) ,
42745	 => std_logic_vector(to_unsigned(0,8) ,
42746	 => std_logic_vector(to_unsigned(0,8) ,
42747	 => std_logic_vector(to_unsigned(17,8) ,
42748	 => std_logic_vector(to_unsigned(66,8) ,
42749	 => std_logic_vector(to_unsigned(47,8) ,
42750	 => std_logic_vector(to_unsigned(27,8) ,
42751	 => std_logic_vector(to_unsigned(14,8) ,
42752	 => std_logic_vector(to_unsigned(6,8) ,
42753	 => std_logic_vector(to_unsigned(1,8) ,
42754	 => std_logic_vector(to_unsigned(0,8) ,
42755	 => std_logic_vector(to_unsigned(1,8) ,
42756	 => std_logic_vector(to_unsigned(2,8) ,
42757	 => std_logic_vector(to_unsigned(2,8) ,
42758	 => std_logic_vector(to_unsigned(3,8) ,
42759	 => std_logic_vector(to_unsigned(3,8) ,
42760	 => std_logic_vector(to_unsigned(4,8) ,
42761	 => std_logic_vector(to_unsigned(4,8) ,
42762	 => std_logic_vector(to_unsigned(3,8) ,
42763	 => std_logic_vector(to_unsigned(4,8) ,
42764	 => std_logic_vector(to_unsigned(3,8) ,
42765	 => std_logic_vector(to_unsigned(3,8) ,
42766	 => std_logic_vector(to_unsigned(2,8) ,
42767	 => std_logic_vector(to_unsigned(10,8) ,
42768	 => std_logic_vector(to_unsigned(37,8) ,
42769	 => std_logic_vector(to_unsigned(20,8) ,
42770	 => std_logic_vector(to_unsigned(4,8) ,
42771	 => std_logic_vector(to_unsigned(1,8) ,
42772	 => std_logic_vector(to_unsigned(2,8) ,
42773	 => std_logic_vector(to_unsigned(10,8) ,
42774	 => std_logic_vector(to_unsigned(8,8) ,
42775	 => std_logic_vector(to_unsigned(12,8) ,
42776	 => std_logic_vector(to_unsigned(24,8) ,
42777	 => std_logic_vector(to_unsigned(24,8) ,
42778	 => std_logic_vector(to_unsigned(5,8) ,
42779	 => std_logic_vector(to_unsigned(2,8) ,
42780	 => std_logic_vector(to_unsigned(0,8) ,
42781	 => std_logic_vector(to_unsigned(0,8) ,
42782	 => std_logic_vector(to_unsigned(0,8) ,
42783	 => std_logic_vector(to_unsigned(0,8) ,
42784	 => std_logic_vector(to_unsigned(1,8) ,
42785	 => std_logic_vector(to_unsigned(1,8) ,
42786	 => std_logic_vector(to_unsigned(1,8) ,
42787	 => std_logic_vector(to_unsigned(1,8) ,
42788	 => std_logic_vector(to_unsigned(1,8) ,
42789	 => std_logic_vector(to_unsigned(2,8) ,
42790	 => std_logic_vector(to_unsigned(2,8) ,
42791	 => std_logic_vector(to_unsigned(0,8) ,
42792	 => std_logic_vector(to_unsigned(44,8) ,
42793	 => std_logic_vector(to_unsigned(206,8) ,
42794	 => std_logic_vector(to_unsigned(33,8) ,
42795	 => std_logic_vector(to_unsigned(0,8) ,
42796	 => std_logic_vector(to_unsigned(0,8) ,
42797	 => std_logic_vector(to_unsigned(0,8) ,
42798	 => std_logic_vector(to_unsigned(1,8) ,
42799	 => std_logic_vector(to_unsigned(3,8) ,
42800	 => std_logic_vector(to_unsigned(5,8) ,
42801	 => std_logic_vector(to_unsigned(6,8) ,
42802	 => std_logic_vector(to_unsigned(2,8) ,
42803	 => std_logic_vector(to_unsigned(3,8) ,
42804	 => std_logic_vector(to_unsigned(3,8) ,
42805	 => std_logic_vector(to_unsigned(2,8) ,
42806	 => std_logic_vector(to_unsigned(2,8) ,
42807	 => std_logic_vector(to_unsigned(1,8) ,
42808	 => std_logic_vector(to_unsigned(8,8) ,
42809	 => std_logic_vector(to_unsigned(10,8) ,
42810	 => std_logic_vector(to_unsigned(3,8) ,
42811	 => std_logic_vector(to_unsigned(1,8) ,
42812	 => std_logic_vector(to_unsigned(1,8) ,
42813	 => std_logic_vector(to_unsigned(1,8) ,
42814	 => std_logic_vector(to_unsigned(1,8) ,
42815	 => std_logic_vector(to_unsigned(1,8) ,
42816	 => std_logic_vector(to_unsigned(2,8) ,
42817	 => std_logic_vector(to_unsigned(1,8) ,
42818	 => std_logic_vector(to_unsigned(3,8) ,
42819	 => std_logic_vector(to_unsigned(3,8) ,
42820	 => std_logic_vector(to_unsigned(3,8) ,
42821	 => std_logic_vector(to_unsigned(2,8) ,
42822	 => std_logic_vector(to_unsigned(0,8) ,
42823	 => std_logic_vector(to_unsigned(0,8) ,
42824	 => std_logic_vector(to_unsigned(0,8) ,
42825	 => std_logic_vector(to_unsigned(6,8) ,
42826	 => std_logic_vector(to_unsigned(51,8) ,
42827	 => std_logic_vector(to_unsigned(49,8) ,
42828	 => std_logic_vector(to_unsigned(41,8) ,
42829	 => std_logic_vector(to_unsigned(24,8) ,
42830	 => std_logic_vector(to_unsigned(18,8) ,
42831	 => std_logic_vector(to_unsigned(9,8) ,
42832	 => std_logic_vector(to_unsigned(4,8) ,
42833	 => std_logic_vector(to_unsigned(8,8) ,
42834	 => std_logic_vector(to_unsigned(31,8) ,
42835	 => std_logic_vector(to_unsigned(15,8) ,
42836	 => std_logic_vector(to_unsigned(0,8) ,
42837	 => std_logic_vector(to_unsigned(1,8) ,
42838	 => std_logic_vector(to_unsigned(1,8) ,
42839	 => std_logic_vector(to_unsigned(1,8) ,
42840	 => std_logic_vector(to_unsigned(1,8) ,
42841	 => std_logic_vector(to_unsigned(1,8) ,
42842	 => std_logic_vector(to_unsigned(1,8) ,
42843	 => std_logic_vector(to_unsigned(2,8) ,
42844	 => std_logic_vector(to_unsigned(1,8) ,
42845	 => std_logic_vector(to_unsigned(2,8) ,
42846	 => std_logic_vector(to_unsigned(6,8) ,
42847	 => std_logic_vector(to_unsigned(2,8) ,
42848	 => std_logic_vector(to_unsigned(2,8) ,
42849	 => std_logic_vector(to_unsigned(3,8) ,
42850	 => std_logic_vector(to_unsigned(1,8) ,
42851	 => std_logic_vector(to_unsigned(1,8) ,
42852	 => std_logic_vector(to_unsigned(1,8) ,
42853	 => std_logic_vector(to_unsigned(1,8) ,
42854	 => std_logic_vector(to_unsigned(1,8) ,
42855	 => std_logic_vector(to_unsigned(1,8) ,
42856	 => std_logic_vector(to_unsigned(1,8) ,
42857	 => std_logic_vector(to_unsigned(1,8) ,
42858	 => std_logic_vector(to_unsigned(1,8) ,
42859	 => std_logic_vector(to_unsigned(2,8) ,
42860	 => std_logic_vector(to_unsigned(1,8) ,
42861	 => std_logic_vector(to_unsigned(1,8) ,
42862	 => std_logic_vector(to_unsigned(2,8) ,
42863	 => std_logic_vector(to_unsigned(2,8) ,
42864	 => std_logic_vector(to_unsigned(2,8) ,
42865	 => std_logic_vector(to_unsigned(1,8) ,
42866	 => std_logic_vector(to_unsigned(1,8) ,
42867	 => std_logic_vector(to_unsigned(1,8) ,
42868	 => std_logic_vector(to_unsigned(2,8) ,
42869	 => std_logic_vector(to_unsigned(1,8) ,
42870	 => std_logic_vector(to_unsigned(2,8) ,
42871	 => std_logic_vector(to_unsigned(1,8) ,
42872	 => std_logic_vector(to_unsigned(2,8) ,
42873	 => std_logic_vector(to_unsigned(2,8) ,
42874	 => std_logic_vector(to_unsigned(2,8) ,
42875	 => std_logic_vector(to_unsigned(3,8) ,
42876	 => std_logic_vector(to_unsigned(1,8) ,
42877	 => std_logic_vector(to_unsigned(1,8) ,
42878	 => std_logic_vector(to_unsigned(2,8) ,
42879	 => std_logic_vector(to_unsigned(2,8) ,
42880	 => std_logic_vector(to_unsigned(2,8) ,
42881	 => std_logic_vector(to_unsigned(90,8) ,
42882	 => std_logic_vector(to_unsigned(79,8) ,
42883	 => std_logic_vector(to_unsigned(84,8) ,
42884	 => std_logic_vector(to_unsigned(85,8) ,
42885	 => std_logic_vector(to_unsigned(87,8) ,
42886	 => std_logic_vector(to_unsigned(87,8) ,
42887	 => std_logic_vector(to_unsigned(93,8) ,
42888	 => std_logic_vector(to_unsigned(69,8) ,
42889	 => std_logic_vector(to_unsigned(52,8) ,
42890	 => std_logic_vector(to_unsigned(57,8) ,
42891	 => std_logic_vector(to_unsigned(52,8) ,
42892	 => std_logic_vector(to_unsigned(58,8) ,
42893	 => std_logic_vector(to_unsigned(61,8) ,
42894	 => std_logic_vector(to_unsigned(80,8) ,
42895	 => std_logic_vector(to_unsigned(95,8) ,
42896	 => std_logic_vector(to_unsigned(99,8) ,
42897	 => std_logic_vector(to_unsigned(97,8) ,
42898	 => std_logic_vector(to_unsigned(74,8) ,
42899	 => std_logic_vector(to_unsigned(100,8) ,
42900	 => std_logic_vector(to_unsigned(139,8) ,
42901	 => std_logic_vector(to_unsigned(133,8) ,
42902	 => std_logic_vector(to_unsigned(136,8) ,
42903	 => std_logic_vector(to_unsigned(131,8) ,
42904	 => std_logic_vector(to_unsigned(131,8) ,
42905	 => std_logic_vector(to_unsigned(146,8) ,
42906	 => std_logic_vector(to_unsigned(138,8) ,
42907	 => std_logic_vector(to_unsigned(152,8) ,
42908	 => std_logic_vector(to_unsigned(142,8) ,
42909	 => std_logic_vector(to_unsigned(112,8) ,
42910	 => std_logic_vector(to_unsigned(133,8) ,
42911	 => std_logic_vector(to_unsigned(149,8) ,
42912	 => std_logic_vector(to_unsigned(156,8) ,
42913	 => std_logic_vector(to_unsigned(161,8) ,
42914	 => std_logic_vector(to_unsigned(147,8) ,
42915	 => std_logic_vector(to_unsigned(144,8) ,
42916	 => std_logic_vector(to_unsigned(147,8) ,
42917	 => std_logic_vector(to_unsigned(151,8) ,
42918	 => std_logic_vector(to_unsigned(152,8) ,
42919	 => std_logic_vector(to_unsigned(156,8) ,
42920	 => std_logic_vector(to_unsigned(138,8) ,
42921	 => std_logic_vector(to_unsigned(105,8) ,
42922	 => std_logic_vector(to_unsigned(125,8) ,
42923	 => std_logic_vector(to_unsigned(105,8) ,
42924	 => std_logic_vector(to_unsigned(119,8) ,
42925	 => std_logic_vector(to_unsigned(119,8) ,
42926	 => std_logic_vector(to_unsigned(116,8) ,
42927	 => std_logic_vector(to_unsigned(133,8) ,
42928	 => std_logic_vector(to_unsigned(134,8) ,
42929	 => std_logic_vector(to_unsigned(154,8) ,
42930	 => std_logic_vector(to_unsigned(146,8) ,
42931	 => std_logic_vector(to_unsigned(141,8) ,
42932	 => std_logic_vector(to_unsigned(156,8) ,
42933	 => std_logic_vector(to_unsigned(146,8) ,
42934	 => std_logic_vector(to_unsigned(121,8) ,
42935	 => std_logic_vector(to_unsigned(111,8) ,
42936	 => std_logic_vector(to_unsigned(111,8) ,
42937	 => std_logic_vector(to_unsigned(118,8) ,
42938	 => std_logic_vector(to_unsigned(118,8) ,
42939	 => std_logic_vector(to_unsigned(116,8) ,
42940	 => std_logic_vector(to_unsigned(119,8) ,
42941	 => std_logic_vector(to_unsigned(124,8) ,
42942	 => std_logic_vector(to_unsigned(118,8) ,
42943	 => std_logic_vector(to_unsigned(108,8) ,
42944	 => std_logic_vector(to_unsigned(112,8) ,
42945	 => std_logic_vector(to_unsigned(105,8) ,
42946	 => std_logic_vector(to_unsigned(100,8) ,
42947	 => std_logic_vector(to_unsigned(111,8) ,
42948	 => std_logic_vector(to_unsigned(100,8) ,
42949	 => std_logic_vector(to_unsigned(90,8) ,
42950	 => std_logic_vector(to_unsigned(101,8) ,
42951	 => std_logic_vector(to_unsigned(97,8) ,
42952	 => std_logic_vector(to_unsigned(86,8) ,
42953	 => std_logic_vector(to_unsigned(78,8) ,
42954	 => std_logic_vector(to_unsigned(18,8) ,
42955	 => std_logic_vector(to_unsigned(4,8) ,
42956	 => std_logic_vector(to_unsigned(14,8) ,
42957	 => std_logic_vector(to_unsigned(17,8) ,
42958	 => std_logic_vector(to_unsigned(8,8) ,
42959	 => std_logic_vector(to_unsigned(2,8) ,
42960	 => std_logic_vector(to_unsigned(9,8) ,
42961	 => std_logic_vector(to_unsigned(70,8) ,
42962	 => std_logic_vector(to_unsigned(125,8) ,
42963	 => std_logic_vector(to_unsigned(121,8) ,
42964	 => std_logic_vector(to_unsigned(114,8) ,
42965	 => std_logic_vector(to_unsigned(112,8) ,
42966	 => std_logic_vector(to_unsigned(109,8) ,
42967	 => std_logic_vector(to_unsigned(103,8) ,
42968	 => std_logic_vector(to_unsigned(87,8) ,
42969	 => std_logic_vector(to_unsigned(85,8) ,
42970	 => std_logic_vector(to_unsigned(86,8) ,
42971	 => std_logic_vector(to_unsigned(99,8) ,
42972	 => std_logic_vector(to_unsigned(60,8) ,
42973	 => std_logic_vector(to_unsigned(3,8) ,
42974	 => std_logic_vector(to_unsigned(7,8) ,
42975	 => std_logic_vector(to_unsigned(80,8) ,
42976	 => std_logic_vector(to_unsigned(51,8) ,
42977	 => std_logic_vector(to_unsigned(38,8) ,
42978	 => std_logic_vector(to_unsigned(48,8) ,
42979	 => std_logic_vector(to_unsigned(12,8) ,
42980	 => std_logic_vector(to_unsigned(2,8) ,
42981	 => std_logic_vector(to_unsigned(5,8) ,
42982	 => std_logic_vector(to_unsigned(7,8) ,
42983	 => std_logic_vector(to_unsigned(10,8) ,
42984	 => std_logic_vector(to_unsigned(5,8) ,
42985	 => std_logic_vector(to_unsigned(0,8) ,
42986	 => std_logic_vector(to_unsigned(2,8) ,
42987	 => std_logic_vector(to_unsigned(21,8) ,
42988	 => std_logic_vector(to_unsigned(34,8) ,
42989	 => std_logic_vector(to_unsigned(13,8) ,
42990	 => std_logic_vector(to_unsigned(38,8) ,
42991	 => std_logic_vector(to_unsigned(121,8) ,
42992	 => std_logic_vector(to_unsigned(133,8) ,
42993	 => std_logic_vector(to_unsigned(100,8) ,
42994	 => std_logic_vector(to_unsigned(105,8) ,
42995	 => std_logic_vector(to_unsigned(107,8) ,
42996	 => std_logic_vector(to_unsigned(118,8) ,
42997	 => std_logic_vector(to_unsigned(115,8) ,
42998	 => std_logic_vector(to_unsigned(109,8) ,
42999	 => std_logic_vector(to_unsigned(104,8) ,
43000	 => std_logic_vector(to_unsigned(104,8) ,
43001	 => std_logic_vector(to_unsigned(105,8) ,
43002	 => std_logic_vector(to_unsigned(103,8) ,
43003	 => std_logic_vector(to_unsigned(115,8) ,
43004	 => std_logic_vector(to_unsigned(37,8) ,
43005	 => std_logic_vector(to_unsigned(3,8) ,
43006	 => std_logic_vector(to_unsigned(4,8) ,
43007	 => std_logic_vector(to_unsigned(2,8) ,
43008	 => std_logic_vector(to_unsigned(2,8) ,
43009	 => std_logic_vector(to_unsigned(30,8) ,
43010	 => std_logic_vector(to_unsigned(128,8) ,
43011	 => std_logic_vector(to_unsigned(122,8) ,
43012	 => std_logic_vector(to_unsigned(115,8) ,
43013	 => std_logic_vector(to_unsigned(118,8) ,
43014	 => std_logic_vector(to_unsigned(125,8) ,
43015	 => std_logic_vector(to_unsigned(22,8) ,
43016	 => std_logic_vector(to_unsigned(1,8) ,
43017	 => std_logic_vector(to_unsigned(5,8) ,
43018	 => std_logic_vector(to_unsigned(3,8) ,
43019	 => std_logic_vector(to_unsigned(4,8) ,
43020	 => std_logic_vector(to_unsigned(43,8) ,
43021	 => std_logic_vector(to_unsigned(125,8) ,
43022	 => std_logic_vector(to_unsigned(124,8) ,
43023	 => std_logic_vector(to_unsigned(116,8) ,
43024	 => std_logic_vector(to_unsigned(116,8) ,
43025	 => std_logic_vector(to_unsigned(121,8) ,
43026	 => std_logic_vector(to_unsigned(116,8) ,
43027	 => std_logic_vector(to_unsigned(125,8) ,
43028	 => std_logic_vector(to_unsigned(133,8) ,
43029	 => std_logic_vector(to_unsigned(146,8) ,
43030	 => std_logic_vector(to_unsigned(118,8) ,
43031	 => std_logic_vector(to_unsigned(11,8) ,
43032	 => std_logic_vector(to_unsigned(3,8) ,
43033	 => std_logic_vector(to_unsigned(6,8) ,
43034	 => std_logic_vector(to_unsigned(7,8) ,
43035	 => std_logic_vector(to_unsigned(6,8) ,
43036	 => std_logic_vector(to_unsigned(0,8) ,
43037	 => std_logic_vector(to_unsigned(16,8) ,
43038	 => std_logic_vector(to_unsigned(101,8) ,
43039	 => std_logic_vector(to_unsigned(10,8) ,
43040	 => std_logic_vector(to_unsigned(4,8) ,
43041	 => std_logic_vector(to_unsigned(10,8) ,
43042	 => std_logic_vector(to_unsigned(12,8) ,
43043	 => std_logic_vector(to_unsigned(3,8) ,
43044	 => std_logic_vector(to_unsigned(5,8) ,
43045	 => std_logic_vector(to_unsigned(95,8) ,
43046	 => std_logic_vector(to_unsigned(139,8) ,
43047	 => std_logic_vector(to_unsigned(124,8) ,
43048	 => std_logic_vector(to_unsigned(127,8) ,
43049	 => std_logic_vector(to_unsigned(133,8) ,
43050	 => std_logic_vector(to_unsigned(121,8) ,
43051	 => std_logic_vector(to_unsigned(114,8) ,
43052	 => std_logic_vector(to_unsigned(118,8) ,
43053	 => std_logic_vector(to_unsigned(115,8) ,
43054	 => std_logic_vector(to_unsigned(99,8) ,
43055	 => std_logic_vector(to_unsigned(76,8) ,
43056	 => std_logic_vector(to_unsigned(48,8) ,
43057	 => std_logic_vector(to_unsigned(3,8) ,
43058	 => std_logic_vector(to_unsigned(1,8) ,
43059	 => std_logic_vector(to_unsigned(6,8) ,
43060	 => std_logic_vector(to_unsigned(5,8) ,
43061	 => std_logic_vector(to_unsigned(2,8) ,
43062	 => std_logic_vector(to_unsigned(2,8) ,
43063	 => std_logic_vector(to_unsigned(4,8) ,
43064	 => std_logic_vector(to_unsigned(5,8) ,
43065	 => std_logic_vector(to_unsigned(2,8) ,
43066	 => std_logic_vector(to_unsigned(2,8) ,
43067	 => std_logic_vector(to_unsigned(13,8) ,
43068	 => std_logic_vector(to_unsigned(42,8) ,
43069	 => std_logic_vector(to_unsigned(41,8) ,
43070	 => std_logic_vector(to_unsigned(33,8) ,
43071	 => std_logic_vector(to_unsigned(6,8) ,
43072	 => std_logic_vector(to_unsigned(0,8) ,
43073	 => std_logic_vector(to_unsigned(0,8) ,
43074	 => std_logic_vector(to_unsigned(0,8) ,
43075	 => std_logic_vector(to_unsigned(0,8) ,
43076	 => std_logic_vector(to_unsigned(1,8) ,
43077	 => std_logic_vector(to_unsigned(1,8) ,
43078	 => std_logic_vector(to_unsigned(1,8) ,
43079	 => std_logic_vector(to_unsigned(2,8) ,
43080	 => std_logic_vector(to_unsigned(2,8) ,
43081	 => std_logic_vector(to_unsigned(2,8) ,
43082	 => std_logic_vector(to_unsigned(4,8) ,
43083	 => std_logic_vector(to_unsigned(4,8) ,
43084	 => std_logic_vector(to_unsigned(4,8) ,
43085	 => std_logic_vector(to_unsigned(5,8) ,
43086	 => std_logic_vector(to_unsigned(2,8) ,
43087	 => std_logic_vector(to_unsigned(13,8) ,
43088	 => std_logic_vector(to_unsigned(32,8) ,
43089	 => std_logic_vector(to_unsigned(12,8) ,
43090	 => std_logic_vector(to_unsigned(4,8) ,
43091	 => std_logic_vector(to_unsigned(2,8) ,
43092	 => std_logic_vector(to_unsigned(0,8) ,
43093	 => std_logic_vector(to_unsigned(0,8) ,
43094	 => std_logic_vector(to_unsigned(0,8) ,
43095	 => std_logic_vector(to_unsigned(0,8) ,
43096	 => std_logic_vector(to_unsigned(1,8) ,
43097	 => std_logic_vector(to_unsigned(1,8) ,
43098	 => std_logic_vector(to_unsigned(1,8) ,
43099	 => std_logic_vector(to_unsigned(1,8) ,
43100	 => std_logic_vector(to_unsigned(1,8) ,
43101	 => std_logic_vector(to_unsigned(1,8) ,
43102	 => std_logic_vector(to_unsigned(0,8) ,
43103	 => std_logic_vector(to_unsigned(1,8) ,
43104	 => std_logic_vector(to_unsigned(1,8) ,
43105	 => std_logic_vector(to_unsigned(1,8) ,
43106	 => std_logic_vector(to_unsigned(1,8) ,
43107	 => std_logic_vector(to_unsigned(2,8) ,
43108	 => std_logic_vector(to_unsigned(1,8) ,
43109	 => std_logic_vector(to_unsigned(1,8) ,
43110	 => std_logic_vector(to_unsigned(2,8) ,
43111	 => std_logic_vector(to_unsigned(0,8) ,
43112	 => std_logic_vector(to_unsigned(18,8) ,
43113	 => std_logic_vector(to_unsigned(78,8) ,
43114	 => std_logic_vector(to_unsigned(2,8) ,
43115	 => std_logic_vector(to_unsigned(0,8) ,
43116	 => std_logic_vector(to_unsigned(0,8) ,
43117	 => std_logic_vector(to_unsigned(0,8) ,
43118	 => std_logic_vector(to_unsigned(1,8) ,
43119	 => std_logic_vector(to_unsigned(3,8) ,
43120	 => std_logic_vector(to_unsigned(3,8) ,
43121	 => std_logic_vector(to_unsigned(4,8) ,
43122	 => std_logic_vector(to_unsigned(3,8) ,
43123	 => std_logic_vector(to_unsigned(2,8) ,
43124	 => std_logic_vector(to_unsigned(3,8) ,
43125	 => std_logic_vector(to_unsigned(2,8) ,
43126	 => std_logic_vector(to_unsigned(2,8) ,
43127	 => std_logic_vector(to_unsigned(2,8) ,
43128	 => std_logic_vector(to_unsigned(9,8) ,
43129	 => std_logic_vector(to_unsigned(10,8) ,
43130	 => std_logic_vector(to_unsigned(2,8) ,
43131	 => std_logic_vector(to_unsigned(1,8) ,
43132	 => std_logic_vector(to_unsigned(1,8) ,
43133	 => std_logic_vector(to_unsigned(2,8) ,
43134	 => std_logic_vector(to_unsigned(1,8) ,
43135	 => std_logic_vector(to_unsigned(1,8) ,
43136	 => std_logic_vector(to_unsigned(2,8) ,
43137	 => std_logic_vector(to_unsigned(3,8) ,
43138	 => std_logic_vector(to_unsigned(3,8) ,
43139	 => std_logic_vector(to_unsigned(3,8) ,
43140	 => std_logic_vector(to_unsigned(3,8) ,
43141	 => std_logic_vector(to_unsigned(2,8) ,
43142	 => std_logic_vector(to_unsigned(0,8) ,
43143	 => std_logic_vector(to_unsigned(0,8) ,
43144	 => std_logic_vector(to_unsigned(0,8) ,
43145	 => std_logic_vector(to_unsigned(9,8) ,
43146	 => std_logic_vector(to_unsigned(39,8) ,
43147	 => std_logic_vector(to_unsigned(43,8) ,
43148	 => std_logic_vector(to_unsigned(38,8) ,
43149	 => std_logic_vector(to_unsigned(30,8) ,
43150	 => std_logic_vector(to_unsigned(22,8) ,
43151	 => std_logic_vector(to_unsigned(12,8) ,
43152	 => std_logic_vector(to_unsigned(5,8) ,
43153	 => std_logic_vector(to_unsigned(8,8) ,
43154	 => std_logic_vector(to_unsigned(22,8) ,
43155	 => std_logic_vector(to_unsigned(23,8) ,
43156	 => std_logic_vector(to_unsigned(1,8) ,
43157	 => std_logic_vector(to_unsigned(1,8) ,
43158	 => std_logic_vector(to_unsigned(2,8) ,
43159	 => std_logic_vector(to_unsigned(1,8) ,
43160	 => std_logic_vector(to_unsigned(1,8) ,
43161	 => std_logic_vector(to_unsigned(1,8) ,
43162	 => std_logic_vector(to_unsigned(1,8) ,
43163	 => std_logic_vector(to_unsigned(2,8) ,
43164	 => std_logic_vector(to_unsigned(2,8) ,
43165	 => std_logic_vector(to_unsigned(5,8) ,
43166	 => std_logic_vector(to_unsigned(7,8) ,
43167	 => std_logic_vector(to_unsigned(4,8) ,
43168	 => std_logic_vector(to_unsigned(2,8) ,
43169	 => std_logic_vector(to_unsigned(3,8) ,
43170	 => std_logic_vector(to_unsigned(3,8) ,
43171	 => std_logic_vector(to_unsigned(3,8) ,
43172	 => std_logic_vector(to_unsigned(1,8) ,
43173	 => std_logic_vector(to_unsigned(0,8) ,
43174	 => std_logic_vector(to_unsigned(1,8) ,
43175	 => std_logic_vector(to_unsigned(1,8) ,
43176	 => std_logic_vector(to_unsigned(1,8) ,
43177	 => std_logic_vector(to_unsigned(1,8) ,
43178	 => std_logic_vector(to_unsigned(1,8) ,
43179	 => std_logic_vector(to_unsigned(1,8) ,
43180	 => std_logic_vector(to_unsigned(1,8) ,
43181	 => std_logic_vector(to_unsigned(1,8) ,
43182	 => std_logic_vector(to_unsigned(2,8) ,
43183	 => std_logic_vector(to_unsigned(1,8) ,
43184	 => std_logic_vector(to_unsigned(2,8) ,
43185	 => std_logic_vector(to_unsigned(2,8) ,
43186	 => std_logic_vector(to_unsigned(2,8) ,
43187	 => std_logic_vector(to_unsigned(2,8) ,
43188	 => std_logic_vector(to_unsigned(2,8) ,
43189	 => std_logic_vector(to_unsigned(2,8) ,
43190	 => std_logic_vector(to_unsigned(3,8) ,
43191	 => std_logic_vector(to_unsigned(2,8) ,
43192	 => std_logic_vector(to_unsigned(2,8) ,
43193	 => std_logic_vector(to_unsigned(2,8) ,
43194	 => std_logic_vector(to_unsigned(2,8) ,
43195	 => std_logic_vector(to_unsigned(3,8) ,
43196	 => std_logic_vector(to_unsigned(2,8) ,
43197	 => std_logic_vector(to_unsigned(1,8) ,
43198	 => std_logic_vector(to_unsigned(2,8) ,
43199	 => std_logic_vector(to_unsigned(2,8) ,
43200	 => std_logic_vector(to_unsigned(2,8) ,
43201	 => std_logic_vector(to_unsigned(81,8) ,
43202	 => std_logic_vector(to_unsigned(78,8) ,
43203	 => std_logic_vector(to_unsigned(84,8) ,
43204	 => std_logic_vector(to_unsigned(90,8) ,
43205	 => std_logic_vector(to_unsigned(82,8) ,
43206	 => std_logic_vector(to_unsigned(73,8) ,
43207	 => std_logic_vector(to_unsigned(81,8) ,
43208	 => std_logic_vector(to_unsigned(61,8) ,
43209	 => std_logic_vector(to_unsigned(53,8) ,
43210	 => std_logic_vector(to_unsigned(53,8) ,
43211	 => std_logic_vector(to_unsigned(56,8) ,
43212	 => std_logic_vector(to_unsigned(56,8) ,
43213	 => std_logic_vector(to_unsigned(58,8) ,
43214	 => std_logic_vector(to_unsigned(105,8) ,
43215	 => std_logic_vector(to_unsigned(133,8) ,
43216	 => std_logic_vector(to_unsigned(118,8) ,
43217	 => std_logic_vector(to_unsigned(111,8) ,
43218	 => std_logic_vector(to_unsigned(119,8) ,
43219	 => std_logic_vector(to_unsigned(130,8) ,
43220	 => std_logic_vector(to_unsigned(133,8) ,
43221	 => std_logic_vector(to_unsigned(138,8) ,
43222	 => std_logic_vector(to_unsigned(138,8) ,
43223	 => std_logic_vector(to_unsigned(131,8) ,
43224	 => std_logic_vector(to_unsigned(125,8) ,
43225	 => std_logic_vector(to_unsigned(134,8) ,
43226	 => std_logic_vector(to_unsigned(138,8) ,
43227	 => std_logic_vector(to_unsigned(133,8) ,
43228	 => std_logic_vector(to_unsigned(131,8) ,
43229	 => std_logic_vector(to_unsigned(112,8) ,
43230	 => std_logic_vector(to_unsigned(130,8) ,
43231	 => std_logic_vector(to_unsigned(139,8) ,
43232	 => std_logic_vector(to_unsigned(130,8) ,
43233	 => std_logic_vector(to_unsigned(133,8) ,
43234	 => std_logic_vector(to_unsigned(138,8) ,
43235	 => std_logic_vector(to_unsigned(144,8) ,
43236	 => std_logic_vector(to_unsigned(146,8) ,
43237	 => std_logic_vector(to_unsigned(147,8) ,
43238	 => std_logic_vector(to_unsigned(147,8) ,
43239	 => std_logic_vector(to_unsigned(161,8) ,
43240	 => std_logic_vector(to_unsigned(144,8) ,
43241	 => std_logic_vector(to_unsigned(99,8) ,
43242	 => std_logic_vector(to_unsigned(119,8) ,
43243	 => std_logic_vector(to_unsigned(99,8) ,
43244	 => std_logic_vector(to_unsigned(116,8) ,
43245	 => std_logic_vector(to_unsigned(122,8) ,
43246	 => std_logic_vector(to_unsigned(108,8) ,
43247	 => std_logic_vector(to_unsigned(121,8) ,
43248	 => std_logic_vector(to_unsigned(128,8) ,
43249	 => std_logic_vector(to_unsigned(144,8) ,
43250	 => std_logic_vector(to_unsigned(134,8) ,
43251	 => std_logic_vector(to_unsigned(131,8) ,
43252	 => std_logic_vector(to_unsigned(152,8) ,
43253	 => std_logic_vector(to_unsigned(146,8) ,
43254	 => std_logic_vector(to_unsigned(121,8) ,
43255	 => std_logic_vector(to_unsigned(109,8) ,
43256	 => std_logic_vector(to_unsigned(100,8) ,
43257	 => std_logic_vector(to_unsigned(105,8) ,
43258	 => std_logic_vector(to_unsigned(115,8) ,
43259	 => std_logic_vector(to_unsigned(115,8) ,
43260	 => std_logic_vector(to_unsigned(115,8) ,
43261	 => std_logic_vector(to_unsigned(112,8) ,
43262	 => std_logic_vector(to_unsigned(109,8) ,
43263	 => std_logic_vector(to_unsigned(111,8) ,
43264	 => std_logic_vector(to_unsigned(114,8) ,
43265	 => std_logic_vector(to_unsigned(105,8) ,
43266	 => std_logic_vector(to_unsigned(105,8) ,
43267	 => std_logic_vector(to_unsigned(104,8) ,
43268	 => std_logic_vector(to_unsigned(100,8) ,
43269	 => std_logic_vector(to_unsigned(96,8) ,
43270	 => std_logic_vector(to_unsigned(95,8) ,
43271	 => std_logic_vector(to_unsigned(97,8) ,
43272	 => std_logic_vector(to_unsigned(91,8) ,
43273	 => std_logic_vector(to_unsigned(24,8) ,
43274	 => std_logic_vector(to_unsigned(6,8) ,
43275	 => std_logic_vector(to_unsigned(8,8) ,
43276	 => std_logic_vector(to_unsigned(12,8) ,
43277	 => std_logic_vector(to_unsigned(6,8) ,
43278	 => std_logic_vector(to_unsigned(1,8) ,
43279	 => std_logic_vector(to_unsigned(3,8) ,
43280	 => std_logic_vector(to_unsigned(66,8) ,
43281	 => std_logic_vector(to_unsigned(139,8) ,
43282	 => std_logic_vector(to_unsigned(99,8) ,
43283	 => std_logic_vector(to_unsigned(99,8) ,
43284	 => std_logic_vector(to_unsigned(103,8) ,
43285	 => std_logic_vector(to_unsigned(107,8) ,
43286	 => std_logic_vector(to_unsigned(111,8) ,
43287	 => std_logic_vector(to_unsigned(99,8) ,
43288	 => std_logic_vector(to_unsigned(82,8) ,
43289	 => std_logic_vector(to_unsigned(73,8) ,
43290	 => std_logic_vector(to_unsigned(96,8) ,
43291	 => std_logic_vector(to_unsigned(68,8) ,
43292	 => std_logic_vector(to_unsigned(16,8) ,
43293	 => std_logic_vector(to_unsigned(11,8) ,
43294	 => std_logic_vector(to_unsigned(23,8) ,
43295	 => std_logic_vector(to_unsigned(46,8) ,
43296	 => std_logic_vector(to_unsigned(77,8) ,
43297	 => std_logic_vector(to_unsigned(53,8) ,
43298	 => std_logic_vector(to_unsigned(14,8) ,
43299	 => std_logic_vector(to_unsigned(5,8) ,
43300	 => std_logic_vector(to_unsigned(4,8) ,
43301	 => std_logic_vector(to_unsigned(4,8) ,
43302	 => std_logic_vector(to_unsigned(8,8) ,
43303	 => std_logic_vector(to_unsigned(7,8) ,
43304	 => std_logic_vector(to_unsigned(3,8) ,
43305	 => std_logic_vector(to_unsigned(2,8) ,
43306	 => std_logic_vector(to_unsigned(35,8) ,
43307	 => std_logic_vector(to_unsigned(96,8) ,
43308	 => std_logic_vector(to_unsigned(96,8) ,
43309	 => std_logic_vector(to_unsigned(97,8) ,
43310	 => std_logic_vector(to_unsigned(101,8) ,
43311	 => std_logic_vector(to_unsigned(103,8) ,
43312	 => std_logic_vector(to_unsigned(107,8) ,
43313	 => std_logic_vector(to_unsigned(114,8) ,
43314	 => std_logic_vector(to_unsigned(97,8) ,
43315	 => std_logic_vector(to_unsigned(101,8) ,
43316	 => std_logic_vector(to_unsigned(100,8) ,
43317	 => std_logic_vector(to_unsigned(105,8) ,
43318	 => std_logic_vector(to_unsigned(111,8) ,
43319	 => std_logic_vector(to_unsigned(107,8) ,
43320	 => std_logic_vector(to_unsigned(111,8) ,
43321	 => std_logic_vector(to_unsigned(115,8) ,
43322	 => std_logic_vector(to_unsigned(101,8) ,
43323	 => std_logic_vector(to_unsigned(109,8) ,
43324	 => std_logic_vector(to_unsigned(37,8) ,
43325	 => std_logic_vector(to_unsigned(5,8) ,
43326	 => std_logic_vector(to_unsigned(4,8) ,
43327	 => std_logic_vector(to_unsigned(2,8) ,
43328	 => std_logic_vector(to_unsigned(1,8) ,
43329	 => std_logic_vector(to_unsigned(32,8) ,
43330	 => std_logic_vector(to_unsigned(131,8) ,
43331	 => std_logic_vector(to_unsigned(133,8) ,
43332	 => std_logic_vector(to_unsigned(125,8) ,
43333	 => std_logic_vector(to_unsigned(108,8) ,
43334	 => std_logic_vector(to_unsigned(100,8) ,
43335	 => std_logic_vector(to_unsigned(56,8) ,
43336	 => std_logic_vector(to_unsigned(18,8) ,
43337	 => std_logic_vector(to_unsigned(16,8) ,
43338	 => std_logic_vector(to_unsigned(23,8) ,
43339	 => std_logic_vector(to_unsigned(51,8) ,
43340	 => std_logic_vector(to_unsigned(105,8) ,
43341	 => std_logic_vector(to_unsigned(112,8) ,
43342	 => std_logic_vector(to_unsigned(96,8) ,
43343	 => std_logic_vector(to_unsigned(103,8) ,
43344	 => std_logic_vector(to_unsigned(114,8) ,
43345	 => std_logic_vector(to_unsigned(112,8) ,
43346	 => std_logic_vector(to_unsigned(92,8) ,
43347	 => std_logic_vector(to_unsigned(108,8) ,
43348	 => std_logic_vector(to_unsigned(124,8) ,
43349	 => std_logic_vector(to_unsigned(141,8) ,
43350	 => std_logic_vector(to_unsigned(77,8) ,
43351	 => std_logic_vector(to_unsigned(5,8) ,
43352	 => std_logic_vector(to_unsigned(6,8) ,
43353	 => std_logic_vector(to_unsigned(10,8) ,
43354	 => std_logic_vector(to_unsigned(5,8) ,
43355	 => std_logic_vector(to_unsigned(1,8) ,
43356	 => std_logic_vector(to_unsigned(3,8) ,
43357	 => std_logic_vector(to_unsigned(79,8) ,
43358	 => std_logic_vector(to_unsigned(66,8) ,
43359	 => std_logic_vector(to_unsigned(3,8) ,
43360	 => std_logic_vector(to_unsigned(9,8) ,
43361	 => std_logic_vector(to_unsigned(12,8) ,
43362	 => std_logic_vector(to_unsigned(12,8) ,
43363	 => std_logic_vector(to_unsigned(4,8) ,
43364	 => std_logic_vector(to_unsigned(4,8) ,
43365	 => std_logic_vector(to_unsigned(84,8) ,
43366	 => std_logic_vector(to_unsigned(105,8) ,
43367	 => std_logic_vector(to_unsigned(104,8) ,
43368	 => std_logic_vector(to_unsigned(108,8) ,
43369	 => std_logic_vector(to_unsigned(101,8) ,
43370	 => std_logic_vector(to_unsigned(112,8) ,
43371	 => std_logic_vector(to_unsigned(107,8) ,
43372	 => std_logic_vector(to_unsigned(100,8) ,
43373	 => std_logic_vector(to_unsigned(103,8) ,
43374	 => std_logic_vector(to_unsigned(100,8) ,
43375	 => std_logic_vector(to_unsigned(97,8) ,
43376	 => std_logic_vector(to_unsigned(87,8) ,
43377	 => std_logic_vector(to_unsigned(4,8) ,
43378	 => std_logic_vector(to_unsigned(2,8) ,
43379	 => std_logic_vector(to_unsigned(12,8) ,
43380	 => std_logic_vector(to_unsigned(4,8) ,
43381	 => std_logic_vector(to_unsigned(4,8) ,
43382	 => std_logic_vector(to_unsigned(1,8) ,
43383	 => std_logic_vector(to_unsigned(32,8) ,
43384	 => std_logic_vector(to_unsigned(100,8) ,
43385	 => std_logic_vector(to_unsigned(38,8) ,
43386	 => std_logic_vector(to_unsigned(8,8) ,
43387	 => std_logic_vector(to_unsigned(13,8) ,
43388	 => std_logic_vector(to_unsigned(27,8) ,
43389	 => std_logic_vector(to_unsigned(29,8) ,
43390	 => std_logic_vector(to_unsigned(13,8) ,
43391	 => std_logic_vector(to_unsigned(17,8) ,
43392	 => std_logic_vector(to_unsigned(22,8) ,
43393	 => std_logic_vector(to_unsigned(12,8) ,
43394	 => std_logic_vector(to_unsigned(7,8) ,
43395	 => std_logic_vector(to_unsigned(6,8) ,
43396	 => std_logic_vector(to_unsigned(5,8) ,
43397	 => std_logic_vector(to_unsigned(3,8) ,
43398	 => std_logic_vector(to_unsigned(2,8) ,
43399	 => std_logic_vector(to_unsigned(2,8) ,
43400	 => std_logic_vector(to_unsigned(2,8) ,
43401	 => std_logic_vector(to_unsigned(2,8) ,
43402	 => std_logic_vector(to_unsigned(1,8) ,
43403	 => std_logic_vector(to_unsigned(1,8) ,
43404	 => std_logic_vector(to_unsigned(1,8) ,
43405	 => std_logic_vector(to_unsigned(0,8) ,
43406	 => std_logic_vector(to_unsigned(1,8) ,
43407	 => std_logic_vector(to_unsigned(12,8) ,
43408	 => std_logic_vector(to_unsigned(29,8) ,
43409	 => std_logic_vector(to_unsigned(37,8) ,
43410	 => std_logic_vector(to_unsigned(6,8) ,
43411	 => std_logic_vector(to_unsigned(2,8) ,
43412	 => std_logic_vector(to_unsigned(1,8) ,
43413	 => std_logic_vector(to_unsigned(0,8) ,
43414	 => std_logic_vector(to_unsigned(0,8) ,
43415	 => std_logic_vector(to_unsigned(1,8) ,
43416	 => std_logic_vector(to_unsigned(1,8) ,
43417	 => std_logic_vector(to_unsigned(1,8) ,
43418	 => std_logic_vector(to_unsigned(5,8) ,
43419	 => std_logic_vector(to_unsigned(1,8) ,
43420	 => std_logic_vector(to_unsigned(0,8) ,
43421	 => std_logic_vector(to_unsigned(0,8) ,
43422	 => std_logic_vector(to_unsigned(0,8) ,
43423	 => std_logic_vector(to_unsigned(2,8) ,
43424	 => std_logic_vector(to_unsigned(2,8) ,
43425	 => std_logic_vector(to_unsigned(2,8) ,
43426	 => std_logic_vector(to_unsigned(3,8) ,
43427	 => std_logic_vector(to_unsigned(3,8) ,
43428	 => std_logic_vector(to_unsigned(3,8) ,
43429	 => std_logic_vector(to_unsigned(2,8) ,
43430	 => std_logic_vector(to_unsigned(2,8) ,
43431	 => std_logic_vector(to_unsigned(1,8) ,
43432	 => std_logic_vector(to_unsigned(3,8) ,
43433	 => std_logic_vector(to_unsigned(8,8) ,
43434	 => std_logic_vector(to_unsigned(1,8) ,
43435	 => std_logic_vector(to_unsigned(0,8) ,
43436	 => std_logic_vector(to_unsigned(0,8) ,
43437	 => std_logic_vector(to_unsigned(0,8) ,
43438	 => std_logic_vector(to_unsigned(3,8) ,
43439	 => std_logic_vector(to_unsigned(5,8) ,
43440	 => std_logic_vector(to_unsigned(6,8) ,
43441	 => std_logic_vector(to_unsigned(4,8) ,
43442	 => std_logic_vector(to_unsigned(3,8) ,
43443	 => std_logic_vector(to_unsigned(3,8) ,
43444	 => std_logic_vector(to_unsigned(2,8) ,
43445	 => std_logic_vector(to_unsigned(1,8) ,
43446	 => std_logic_vector(to_unsigned(1,8) ,
43447	 => std_logic_vector(to_unsigned(2,8) ,
43448	 => std_logic_vector(to_unsigned(10,8) ,
43449	 => std_logic_vector(to_unsigned(10,8) ,
43450	 => std_logic_vector(to_unsigned(4,8) ,
43451	 => std_logic_vector(to_unsigned(1,8) ,
43452	 => std_logic_vector(to_unsigned(1,8) ,
43453	 => std_logic_vector(to_unsigned(1,8) ,
43454	 => std_logic_vector(to_unsigned(1,8) ,
43455	 => std_logic_vector(to_unsigned(1,8) ,
43456	 => std_logic_vector(to_unsigned(1,8) ,
43457	 => std_logic_vector(to_unsigned(2,8) ,
43458	 => std_logic_vector(to_unsigned(4,8) ,
43459	 => std_logic_vector(to_unsigned(4,8) ,
43460	 => std_logic_vector(to_unsigned(3,8) ,
43461	 => std_logic_vector(to_unsigned(2,8) ,
43462	 => std_logic_vector(to_unsigned(1,8) ,
43463	 => std_logic_vector(to_unsigned(0,8) ,
43464	 => std_logic_vector(to_unsigned(1,8) ,
43465	 => std_logic_vector(to_unsigned(24,8) ,
43466	 => std_logic_vector(to_unsigned(51,8) ,
43467	 => std_logic_vector(to_unsigned(47,8) ,
43468	 => std_logic_vector(to_unsigned(41,8) ,
43469	 => std_logic_vector(to_unsigned(34,8) ,
43470	 => std_logic_vector(to_unsigned(17,8) ,
43471	 => std_logic_vector(to_unsigned(10,8) ,
43472	 => std_logic_vector(to_unsigned(7,8) ,
43473	 => std_logic_vector(to_unsigned(6,8) ,
43474	 => std_logic_vector(to_unsigned(11,8) ,
43475	 => std_logic_vector(to_unsigned(19,8) ,
43476	 => std_logic_vector(to_unsigned(2,8) ,
43477	 => std_logic_vector(to_unsigned(0,8) ,
43478	 => std_logic_vector(to_unsigned(1,8) ,
43479	 => std_logic_vector(to_unsigned(1,8) ,
43480	 => std_logic_vector(to_unsigned(1,8) ,
43481	 => std_logic_vector(to_unsigned(1,8) ,
43482	 => std_logic_vector(to_unsigned(1,8) ,
43483	 => std_logic_vector(to_unsigned(1,8) ,
43484	 => std_logic_vector(to_unsigned(2,8) ,
43485	 => std_logic_vector(to_unsigned(6,8) ,
43486	 => std_logic_vector(to_unsigned(5,8) ,
43487	 => std_logic_vector(to_unsigned(5,8) ,
43488	 => std_logic_vector(to_unsigned(3,8) ,
43489	 => std_logic_vector(to_unsigned(3,8) ,
43490	 => std_logic_vector(to_unsigned(3,8) ,
43491	 => std_logic_vector(to_unsigned(2,8) ,
43492	 => std_logic_vector(to_unsigned(1,8) ,
43493	 => std_logic_vector(to_unsigned(1,8) ,
43494	 => std_logic_vector(to_unsigned(1,8) ,
43495	 => std_logic_vector(to_unsigned(1,8) ,
43496	 => std_logic_vector(to_unsigned(1,8) ,
43497	 => std_logic_vector(to_unsigned(1,8) ,
43498	 => std_logic_vector(to_unsigned(1,8) ,
43499	 => std_logic_vector(to_unsigned(1,8) ,
43500	 => std_logic_vector(to_unsigned(1,8) ,
43501	 => std_logic_vector(to_unsigned(1,8) ,
43502	 => std_logic_vector(to_unsigned(1,8) ,
43503	 => std_logic_vector(to_unsigned(1,8) ,
43504	 => std_logic_vector(to_unsigned(2,8) ,
43505	 => std_logic_vector(to_unsigned(1,8) ,
43506	 => std_logic_vector(to_unsigned(1,8) ,
43507	 => std_logic_vector(to_unsigned(1,8) ,
43508	 => std_logic_vector(to_unsigned(2,8) ,
43509	 => std_logic_vector(to_unsigned(2,8) ,
43510	 => std_logic_vector(to_unsigned(3,8) ,
43511	 => std_logic_vector(to_unsigned(4,8) ,
43512	 => std_logic_vector(to_unsigned(2,8) ,
43513	 => std_logic_vector(to_unsigned(2,8) ,
43514	 => std_logic_vector(to_unsigned(2,8) ,
43515	 => std_logic_vector(to_unsigned(3,8) ,
43516	 => std_logic_vector(to_unsigned(3,8) ,
43517	 => std_logic_vector(to_unsigned(3,8) ,
43518	 => std_logic_vector(to_unsigned(3,8) ,
43519	 => std_logic_vector(to_unsigned(2,8) ,
43520	 => std_logic_vector(to_unsigned(3,8) ,
43521	 => std_logic_vector(to_unsigned(87,8) ,
43522	 => std_logic_vector(to_unsigned(84,8) ,
43523	 => std_logic_vector(to_unsigned(84,8) ,
43524	 => std_logic_vector(to_unsigned(78,8) ,
43525	 => std_logic_vector(to_unsigned(79,8) ,
43526	 => std_logic_vector(to_unsigned(84,8) ,
43527	 => std_logic_vector(to_unsigned(86,8) ,
43528	 => std_logic_vector(to_unsigned(53,8) ,
43529	 => std_logic_vector(to_unsigned(45,8) ,
43530	 => std_logic_vector(to_unsigned(49,8) ,
43531	 => std_logic_vector(to_unsigned(48,8) ,
43532	 => std_logic_vector(to_unsigned(49,8) ,
43533	 => std_logic_vector(to_unsigned(48,8) ,
43534	 => std_logic_vector(to_unsigned(93,8) ,
43535	 => std_logic_vector(to_unsigned(122,8) ,
43536	 => std_logic_vector(to_unsigned(118,8) ,
43537	 => std_logic_vector(to_unsigned(101,8) ,
43538	 => std_logic_vector(to_unsigned(116,8) ,
43539	 => std_logic_vector(to_unsigned(138,8) ,
43540	 => std_logic_vector(to_unsigned(131,8) ,
43541	 => std_logic_vector(to_unsigned(141,8) ,
43542	 => std_logic_vector(to_unsigned(133,8) ,
43543	 => std_logic_vector(to_unsigned(128,8) ,
43544	 => std_logic_vector(to_unsigned(138,8) ,
43545	 => std_logic_vector(to_unsigned(141,8) ,
43546	 => std_logic_vector(to_unsigned(136,8) ,
43547	 => std_logic_vector(to_unsigned(141,8) ,
43548	 => std_logic_vector(to_unsigned(138,8) ,
43549	 => std_logic_vector(to_unsigned(125,8) ,
43550	 => std_logic_vector(to_unsigned(138,8) ,
43551	 => std_logic_vector(to_unsigned(131,8) ,
43552	 => std_logic_vector(to_unsigned(133,8) ,
43553	 => std_logic_vector(to_unsigned(134,8) ,
43554	 => std_logic_vector(to_unsigned(141,8) ,
43555	 => std_logic_vector(to_unsigned(144,8) ,
43556	 => std_logic_vector(to_unsigned(154,8) ,
43557	 => std_logic_vector(to_unsigned(156,8) ,
43558	 => std_logic_vector(to_unsigned(156,8) ,
43559	 => std_logic_vector(to_unsigned(157,8) ,
43560	 => std_logic_vector(to_unsigned(146,8) ,
43561	 => std_logic_vector(to_unsigned(96,8) ,
43562	 => std_logic_vector(to_unsigned(109,8) ,
43563	 => std_logic_vector(to_unsigned(91,8) ,
43564	 => std_logic_vector(to_unsigned(105,8) ,
43565	 => std_logic_vector(to_unsigned(119,8) ,
43566	 => std_logic_vector(to_unsigned(103,8) ,
43567	 => std_logic_vector(to_unsigned(111,8) ,
43568	 => std_logic_vector(to_unsigned(130,8) ,
43569	 => std_logic_vector(to_unsigned(142,8) ,
43570	 => std_logic_vector(to_unsigned(144,8) ,
43571	 => std_logic_vector(to_unsigned(138,8) ,
43572	 => std_logic_vector(to_unsigned(142,8) ,
43573	 => std_logic_vector(to_unsigned(136,8) ,
43574	 => std_logic_vector(to_unsigned(114,8) ,
43575	 => std_logic_vector(to_unsigned(103,8) ,
43576	 => std_logic_vector(to_unsigned(96,8) ,
43577	 => std_logic_vector(to_unsigned(100,8) ,
43578	 => std_logic_vector(to_unsigned(105,8) ,
43579	 => std_logic_vector(to_unsigned(100,8) ,
43580	 => std_logic_vector(to_unsigned(92,8) ,
43581	 => std_logic_vector(to_unsigned(97,8) ,
43582	 => std_logic_vector(to_unsigned(99,8) ,
43583	 => std_logic_vector(to_unsigned(85,8) ,
43584	 => std_logic_vector(to_unsigned(100,8) ,
43585	 => std_logic_vector(to_unsigned(105,8) ,
43586	 => std_logic_vector(to_unsigned(99,8) ,
43587	 => std_logic_vector(to_unsigned(88,8) ,
43588	 => std_logic_vector(to_unsigned(85,8) ,
43589	 => std_logic_vector(to_unsigned(90,8) ,
43590	 => std_logic_vector(to_unsigned(90,8) ,
43591	 => std_logic_vector(to_unsigned(90,8) ,
43592	 => std_logic_vector(to_unsigned(69,8) ,
43593	 => std_logic_vector(to_unsigned(8,8) ,
43594	 => std_logic_vector(to_unsigned(6,8) ,
43595	 => std_logic_vector(to_unsigned(8,8) ,
43596	 => std_logic_vector(to_unsigned(3,8) ,
43597	 => std_logic_vector(to_unsigned(4,8) ,
43598	 => std_logic_vector(to_unsigned(14,8) ,
43599	 => std_logic_vector(to_unsigned(60,8) ,
43600	 => std_logic_vector(to_unsigned(107,8) ,
43601	 => std_logic_vector(to_unsigned(100,8) ,
43602	 => std_logic_vector(to_unsigned(93,8) ,
43603	 => std_logic_vector(to_unsigned(103,8) ,
43604	 => std_logic_vector(to_unsigned(108,8) ,
43605	 => std_logic_vector(to_unsigned(118,8) ,
43606	 => std_logic_vector(to_unsigned(100,8) ,
43607	 => std_logic_vector(to_unsigned(81,8) ,
43608	 => std_logic_vector(to_unsigned(76,8) ,
43609	 => std_logic_vector(to_unsigned(76,8) ,
43610	 => std_logic_vector(to_unsigned(81,8) ,
43611	 => std_logic_vector(to_unsigned(23,8) ,
43612	 => std_logic_vector(to_unsigned(8,8) ,
43613	 => std_logic_vector(to_unsigned(21,8) ,
43614	 => std_logic_vector(to_unsigned(12,8) ,
43615	 => std_logic_vector(to_unsigned(23,8) ,
43616	 => std_logic_vector(to_unsigned(57,8) ,
43617	 => std_logic_vector(to_unsigned(14,8) ,
43618	 => std_logic_vector(to_unsigned(6,8) ,
43619	 => std_logic_vector(to_unsigned(9,8) ,
43620	 => std_logic_vector(to_unsigned(6,8) ,
43621	 => std_logic_vector(to_unsigned(4,8) ,
43622	 => std_logic_vector(to_unsigned(5,8) ,
43623	 => std_logic_vector(to_unsigned(6,8) ,
43624	 => std_logic_vector(to_unsigned(1,8) ,
43625	 => std_logic_vector(to_unsigned(10,8) ,
43626	 => std_logic_vector(to_unsigned(115,8) ,
43627	 => std_logic_vector(to_unsigned(100,8) ,
43628	 => std_logic_vector(to_unsigned(93,8) ,
43629	 => std_logic_vector(to_unsigned(109,8) ,
43630	 => std_logic_vector(to_unsigned(104,8) ,
43631	 => std_logic_vector(to_unsigned(105,8) ,
43632	 => std_logic_vector(to_unsigned(101,8) ,
43633	 => std_logic_vector(to_unsigned(100,8) ,
43634	 => std_logic_vector(to_unsigned(88,8) ,
43635	 => std_logic_vector(to_unsigned(96,8) ,
43636	 => std_logic_vector(to_unsigned(99,8) ,
43637	 => std_logic_vector(to_unsigned(97,8) ,
43638	 => std_logic_vector(to_unsigned(104,8) ,
43639	 => std_logic_vector(to_unsigned(99,8) ,
43640	 => std_logic_vector(to_unsigned(107,8) ,
43641	 => std_logic_vector(to_unsigned(104,8) ,
43642	 => std_logic_vector(to_unsigned(95,8) ,
43643	 => std_logic_vector(to_unsigned(114,8) ,
43644	 => std_logic_vector(to_unsigned(37,8) ,
43645	 => std_logic_vector(to_unsigned(4,8) ,
43646	 => std_logic_vector(to_unsigned(3,8) ,
43647	 => std_logic_vector(to_unsigned(2,8) ,
43648	 => std_logic_vector(to_unsigned(1,8) ,
43649	 => std_logic_vector(to_unsigned(26,8) ,
43650	 => std_logic_vector(to_unsigned(133,8) ,
43651	 => std_logic_vector(to_unsigned(138,8) ,
43652	 => std_logic_vector(to_unsigned(131,8) ,
43653	 => std_logic_vector(to_unsigned(121,8) ,
43654	 => std_logic_vector(to_unsigned(105,8) ,
43655	 => std_logic_vector(to_unsigned(95,8) ,
43656	 => std_logic_vector(to_unsigned(99,8) ,
43657	 => std_logic_vector(to_unsigned(90,8) ,
43658	 => std_logic_vector(to_unsigned(88,8) ,
43659	 => std_logic_vector(to_unsigned(81,8) ,
43660	 => std_logic_vector(to_unsigned(85,8) ,
43661	 => std_logic_vector(to_unsigned(87,8) ,
43662	 => std_logic_vector(to_unsigned(87,8) ,
43663	 => std_logic_vector(to_unsigned(88,8) ,
43664	 => std_logic_vector(to_unsigned(103,8) ,
43665	 => std_logic_vector(to_unsigned(107,8) ,
43666	 => std_logic_vector(to_unsigned(97,8) ,
43667	 => std_logic_vector(to_unsigned(111,8) ,
43668	 => std_logic_vector(to_unsigned(122,8) ,
43669	 => std_logic_vector(to_unsigned(144,8) ,
43670	 => std_logic_vector(to_unsigned(45,8) ,
43671	 => std_logic_vector(to_unsigned(1,8) ,
43672	 => std_logic_vector(to_unsigned(4,8) ,
43673	 => std_logic_vector(to_unsigned(2,8) ,
43674	 => std_logic_vector(to_unsigned(1,8) ,
43675	 => std_logic_vector(to_unsigned(8,8) ,
43676	 => std_logic_vector(to_unsigned(61,8) ,
43677	 => std_logic_vector(to_unsigned(133,8) ,
43678	 => std_logic_vector(to_unsigned(35,8) ,
43679	 => std_logic_vector(to_unsigned(3,8) ,
43680	 => std_logic_vector(to_unsigned(8,8) ,
43681	 => std_logic_vector(to_unsigned(8,8) ,
43682	 => std_logic_vector(to_unsigned(8,8) ,
43683	 => std_logic_vector(to_unsigned(2,8) ,
43684	 => std_logic_vector(to_unsigned(4,8) ,
43685	 => std_logic_vector(to_unsigned(82,8) ,
43686	 => std_logic_vector(to_unsigned(100,8) ,
43687	 => std_logic_vector(to_unsigned(105,8) ,
43688	 => std_logic_vector(to_unsigned(114,8) ,
43689	 => std_logic_vector(to_unsigned(104,8) ,
43690	 => std_logic_vector(to_unsigned(114,8) ,
43691	 => std_logic_vector(to_unsigned(108,8) ,
43692	 => std_logic_vector(to_unsigned(97,8) ,
43693	 => std_logic_vector(to_unsigned(95,8) ,
43694	 => std_logic_vector(to_unsigned(91,8) ,
43695	 => std_logic_vector(to_unsigned(64,8) ,
43696	 => std_logic_vector(to_unsigned(47,8) ,
43697	 => std_logic_vector(to_unsigned(5,8) ,
43698	 => std_logic_vector(to_unsigned(6,8) ,
43699	 => std_logic_vector(to_unsigned(13,8) ,
43700	 => std_logic_vector(to_unsigned(5,8) ,
43701	 => std_logic_vector(to_unsigned(4,8) ,
43702	 => std_logic_vector(to_unsigned(1,8) ,
43703	 => std_logic_vector(to_unsigned(25,8) ,
43704	 => std_logic_vector(to_unsigned(105,8) ,
43705	 => std_logic_vector(to_unsigned(28,8) ,
43706	 => std_logic_vector(to_unsigned(6,8) ,
43707	 => std_logic_vector(to_unsigned(11,8) ,
43708	 => std_logic_vector(to_unsigned(30,8) ,
43709	 => std_logic_vector(to_unsigned(28,8) ,
43710	 => std_logic_vector(to_unsigned(17,8) ,
43711	 => std_logic_vector(to_unsigned(93,8) ,
43712	 => std_logic_vector(to_unsigned(118,8) ,
43713	 => std_logic_vector(to_unsigned(91,8) ,
43714	 => std_logic_vector(to_unsigned(93,8) ,
43715	 => std_logic_vector(to_unsigned(82,8) ,
43716	 => std_logic_vector(to_unsigned(67,8) ,
43717	 => std_logic_vector(to_unsigned(61,8) ,
43718	 => std_logic_vector(to_unsigned(54,8) ,
43719	 => std_logic_vector(to_unsigned(43,8) ,
43720	 => std_logic_vector(to_unsigned(36,8) ,
43721	 => std_logic_vector(to_unsigned(25,8) ,
43722	 => std_logic_vector(to_unsigned(16,8) ,
43723	 => std_logic_vector(to_unsigned(10,8) ,
43724	 => std_logic_vector(to_unsigned(6,8) ,
43725	 => std_logic_vector(to_unsigned(2,8) ,
43726	 => std_logic_vector(to_unsigned(2,8) ,
43727	 => std_logic_vector(to_unsigned(10,8) ,
43728	 => std_logic_vector(to_unsigned(37,8) ,
43729	 => std_logic_vector(to_unsigned(41,8) ,
43730	 => std_logic_vector(to_unsigned(7,8) ,
43731	 => std_logic_vector(to_unsigned(3,8) ,
43732	 => std_logic_vector(to_unsigned(1,8) ,
43733	 => std_logic_vector(to_unsigned(0,8) ,
43734	 => std_logic_vector(to_unsigned(0,8) ,
43735	 => std_logic_vector(to_unsigned(1,8) ,
43736	 => std_logic_vector(to_unsigned(0,8) ,
43737	 => std_logic_vector(to_unsigned(6,8) ,
43738	 => std_logic_vector(to_unsigned(13,8) ,
43739	 => std_logic_vector(to_unsigned(1,8) ,
43740	 => std_logic_vector(to_unsigned(0,8) ,
43741	 => std_logic_vector(to_unsigned(0,8) ,
43742	 => std_logic_vector(to_unsigned(1,8) ,
43743	 => std_logic_vector(to_unsigned(2,8) ,
43744	 => std_logic_vector(to_unsigned(3,8) ,
43745	 => std_logic_vector(to_unsigned(4,8) ,
43746	 => std_logic_vector(to_unsigned(5,8) ,
43747	 => std_logic_vector(to_unsigned(3,8) ,
43748	 => std_logic_vector(to_unsigned(3,8) ,
43749	 => std_logic_vector(to_unsigned(4,8) ,
43750	 => std_logic_vector(to_unsigned(5,8) ,
43751	 => std_logic_vector(to_unsigned(2,8) ,
43752	 => std_logic_vector(to_unsigned(2,8) ,
43753	 => std_logic_vector(to_unsigned(9,8) ,
43754	 => std_logic_vector(to_unsigned(4,8) ,
43755	 => std_logic_vector(to_unsigned(0,8) ,
43756	 => std_logic_vector(to_unsigned(1,8) ,
43757	 => std_logic_vector(to_unsigned(0,8) ,
43758	 => std_logic_vector(to_unsigned(1,8) ,
43759	 => std_logic_vector(to_unsigned(2,8) ,
43760	 => std_logic_vector(to_unsigned(3,8) ,
43761	 => std_logic_vector(to_unsigned(4,8) ,
43762	 => std_logic_vector(to_unsigned(6,8) ,
43763	 => std_logic_vector(to_unsigned(3,8) ,
43764	 => std_logic_vector(to_unsigned(1,8) ,
43765	 => std_logic_vector(to_unsigned(1,8) ,
43766	 => std_logic_vector(to_unsigned(1,8) ,
43767	 => std_logic_vector(to_unsigned(2,8) ,
43768	 => std_logic_vector(to_unsigned(9,8) ,
43769	 => std_logic_vector(to_unsigned(10,8) ,
43770	 => std_logic_vector(to_unsigned(3,8) ,
43771	 => std_logic_vector(to_unsigned(1,8) ,
43772	 => std_logic_vector(to_unsigned(1,8) ,
43773	 => std_logic_vector(to_unsigned(1,8) ,
43774	 => std_logic_vector(to_unsigned(1,8) ,
43775	 => std_logic_vector(to_unsigned(1,8) ,
43776	 => std_logic_vector(to_unsigned(1,8) ,
43777	 => std_logic_vector(to_unsigned(2,8) ,
43778	 => std_logic_vector(to_unsigned(2,8) ,
43779	 => std_logic_vector(to_unsigned(3,8) ,
43780	 => std_logic_vector(to_unsigned(2,8) ,
43781	 => std_logic_vector(to_unsigned(2,8) ,
43782	 => std_logic_vector(to_unsigned(0,8) ,
43783	 => std_logic_vector(to_unsigned(0,8) ,
43784	 => std_logic_vector(to_unsigned(8,8) ,
43785	 => std_logic_vector(to_unsigned(27,8) ,
43786	 => std_logic_vector(to_unsigned(38,8) ,
43787	 => std_logic_vector(to_unsigned(55,8) ,
43788	 => std_logic_vector(to_unsigned(39,8) ,
43789	 => std_logic_vector(to_unsigned(34,8) ,
43790	 => std_logic_vector(to_unsigned(22,8) ,
43791	 => std_logic_vector(to_unsigned(10,8) ,
43792	 => std_logic_vector(to_unsigned(6,8) ,
43793	 => std_logic_vector(to_unsigned(5,8) ,
43794	 => std_logic_vector(to_unsigned(11,8) ,
43795	 => std_logic_vector(to_unsigned(21,8) ,
43796	 => std_logic_vector(to_unsigned(5,8) ,
43797	 => std_logic_vector(to_unsigned(0,8) ,
43798	 => std_logic_vector(to_unsigned(1,8) ,
43799	 => std_logic_vector(to_unsigned(1,8) ,
43800	 => std_logic_vector(to_unsigned(1,8) ,
43801	 => std_logic_vector(to_unsigned(1,8) ,
43802	 => std_logic_vector(to_unsigned(0,8) ,
43803	 => std_logic_vector(to_unsigned(1,8) ,
43804	 => std_logic_vector(to_unsigned(3,8) ,
43805	 => std_logic_vector(to_unsigned(4,8) ,
43806	 => std_logic_vector(to_unsigned(5,8) ,
43807	 => std_logic_vector(to_unsigned(3,8) ,
43808	 => std_logic_vector(to_unsigned(3,8) ,
43809	 => std_logic_vector(to_unsigned(2,8) ,
43810	 => std_logic_vector(to_unsigned(2,8) ,
43811	 => std_logic_vector(to_unsigned(1,8) ,
43812	 => std_logic_vector(to_unsigned(0,8) ,
43813	 => std_logic_vector(to_unsigned(1,8) ,
43814	 => std_logic_vector(to_unsigned(1,8) ,
43815	 => std_logic_vector(to_unsigned(1,8) ,
43816	 => std_logic_vector(to_unsigned(1,8) ,
43817	 => std_logic_vector(to_unsigned(1,8) ,
43818	 => std_logic_vector(to_unsigned(1,8) ,
43819	 => std_logic_vector(to_unsigned(1,8) ,
43820	 => std_logic_vector(to_unsigned(1,8) ,
43821	 => std_logic_vector(to_unsigned(1,8) ,
43822	 => std_logic_vector(to_unsigned(1,8) ,
43823	 => std_logic_vector(to_unsigned(1,8) ,
43824	 => std_logic_vector(to_unsigned(1,8) ,
43825	 => std_logic_vector(to_unsigned(1,8) ,
43826	 => std_logic_vector(to_unsigned(1,8) ,
43827	 => std_logic_vector(to_unsigned(2,8) ,
43828	 => std_logic_vector(to_unsigned(2,8) ,
43829	 => std_logic_vector(to_unsigned(1,8) ,
43830	 => std_logic_vector(to_unsigned(2,8) ,
43831	 => std_logic_vector(to_unsigned(2,8) ,
43832	 => std_logic_vector(to_unsigned(3,8) ,
43833	 => std_logic_vector(to_unsigned(2,8) ,
43834	 => std_logic_vector(to_unsigned(2,8) ,
43835	 => std_logic_vector(to_unsigned(3,8) ,
43836	 => std_logic_vector(to_unsigned(2,8) ,
43837	 => std_logic_vector(to_unsigned(2,8) ,
43838	 => std_logic_vector(to_unsigned(2,8) ,
43839	 => std_logic_vector(to_unsigned(2,8) ,
43840	 => std_logic_vector(to_unsigned(2,8) ,
43841	 => std_logic_vector(to_unsigned(77,8) ,
43842	 => std_logic_vector(to_unsigned(71,8) ,
43843	 => std_logic_vector(to_unsigned(71,8) ,
43844	 => std_logic_vector(to_unsigned(86,8) ,
43845	 => std_logic_vector(to_unsigned(87,8) ,
43846	 => std_logic_vector(to_unsigned(80,8) ,
43847	 => std_logic_vector(to_unsigned(84,8) ,
43848	 => std_logic_vector(to_unsigned(57,8) ,
43849	 => std_logic_vector(to_unsigned(41,8) ,
43850	 => std_logic_vector(to_unsigned(45,8) ,
43851	 => std_logic_vector(to_unsigned(47,8) ,
43852	 => std_logic_vector(to_unsigned(49,8) ,
43853	 => std_logic_vector(to_unsigned(45,8) ,
43854	 => std_logic_vector(to_unsigned(82,8) ,
43855	 => std_logic_vector(to_unsigned(115,8) ,
43856	 => std_logic_vector(to_unsigned(108,8) ,
43857	 => std_logic_vector(to_unsigned(111,8) ,
43858	 => std_logic_vector(to_unsigned(114,8) ,
43859	 => std_logic_vector(to_unsigned(112,8) ,
43860	 => std_logic_vector(to_unsigned(128,8) ,
43861	 => std_logic_vector(to_unsigned(128,8) ,
43862	 => std_logic_vector(to_unsigned(124,8) ,
43863	 => std_logic_vector(to_unsigned(128,8) ,
43864	 => std_logic_vector(to_unsigned(138,8) ,
43865	 => std_logic_vector(to_unsigned(136,8) ,
43866	 => std_logic_vector(to_unsigned(151,8) ,
43867	 => std_logic_vector(to_unsigned(149,8) ,
43868	 => std_logic_vector(to_unsigned(144,8) ,
43869	 => std_logic_vector(to_unsigned(149,8) ,
43870	 => std_logic_vector(to_unsigned(151,8) ,
43871	 => std_logic_vector(to_unsigned(144,8) ,
43872	 => std_logic_vector(to_unsigned(146,8) ,
43873	 => std_logic_vector(to_unsigned(151,8) ,
43874	 => std_logic_vector(to_unsigned(146,8) ,
43875	 => std_logic_vector(to_unsigned(154,8) ,
43876	 => std_logic_vector(to_unsigned(154,8) ,
43877	 => std_logic_vector(to_unsigned(156,8) ,
43878	 => std_logic_vector(to_unsigned(156,8) ,
43879	 => std_logic_vector(to_unsigned(157,8) ,
43880	 => std_logic_vector(to_unsigned(149,8) ,
43881	 => std_logic_vector(to_unsigned(100,8) ,
43882	 => std_logic_vector(to_unsigned(109,8) ,
43883	 => std_logic_vector(to_unsigned(96,8) ,
43884	 => std_logic_vector(to_unsigned(91,8) ,
43885	 => std_logic_vector(to_unsigned(103,8) ,
43886	 => std_logic_vector(to_unsigned(99,8) ,
43887	 => std_logic_vector(to_unsigned(111,8) ,
43888	 => std_logic_vector(to_unsigned(136,8) ,
43889	 => std_logic_vector(to_unsigned(147,8) ,
43890	 => std_logic_vector(to_unsigned(130,8) ,
43891	 => std_logic_vector(to_unsigned(128,8) ,
43892	 => std_logic_vector(to_unsigned(131,8) ,
43893	 => std_logic_vector(to_unsigned(125,8) ,
43894	 => std_logic_vector(to_unsigned(108,8) ,
43895	 => std_logic_vector(to_unsigned(92,8) ,
43896	 => std_logic_vector(to_unsigned(99,8) ,
43897	 => std_logic_vector(to_unsigned(103,8) ,
43898	 => std_logic_vector(to_unsigned(103,8) ,
43899	 => std_logic_vector(to_unsigned(99,8) ,
43900	 => std_logic_vector(to_unsigned(92,8) ,
43901	 => std_logic_vector(to_unsigned(100,8) ,
43902	 => std_logic_vector(to_unsigned(92,8) ,
43903	 => std_logic_vector(to_unsigned(78,8) ,
43904	 => std_logic_vector(to_unsigned(93,8) ,
43905	 => std_logic_vector(to_unsigned(97,8) ,
43906	 => std_logic_vector(to_unsigned(81,8) ,
43907	 => std_logic_vector(to_unsigned(80,8) ,
43908	 => std_logic_vector(to_unsigned(79,8) ,
43909	 => std_logic_vector(to_unsigned(82,8) ,
43910	 => std_logic_vector(to_unsigned(81,8) ,
43911	 => std_logic_vector(to_unsigned(85,8) ,
43912	 => std_logic_vector(to_unsigned(69,8) ,
43913	 => std_logic_vector(to_unsigned(16,8) ,
43914	 => std_logic_vector(to_unsigned(11,8) ,
43915	 => std_logic_vector(to_unsigned(19,8) ,
43916	 => std_logic_vector(to_unsigned(26,8) ,
43917	 => std_logic_vector(to_unsigned(69,8) ,
43918	 => std_logic_vector(to_unsigned(109,8) ,
43919	 => std_logic_vector(to_unsigned(125,8) ,
43920	 => std_logic_vector(to_unsigned(112,8) ,
43921	 => std_logic_vector(to_unsigned(107,8) ,
43922	 => std_logic_vector(to_unsigned(103,8) ,
43923	 => std_logic_vector(to_unsigned(103,8) ,
43924	 => std_logic_vector(to_unsigned(99,8) ,
43925	 => std_logic_vector(to_unsigned(114,8) ,
43926	 => std_logic_vector(to_unsigned(96,8) ,
43927	 => std_logic_vector(to_unsigned(82,8) ,
43928	 => std_logic_vector(to_unsigned(87,8) ,
43929	 => std_logic_vector(to_unsigned(69,8) ,
43930	 => std_logic_vector(to_unsigned(15,8) ,
43931	 => std_logic_vector(to_unsigned(7,8) ,
43932	 => std_logic_vector(to_unsigned(10,8) ,
43933	 => std_logic_vector(to_unsigned(12,8) ,
43934	 => std_logic_vector(to_unsigned(12,8) ,
43935	 => std_logic_vector(to_unsigned(15,8) ,
43936	 => std_logic_vector(to_unsigned(10,8) ,
43937	 => std_logic_vector(to_unsigned(6,8) ,
43938	 => std_logic_vector(to_unsigned(8,8) ,
43939	 => std_logic_vector(to_unsigned(6,8) ,
43940	 => std_logic_vector(to_unsigned(8,8) ,
43941	 => std_logic_vector(to_unsigned(5,8) ,
43942	 => std_logic_vector(to_unsigned(2,8) ,
43943	 => std_logic_vector(to_unsigned(1,8) ,
43944	 => std_logic_vector(to_unsigned(8,8) ,
43945	 => std_logic_vector(to_unsigned(66,8) ,
43946	 => std_logic_vector(to_unsigned(103,8) ,
43947	 => std_logic_vector(to_unsigned(88,8) ,
43948	 => std_logic_vector(to_unsigned(95,8) ,
43949	 => std_logic_vector(to_unsigned(92,8) ,
43950	 => std_logic_vector(to_unsigned(103,8) ,
43951	 => std_logic_vector(to_unsigned(100,8) ,
43952	 => std_logic_vector(to_unsigned(101,8) ,
43953	 => std_logic_vector(to_unsigned(111,8) ,
43954	 => std_logic_vector(to_unsigned(81,8) ,
43955	 => std_logic_vector(to_unsigned(79,8) ,
43956	 => std_logic_vector(to_unsigned(103,8) ,
43957	 => std_logic_vector(to_unsigned(91,8) ,
43958	 => std_logic_vector(to_unsigned(87,8) ,
43959	 => std_logic_vector(to_unsigned(93,8) ,
43960	 => std_logic_vector(to_unsigned(97,8) ,
43961	 => std_logic_vector(to_unsigned(91,8) ,
43962	 => std_logic_vector(to_unsigned(92,8) ,
43963	 => std_logic_vector(to_unsigned(97,8) ,
43964	 => std_logic_vector(to_unsigned(20,8) ,
43965	 => std_logic_vector(to_unsigned(3,8) ,
43966	 => std_logic_vector(to_unsigned(4,8) ,
43967	 => std_logic_vector(to_unsigned(4,8) ,
43968	 => std_logic_vector(to_unsigned(1,8) ,
43969	 => std_logic_vector(to_unsigned(13,8) ,
43970	 => std_logic_vector(to_unsigned(111,8) ,
43971	 => std_logic_vector(to_unsigned(125,8) ,
43972	 => std_logic_vector(to_unsigned(118,8) ,
43973	 => std_logic_vector(to_unsigned(116,8) ,
43974	 => std_logic_vector(to_unsigned(103,8) ,
43975	 => std_logic_vector(to_unsigned(79,8) ,
43976	 => std_logic_vector(to_unsigned(96,8) ,
43977	 => std_logic_vector(to_unsigned(104,8) ,
43978	 => std_logic_vector(to_unsigned(99,8) ,
43979	 => std_logic_vector(to_unsigned(90,8) ,
43980	 => std_logic_vector(to_unsigned(88,8) ,
43981	 => std_logic_vector(to_unsigned(87,8) ,
43982	 => std_logic_vector(to_unsigned(91,8) ,
43983	 => std_logic_vector(to_unsigned(91,8) ,
43984	 => std_logic_vector(to_unsigned(86,8) ,
43985	 => std_logic_vector(to_unsigned(81,8) ,
43986	 => std_logic_vector(to_unsigned(93,8) ,
43987	 => std_logic_vector(to_unsigned(91,8) ,
43988	 => std_logic_vector(to_unsigned(99,8) ,
43989	 => std_logic_vector(to_unsigned(130,8) ,
43990	 => std_logic_vector(to_unsigned(70,8) ,
43991	 => std_logic_vector(to_unsigned(12,8) ,
43992	 => std_logic_vector(to_unsigned(8,8) ,
43993	 => std_logic_vector(to_unsigned(11,8) ,
43994	 => std_logic_vector(to_unsigned(37,8) ,
43995	 => std_logic_vector(to_unsigned(97,8) ,
43996	 => std_logic_vector(to_unsigned(103,8) ,
43997	 => std_logic_vector(to_unsigned(118,8) ,
43998	 => std_logic_vector(to_unsigned(20,8) ,
43999	 => std_logic_vector(to_unsigned(2,8) ,
44000	 => std_logic_vector(to_unsigned(9,8) ,
44001	 => std_logic_vector(to_unsigned(6,8) ,
44002	 => std_logic_vector(to_unsigned(4,8) ,
44003	 => std_logic_vector(to_unsigned(0,8) ,
44004	 => std_logic_vector(to_unsigned(25,8) ,
44005	 => std_logic_vector(to_unsigned(122,8) ,
44006	 => std_logic_vector(to_unsigned(96,8) ,
44007	 => std_logic_vector(to_unsigned(96,8) ,
44008	 => std_logic_vector(to_unsigned(100,8) ,
44009	 => std_logic_vector(to_unsigned(101,8) ,
44010	 => std_logic_vector(to_unsigned(99,8) ,
44011	 => std_logic_vector(to_unsigned(96,8) ,
44012	 => std_logic_vector(to_unsigned(101,8) ,
44013	 => std_logic_vector(to_unsigned(101,8) ,
44014	 => std_logic_vector(to_unsigned(86,8) ,
44015	 => std_logic_vector(to_unsigned(69,8) ,
44016	 => std_logic_vector(to_unsigned(37,8) ,
44017	 => std_logic_vector(to_unsigned(4,8) ,
44018	 => std_logic_vector(to_unsigned(6,8) ,
44019	 => std_logic_vector(to_unsigned(6,8) ,
44020	 => std_logic_vector(to_unsigned(4,8) ,
44021	 => std_logic_vector(to_unsigned(5,8) ,
44022	 => std_logic_vector(to_unsigned(1,8) ,
44023	 => std_logic_vector(to_unsigned(21,8) ,
44024	 => std_logic_vector(to_unsigned(81,8) ,
44025	 => std_logic_vector(to_unsigned(10,8) ,
44026	 => std_logic_vector(to_unsigned(7,8) ,
44027	 => std_logic_vector(to_unsigned(10,8) ,
44028	 => std_logic_vector(to_unsigned(29,8) ,
44029	 => std_logic_vector(to_unsigned(22,8) ,
44030	 => std_logic_vector(to_unsigned(21,8) ,
44031	 => std_logic_vector(to_unsigned(104,8) ,
44032	 => std_logic_vector(to_unsigned(84,8) ,
44033	 => std_logic_vector(to_unsigned(78,8) ,
44034	 => std_logic_vector(to_unsigned(115,8) ,
44035	 => std_logic_vector(to_unsigned(93,8) ,
44036	 => std_logic_vector(to_unsigned(78,8) ,
44037	 => std_logic_vector(to_unsigned(104,8) ,
44038	 => std_logic_vector(to_unsigned(107,8) ,
44039	 => std_logic_vector(to_unsigned(77,8) ,
44040	 => std_logic_vector(to_unsigned(99,8) ,
44041	 => std_logic_vector(to_unsigned(122,8) ,
44042	 => std_logic_vector(to_unsigned(133,8) ,
44043	 => std_logic_vector(to_unsigned(105,8) ,
44044	 => std_logic_vector(to_unsigned(92,8) ,
44045	 => std_logic_vector(to_unsigned(72,8) ,
44046	 => std_logic_vector(to_unsigned(25,8) ,
44047	 => std_logic_vector(to_unsigned(14,8) ,
44048	 => std_logic_vector(to_unsigned(49,8) ,
44049	 => std_logic_vector(to_unsigned(25,8) ,
44050	 => std_logic_vector(to_unsigned(13,8) ,
44051	 => std_logic_vector(to_unsigned(3,8) ,
44052	 => std_logic_vector(to_unsigned(1,8) ,
44053	 => std_logic_vector(to_unsigned(2,8) ,
44054	 => std_logic_vector(to_unsigned(1,8) ,
44055	 => std_logic_vector(to_unsigned(1,8) ,
44056	 => std_logic_vector(to_unsigned(1,8) ,
44057	 => std_logic_vector(to_unsigned(12,8) ,
44058	 => std_logic_vector(to_unsigned(9,8) ,
44059	 => std_logic_vector(to_unsigned(0,8) ,
44060	 => std_logic_vector(to_unsigned(0,8) ,
44061	 => std_logic_vector(to_unsigned(0,8) ,
44062	 => std_logic_vector(to_unsigned(1,8) ,
44063	 => std_logic_vector(to_unsigned(1,8) ,
44064	 => std_logic_vector(to_unsigned(1,8) ,
44065	 => std_logic_vector(to_unsigned(1,8) ,
44066	 => std_logic_vector(to_unsigned(1,8) ,
44067	 => std_logic_vector(to_unsigned(1,8) ,
44068	 => std_logic_vector(to_unsigned(1,8) ,
44069	 => std_logic_vector(to_unsigned(2,8) ,
44070	 => std_logic_vector(to_unsigned(2,8) ,
44071	 => std_logic_vector(to_unsigned(2,8) ,
44072	 => std_logic_vector(to_unsigned(2,8) ,
44073	 => std_logic_vector(to_unsigned(4,8) ,
44074	 => std_logic_vector(to_unsigned(6,8) ,
44075	 => std_logic_vector(to_unsigned(0,8) ,
44076	 => std_logic_vector(to_unsigned(1,8) ,
44077	 => std_logic_vector(to_unsigned(1,8) ,
44078	 => std_logic_vector(to_unsigned(0,8) ,
44079	 => std_logic_vector(to_unsigned(0,8) ,
44080	 => std_logic_vector(to_unsigned(0,8) ,
44081	 => std_logic_vector(to_unsigned(0,8) ,
44082	 => std_logic_vector(to_unsigned(1,8) ,
44083	 => std_logic_vector(to_unsigned(1,8) ,
44084	 => std_logic_vector(to_unsigned(2,8) ,
44085	 => std_logic_vector(to_unsigned(1,8) ,
44086	 => std_logic_vector(to_unsigned(1,8) ,
44087	 => std_logic_vector(to_unsigned(1,8) ,
44088	 => std_logic_vector(to_unsigned(6,8) ,
44089	 => std_logic_vector(to_unsigned(10,8) ,
44090	 => std_logic_vector(to_unsigned(3,8) ,
44091	 => std_logic_vector(to_unsigned(1,8) ,
44092	 => std_logic_vector(to_unsigned(1,8) ,
44093	 => std_logic_vector(to_unsigned(1,8) ,
44094	 => std_logic_vector(to_unsigned(1,8) ,
44095	 => std_logic_vector(to_unsigned(1,8) ,
44096	 => std_logic_vector(to_unsigned(2,8) ,
44097	 => std_logic_vector(to_unsigned(3,8) ,
44098	 => std_logic_vector(to_unsigned(5,8) ,
44099	 => std_logic_vector(to_unsigned(4,8) ,
44100	 => std_logic_vector(to_unsigned(3,8) ,
44101	 => std_logic_vector(to_unsigned(1,8) ,
44102	 => std_logic_vector(to_unsigned(0,8) ,
44103	 => std_logic_vector(to_unsigned(6,8) ,
44104	 => std_logic_vector(to_unsigned(18,8) ,
44105	 => std_logic_vector(to_unsigned(30,8) ,
44106	 => std_logic_vector(to_unsigned(31,8) ,
44107	 => std_logic_vector(to_unsigned(37,8) ,
44108	 => std_logic_vector(to_unsigned(32,8) ,
44109	 => std_logic_vector(to_unsigned(30,8) ,
44110	 => std_logic_vector(to_unsigned(30,8) ,
44111	 => std_logic_vector(to_unsigned(14,8) ,
44112	 => std_logic_vector(to_unsigned(7,8) ,
44113	 => std_logic_vector(to_unsigned(5,8) ,
44114	 => std_logic_vector(to_unsigned(9,8) ,
44115	 => std_logic_vector(to_unsigned(16,8) ,
44116	 => std_logic_vector(to_unsigned(9,8) ,
44117	 => std_logic_vector(to_unsigned(0,8) ,
44118	 => std_logic_vector(to_unsigned(0,8) ,
44119	 => std_logic_vector(to_unsigned(0,8) ,
44120	 => std_logic_vector(to_unsigned(0,8) ,
44121	 => std_logic_vector(to_unsigned(1,8) ,
44122	 => std_logic_vector(to_unsigned(1,8) ,
44123	 => std_logic_vector(to_unsigned(1,8) ,
44124	 => std_logic_vector(to_unsigned(4,8) ,
44125	 => std_logic_vector(to_unsigned(3,8) ,
44126	 => std_logic_vector(to_unsigned(6,8) ,
44127	 => std_logic_vector(to_unsigned(2,8) ,
44128	 => std_logic_vector(to_unsigned(1,8) ,
44129	 => std_logic_vector(to_unsigned(2,8) ,
44130	 => std_logic_vector(to_unsigned(1,8) ,
44131	 => std_logic_vector(to_unsigned(0,8) ,
44132	 => std_logic_vector(to_unsigned(1,8) ,
44133	 => std_logic_vector(to_unsigned(1,8) ,
44134	 => std_logic_vector(to_unsigned(1,8) ,
44135	 => std_logic_vector(to_unsigned(1,8) ,
44136	 => std_logic_vector(to_unsigned(1,8) ,
44137	 => std_logic_vector(to_unsigned(1,8) ,
44138	 => std_logic_vector(to_unsigned(1,8) ,
44139	 => std_logic_vector(to_unsigned(1,8) ,
44140	 => std_logic_vector(to_unsigned(1,8) ,
44141	 => std_logic_vector(to_unsigned(1,8) ,
44142	 => std_logic_vector(to_unsigned(1,8) ,
44143	 => std_logic_vector(to_unsigned(1,8) ,
44144	 => std_logic_vector(to_unsigned(1,8) ,
44145	 => std_logic_vector(to_unsigned(1,8) ,
44146	 => std_logic_vector(to_unsigned(2,8) ,
44147	 => std_logic_vector(to_unsigned(1,8) ,
44148	 => std_logic_vector(to_unsigned(2,8) ,
44149	 => std_logic_vector(to_unsigned(2,8) ,
44150	 => std_logic_vector(to_unsigned(1,8) ,
44151	 => std_logic_vector(to_unsigned(2,8) ,
44152	 => std_logic_vector(to_unsigned(3,8) ,
44153	 => std_logic_vector(to_unsigned(3,8) ,
44154	 => std_logic_vector(to_unsigned(2,8) ,
44155	 => std_logic_vector(to_unsigned(2,8) ,
44156	 => std_logic_vector(to_unsigned(2,8) ,
44157	 => std_logic_vector(to_unsigned(2,8) ,
44158	 => std_logic_vector(to_unsigned(3,8) ,
44159	 => std_logic_vector(to_unsigned(3,8) ,
44160	 => std_logic_vector(to_unsigned(3,8) ,
44161	 => std_logic_vector(to_unsigned(73,8) ,
44162	 => std_logic_vector(to_unsigned(81,8) ,
44163	 => std_logic_vector(to_unsigned(78,8) ,
44164	 => std_logic_vector(to_unsigned(61,8) ,
44165	 => std_logic_vector(to_unsigned(66,8) ,
44166	 => std_logic_vector(to_unsigned(65,8) ,
44167	 => std_logic_vector(to_unsigned(76,8) ,
44168	 => std_logic_vector(to_unsigned(52,8) ,
44169	 => std_logic_vector(to_unsigned(37,8) ,
44170	 => std_logic_vector(to_unsigned(43,8) ,
44171	 => std_logic_vector(to_unsigned(41,8) ,
44172	 => std_logic_vector(to_unsigned(48,8) ,
44173	 => std_logic_vector(to_unsigned(54,8) ,
44174	 => std_logic_vector(to_unsigned(82,8) ,
44175	 => std_logic_vector(to_unsigned(125,8) ,
44176	 => std_logic_vector(to_unsigned(125,8) ,
44177	 => std_logic_vector(to_unsigned(107,8) ,
44178	 => std_logic_vector(to_unsigned(119,8) ,
44179	 => std_logic_vector(to_unsigned(118,8) ,
44180	 => std_logic_vector(to_unsigned(124,8) ,
44181	 => std_logic_vector(to_unsigned(121,8) ,
44182	 => std_logic_vector(to_unsigned(125,8) ,
44183	 => std_logic_vector(to_unsigned(133,8) ,
44184	 => std_logic_vector(to_unsigned(134,8) ,
44185	 => std_logic_vector(to_unsigned(138,8) ,
44186	 => std_logic_vector(to_unsigned(146,8) ,
44187	 => std_logic_vector(to_unsigned(142,8) ,
44188	 => std_logic_vector(to_unsigned(141,8) ,
44189	 => std_logic_vector(to_unsigned(144,8) ,
44190	 => std_logic_vector(to_unsigned(151,8) ,
44191	 => std_logic_vector(to_unsigned(142,8) ,
44192	 => std_logic_vector(to_unsigned(151,8) ,
44193	 => std_logic_vector(to_unsigned(149,8) ,
44194	 => std_logic_vector(to_unsigned(144,8) ,
44195	 => std_logic_vector(to_unsigned(151,8) ,
44196	 => std_logic_vector(to_unsigned(147,8) ,
44197	 => std_logic_vector(to_unsigned(154,8) ,
44198	 => std_logic_vector(to_unsigned(147,8) ,
44199	 => std_logic_vector(to_unsigned(159,8) ,
44200	 => std_logic_vector(to_unsigned(147,8) ,
44201	 => std_logic_vector(to_unsigned(88,8) ,
44202	 => std_logic_vector(to_unsigned(93,8) ,
44203	 => std_logic_vector(to_unsigned(97,8) ,
44204	 => std_logic_vector(to_unsigned(93,8) ,
44205	 => std_logic_vector(to_unsigned(109,8) ,
44206	 => std_logic_vector(to_unsigned(90,8) ,
44207	 => std_logic_vector(to_unsigned(104,8) ,
44208	 => std_logic_vector(to_unsigned(121,8) ,
44209	 => std_logic_vector(to_unsigned(118,8) ,
44210	 => std_logic_vector(to_unsigned(111,8) ,
44211	 => std_logic_vector(to_unsigned(128,8) ,
44212	 => std_logic_vector(to_unsigned(136,8) ,
44213	 => std_logic_vector(to_unsigned(118,8) ,
44214	 => std_logic_vector(to_unsigned(104,8) ,
44215	 => std_logic_vector(to_unsigned(90,8) ,
44216	 => std_logic_vector(to_unsigned(82,8) ,
44217	 => std_logic_vector(to_unsigned(88,8) ,
44218	 => std_logic_vector(to_unsigned(90,8) ,
44219	 => std_logic_vector(to_unsigned(92,8) ,
44220	 => std_logic_vector(to_unsigned(92,8) ,
44221	 => std_logic_vector(to_unsigned(91,8) ,
44222	 => std_logic_vector(to_unsigned(91,8) ,
44223	 => std_logic_vector(to_unsigned(92,8) ,
44224	 => std_logic_vector(to_unsigned(95,8) ,
44225	 => std_logic_vector(to_unsigned(97,8) ,
44226	 => std_logic_vector(to_unsigned(91,8) ,
44227	 => std_logic_vector(to_unsigned(87,8) ,
44228	 => std_logic_vector(to_unsigned(87,8) ,
44229	 => std_logic_vector(to_unsigned(84,8) ,
44230	 => std_logic_vector(to_unsigned(82,8) ,
44231	 => std_logic_vector(to_unsigned(82,8) ,
44232	 => std_logic_vector(to_unsigned(76,8) ,
44233	 => std_logic_vector(to_unsigned(65,8) ,
44234	 => std_logic_vector(to_unsigned(72,8) ,
44235	 => std_logic_vector(to_unsigned(93,8) ,
44236	 => std_logic_vector(to_unsigned(90,8) ,
44237	 => std_logic_vector(to_unsigned(112,8) ,
44238	 => std_logic_vector(to_unsigned(107,8) ,
44239	 => std_logic_vector(to_unsigned(111,8) ,
44240	 => std_logic_vector(to_unsigned(108,8) ,
44241	 => std_logic_vector(to_unsigned(95,8) ,
44242	 => std_logic_vector(to_unsigned(84,8) ,
44243	 => std_logic_vector(to_unsigned(86,8) ,
44244	 => std_logic_vector(to_unsigned(92,8) ,
44245	 => std_logic_vector(to_unsigned(108,8) ,
44246	 => std_logic_vector(to_unsigned(100,8) ,
44247	 => std_logic_vector(to_unsigned(91,8) ,
44248	 => std_logic_vector(to_unsigned(87,8) ,
44249	 => std_logic_vector(to_unsigned(25,8) ,
44250	 => std_logic_vector(to_unsigned(2,8) ,
44251	 => std_logic_vector(to_unsigned(5,8) ,
44252	 => std_logic_vector(to_unsigned(11,8) ,
44253	 => std_logic_vector(to_unsigned(8,8) ,
44254	 => std_logic_vector(to_unsigned(10,8) ,
44255	 => std_logic_vector(to_unsigned(12,8) ,
44256	 => std_logic_vector(to_unsigned(15,8) ,
44257	 => std_logic_vector(to_unsigned(10,8) ,
44258	 => std_logic_vector(to_unsigned(5,8) ,
44259	 => std_logic_vector(to_unsigned(8,8) ,
44260	 => std_logic_vector(to_unsigned(9,8) ,
44261	 => std_logic_vector(to_unsigned(3,8) ,
44262	 => std_logic_vector(to_unsigned(3,8) ,
44263	 => std_logic_vector(to_unsigned(17,8) ,
44264	 => std_logic_vector(to_unsigned(72,8) ,
44265	 => std_logic_vector(to_unsigned(93,8) ,
44266	 => std_logic_vector(to_unsigned(68,8) ,
44267	 => std_logic_vector(to_unsigned(59,8) ,
44268	 => std_logic_vector(to_unsigned(55,8) ,
44269	 => std_logic_vector(to_unsigned(62,8) ,
44270	 => std_logic_vector(to_unsigned(67,8) ,
44271	 => std_logic_vector(to_unsigned(69,8) ,
44272	 => std_logic_vector(to_unsigned(95,8) ,
44273	 => std_logic_vector(to_unsigned(107,8) ,
44274	 => std_logic_vector(to_unsigned(68,8) ,
44275	 => std_logic_vector(to_unsigned(67,8) ,
44276	 => std_logic_vector(to_unsigned(92,8) ,
44277	 => std_logic_vector(to_unsigned(90,8) ,
44278	 => std_logic_vector(to_unsigned(91,8) ,
44279	 => std_logic_vector(to_unsigned(91,8) ,
44280	 => std_logic_vector(to_unsigned(93,8) ,
44281	 => std_logic_vector(to_unsigned(85,8) ,
44282	 => std_logic_vector(to_unsigned(81,8) ,
44283	 => std_logic_vector(to_unsigned(77,8) ,
44284	 => std_logic_vector(to_unsigned(13,8) ,
44285	 => std_logic_vector(to_unsigned(3,8) ,
44286	 => std_logic_vector(to_unsigned(5,8) ,
44287	 => std_logic_vector(to_unsigned(3,8) ,
44288	 => std_logic_vector(to_unsigned(2,8) ,
44289	 => std_logic_vector(to_unsigned(15,8) ,
44290	 => std_logic_vector(to_unsigned(100,8) ,
44291	 => std_logic_vector(to_unsigned(114,8) ,
44292	 => std_logic_vector(to_unsigned(96,8) ,
44293	 => std_logic_vector(to_unsigned(105,8) ,
44294	 => std_logic_vector(to_unsigned(95,8) ,
44295	 => std_logic_vector(to_unsigned(80,8) ,
44296	 => std_logic_vector(to_unsigned(90,8) ,
44297	 => std_logic_vector(to_unsigned(86,8) ,
44298	 => std_logic_vector(to_unsigned(96,8) ,
44299	 => std_logic_vector(to_unsigned(108,8) ,
44300	 => std_logic_vector(to_unsigned(96,8) ,
44301	 => std_logic_vector(to_unsigned(84,8) ,
44302	 => std_logic_vector(to_unsigned(84,8) ,
44303	 => std_logic_vector(to_unsigned(76,8) ,
44304	 => std_logic_vector(to_unsigned(63,8) ,
44305	 => std_logic_vector(to_unsigned(62,8) ,
44306	 => std_logic_vector(to_unsigned(79,8) ,
44307	 => std_logic_vector(to_unsigned(73,8) ,
44308	 => std_logic_vector(to_unsigned(76,8) ,
44309	 => std_logic_vector(to_unsigned(92,8) ,
44310	 => std_logic_vector(to_unsigned(100,8) ,
44311	 => std_logic_vector(to_unsigned(97,8) ,
44312	 => std_logic_vector(to_unsigned(86,8) ,
44313	 => std_logic_vector(to_unsigned(92,8) ,
44314	 => std_logic_vector(to_unsigned(95,8) ,
44315	 => std_logic_vector(to_unsigned(100,8) ,
44316	 => std_logic_vector(to_unsigned(121,8) ,
44317	 => std_logic_vector(to_unsigned(141,8) ,
44318	 => std_logic_vector(to_unsigned(20,8) ,
44319	 => std_logic_vector(to_unsigned(0,8) ,
44320	 => std_logic_vector(to_unsigned(4,8) ,
44321	 => std_logic_vector(to_unsigned(3,8) ,
44322	 => std_logic_vector(to_unsigned(1,8) ,
44323	 => std_logic_vector(to_unsigned(13,8) ,
44324	 => std_logic_vector(to_unsigned(112,8) ,
44325	 => std_logic_vector(to_unsigned(122,8) ,
44326	 => std_logic_vector(to_unsigned(80,8) ,
44327	 => std_logic_vector(to_unsigned(60,8) ,
44328	 => std_logic_vector(to_unsigned(70,8) ,
44329	 => std_logic_vector(to_unsigned(103,8) ,
44330	 => std_logic_vector(to_unsigned(101,8) ,
44331	 => std_logic_vector(to_unsigned(96,8) ,
44332	 => std_logic_vector(to_unsigned(100,8) ,
44333	 => std_logic_vector(to_unsigned(108,8) ,
44334	 => std_logic_vector(to_unsigned(91,8) ,
44335	 => std_logic_vector(to_unsigned(59,8) ,
44336	 => std_logic_vector(to_unsigned(25,8) ,
44337	 => std_logic_vector(to_unsigned(2,8) ,
44338	 => std_logic_vector(to_unsigned(5,8) ,
44339	 => std_logic_vector(to_unsigned(5,8) ,
44340	 => std_logic_vector(to_unsigned(5,8) ,
44341	 => std_logic_vector(to_unsigned(3,8) ,
44342	 => std_logic_vector(to_unsigned(1,8) ,
44343	 => std_logic_vector(to_unsigned(47,8) ,
44344	 => std_logic_vector(to_unsigned(43,8) ,
44345	 => std_logic_vector(to_unsigned(5,8) ,
44346	 => std_logic_vector(to_unsigned(10,8) ,
44347	 => std_logic_vector(to_unsigned(21,8) ,
44348	 => std_logic_vector(to_unsigned(48,8) ,
44349	 => std_logic_vector(to_unsigned(13,8) ,
44350	 => std_logic_vector(to_unsigned(18,8) ,
44351	 => std_logic_vector(to_unsigned(121,8) ,
44352	 => std_logic_vector(to_unsigned(118,8) ,
44353	 => std_logic_vector(to_unsigned(108,8) ,
44354	 => std_logic_vector(to_unsigned(116,8) ,
44355	 => std_logic_vector(to_unsigned(108,8) ,
44356	 => std_logic_vector(to_unsigned(97,8) ,
44357	 => std_logic_vector(to_unsigned(107,8) ,
44358	 => std_logic_vector(to_unsigned(107,8) ,
44359	 => std_logic_vector(to_unsigned(80,8) ,
44360	 => std_logic_vector(to_unsigned(87,8) ,
44361	 => std_logic_vector(to_unsigned(130,8) ,
44362	 => std_logic_vector(to_unsigned(144,8) ,
44363	 => std_logic_vector(to_unsigned(125,8) ,
44364	 => std_logic_vector(to_unsigned(114,8) ,
44365	 => std_logic_vector(to_unsigned(97,8) ,
44366	 => std_logic_vector(to_unsigned(46,8) ,
44367	 => std_logic_vector(to_unsigned(19,8) ,
44368	 => std_logic_vector(to_unsigned(65,8) ,
44369	 => std_logic_vector(to_unsigned(29,8) ,
44370	 => std_logic_vector(to_unsigned(22,8) ,
44371	 => std_logic_vector(to_unsigned(3,8) ,
44372	 => std_logic_vector(to_unsigned(10,8) ,
44373	 => std_logic_vector(to_unsigned(39,8) ,
44374	 => std_logic_vector(to_unsigned(2,8) ,
44375	 => std_logic_vector(to_unsigned(1,8) ,
44376	 => std_logic_vector(to_unsigned(3,8) ,
44377	 => std_logic_vector(to_unsigned(21,8) ,
44378	 => std_logic_vector(to_unsigned(3,8) ,
44379	 => std_logic_vector(to_unsigned(3,8) ,
44380	 => std_logic_vector(to_unsigned(12,8) ,
44381	 => std_logic_vector(to_unsigned(8,8) ,
44382	 => std_logic_vector(to_unsigned(6,8) ,
44383	 => std_logic_vector(to_unsigned(5,8) ,
44384	 => std_logic_vector(to_unsigned(2,8) ,
44385	 => std_logic_vector(to_unsigned(1,8) ,
44386	 => std_logic_vector(to_unsigned(1,8) ,
44387	 => std_logic_vector(to_unsigned(1,8) ,
44388	 => std_logic_vector(to_unsigned(1,8) ,
44389	 => std_logic_vector(to_unsigned(1,8) ,
44390	 => std_logic_vector(to_unsigned(0,8) ,
44391	 => std_logic_vector(to_unsigned(1,8) ,
44392	 => std_logic_vector(to_unsigned(3,8) ,
44393	 => std_logic_vector(to_unsigned(5,8) ,
44394	 => std_logic_vector(to_unsigned(11,8) ,
44395	 => std_logic_vector(to_unsigned(1,8) ,
44396	 => std_logic_vector(to_unsigned(1,8) ,
44397	 => std_logic_vector(to_unsigned(1,8) ,
44398	 => std_logic_vector(to_unsigned(0,8) ,
44399	 => std_logic_vector(to_unsigned(0,8) ,
44400	 => std_logic_vector(to_unsigned(0,8) ,
44401	 => std_logic_vector(to_unsigned(1,8) ,
44402	 => std_logic_vector(to_unsigned(2,8) ,
44403	 => std_logic_vector(to_unsigned(2,8) ,
44404	 => std_logic_vector(to_unsigned(2,8) ,
44405	 => std_logic_vector(to_unsigned(1,8) ,
44406	 => std_logic_vector(to_unsigned(1,8) ,
44407	 => std_logic_vector(to_unsigned(1,8) ,
44408	 => std_logic_vector(to_unsigned(7,8) ,
44409	 => std_logic_vector(to_unsigned(8,8) ,
44410	 => std_logic_vector(to_unsigned(4,8) ,
44411	 => std_logic_vector(to_unsigned(4,8) ,
44412	 => std_logic_vector(to_unsigned(3,8) ,
44413	 => std_logic_vector(to_unsigned(3,8) ,
44414	 => std_logic_vector(to_unsigned(3,8) ,
44415	 => std_logic_vector(to_unsigned(2,8) ,
44416	 => std_logic_vector(to_unsigned(1,8) ,
44417	 => std_logic_vector(to_unsigned(1,8) ,
44418	 => std_logic_vector(to_unsigned(2,8) ,
44419	 => std_logic_vector(to_unsigned(3,8) ,
44420	 => std_logic_vector(to_unsigned(2,8) ,
44421	 => std_logic_vector(to_unsigned(1,8) ,
44422	 => std_logic_vector(to_unsigned(1,8) ,
44423	 => std_logic_vector(to_unsigned(19,8) ,
44424	 => std_logic_vector(to_unsigned(21,8) ,
44425	 => std_logic_vector(to_unsigned(40,8) ,
44426	 => std_logic_vector(to_unsigned(64,8) ,
44427	 => std_logic_vector(to_unsigned(23,8) ,
44428	 => std_logic_vector(to_unsigned(5,8) ,
44429	 => std_logic_vector(to_unsigned(20,8) ,
44430	 => std_logic_vector(to_unsigned(36,8) ,
44431	 => std_logic_vector(to_unsigned(16,8) ,
44432	 => std_logic_vector(to_unsigned(7,8) ,
44433	 => std_logic_vector(to_unsigned(4,8) ,
44434	 => std_logic_vector(to_unsigned(5,8) ,
44435	 => std_logic_vector(to_unsigned(10,8) ,
44436	 => std_logic_vector(to_unsigned(14,8) ,
44437	 => std_logic_vector(to_unsigned(2,8) ,
44438	 => std_logic_vector(to_unsigned(0,8) ,
44439	 => std_logic_vector(to_unsigned(0,8) ,
44440	 => std_logic_vector(to_unsigned(0,8) ,
44441	 => std_logic_vector(to_unsigned(0,8) ,
44442	 => std_logic_vector(to_unsigned(1,8) ,
44443	 => std_logic_vector(to_unsigned(3,8) ,
44444	 => std_logic_vector(to_unsigned(5,8) ,
44445	 => std_logic_vector(to_unsigned(4,8) ,
44446	 => std_logic_vector(to_unsigned(6,8) ,
44447	 => std_logic_vector(to_unsigned(5,8) ,
44448	 => std_logic_vector(to_unsigned(4,8) ,
44449	 => std_logic_vector(to_unsigned(7,8) ,
44450	 => std_logic_vector(to_unsigned(1,8) ,
44451	 => std_logic_vector(to_unsigned(0,8) ,
44452	 => std_logic_vector(to_unsigned(1,8) ,
44453	 => std_logic_vector(to_unsigned(1,8) ,
44454	 => std_logic_vector(to_unsigned(1,8) ,
44455	 => std_logic_vector(to_unsigned(1,8) ,
44456	 => std_logic_vector(to_unsigned(1,8) ,
44457	 => std_logic_vector(to_unsigned(1,8) ,
44458	 => std_logic_vector(to_unsigned(1,8) ,
44459	 => std_logic_vector(to_unsigned(2,8) ,
44460	 => std_logic_vector(to_unsigned(1,8) ,
44461	 => std_logic_vector(to_unsigned(1,8) ,
44462	 => std_logic_vector(to_unsigned(1,8) ,
44463	 => std_logic_vector(to_unsigned(1,8) ,
44464	 => std_logic_vector(to_unsigned(1,8) ,
44465	 => std_logic_vector(to_unsigned(1,8) ,
44466	 => std_logic_vector(to_unsigned(2,8) ,
44467	 => std_logic_vector(to_unsigned(1,8) ,
44468	 => std_logic_vector(to_unsigned(2,8) ,
44469	 => std_logic_vector(to_unsigned(2,8) ,
44470	 => std_logic_vector(to_unsigned(3,8) ,
44471	 => std_logic_vector(to_unsigned(2,8) ,
44472	 => std_logic_vector(to_unsigned(1,8) ,
44473	 => std_logic_vector(to_unsigned(2,8) ,
44474	 => std_logic_vector(to_unsigned(2,8) ,
44475	 => std_logic_vector(to_unsigned(2,8) ,
44476	 => std_logic_vector(to_unsigned(2,8) ,
44477	 => std_logic_vector(to_unsigned(2,8) ,
44478	 => std_logic_vector(to_unsigned(2,8) ,
44479	 => std_logic_vector(to_unsigned(2,8) ,
44480	 => std_logic_vector(to_unsigned(2,8) ,
44481	 => std_logic_vector(to_unsigned(66,8) ,
44482	 => std_logic_vector(to_unsigned(53,8) ,
44483	 => std_logic_vector(to_unsigned(60,8) ,
44484	 => std_logic_vector(to_unsigned(59,8) ,
44485	 => std_logic_vector(to_unsigned(61,8) ,
44486	 => std_logic_vector(to_unsigned(56,8) ,
44487	 => std_logic_vector(to_unsigned(61,8) ,
44488	 => std_logic_vector(to_unsigned(58,8) ,
44489	 => std_logic_vector(to_unsigned(36,8) ,
44490	 => std_logic_vector(to_unsigned(38,8) ,
44491	 => std_logic_vector(to_unsigned(38,8) ,
44492	 => std_logic_vector(to_unsigned(44,8) ,
44493	 => std_logic_vector(to_unsigned(53,8) ,
44494	 => std_logic_vector(to_unsigned(87,8) ,
44495	 => std_logic_vector(to_unsigned(115,8) ,
44496	 => std_logic_vector(to_unsigned(108,8) ,
44497	 => std_logic_vector(to_unsigned(111,8) ,
44498	 => std_logic_vector(to_unsigned(114,8) ,
44499	 => std_logic_vector(to_unsigned(115,8) ,
44500	 => std_logic_vector(to_unsigned(116,8) ,
44501	 => std_logic_vector(to_unsigned(116,8) ,
44502	 => std_logic_vector(to_unsigned(118,8) ,
44503	 => std_logic_vector(to_unsigned(136,8) ,
44504	 => std_logic_vector(to_unsigned(139,8) ,
44505	 => std_logic_vector(to_unsigned(134,8) ,
44506	 => std_logic_vector(to_unsigned(146,8) ,
44507	 => std_logic_vector(to_unsigned(154,8) ,
44508	 => std_logic_vector(to_unsigned(141,8) ,
44509	 => std_logic_vector(to_unsigned(134,8) ,
44510	 => std_logic_vector(to_unsigned(142,8) ,
44511	 => std_logic_vector(to_unsigned(138,8) ,
44512	 => std_logic_vector(to_unsigned(144,8) ,
44513	 => std_logic_vector(to_unsigned(151,8) ,
44514	 => std_logic_vector(to_unsigned(144,8) ,
44515	 => std_logic_vector(to_unsigned(151,8) ,
44516	 => std_logic_vector(to_unsigned(149,8) ,
44517	 => std_logic_vector(to_unsigned(151,8) ,
44518	 => std_logic_vector(to_unsigned(152,8) ,
44519	 => std_logic_vector(to_unsigned(156,8) ,
44520	 => std_logic_vector(to_unsigned(154,8) ,
44521	 => std_logic_vector(to_unsigned(93,8) ,
44522	 => std_logic_vector(to_unsigned(91,8) ,
44523	 => std_logic_vector(to_unsigned(109,8) ,
44524	 => std_logic_vector(to_unsigned(114,8) ,
44525	 => std_logic_vector(to_unsigned(109,8) ,
44526	 => std_logic_vector(to_unsigned(77,8) ,
44527	 => std_logic_vector(to_unsigned(80,8) ,
44528	 => std_logic_vector(to_unsigned(85,8) ,
44529	 => std_logic_vector(to_unsigned(86,8) ,
44530	 => std_logic_vector(to_unsigned(111,8) ,
44531	 => std_logic_vector(to_unsigned(115,8) ,
44532	 => std_logic_vector(to_unsigned(119,8) ,
44533	 => std_logic_vector(to_unsigned(133,8) ,
44534	 => std_logic_vector(to_unsigned(133,8) ,
44535	 => std_logic_vector(to_unsigned(125,8) ,
44536	 => std_logic_vector(to_unsigned(115,8) ,
44537	 => std_logic_vector(to_unsigned(104,8) ,
44538	 => std_logic_vector(to_unsigned(95,8) ,
44539	 => std_logic_vector(to_unsigned(92,8) ,
44540	 => std_logic_vector(to_unsigned(85,8) ,
44541	 => std_logic_vector(to_unsigned(80,8) ,
44542	 => std_logic_vector(to_unsigned(93,8) ,
44543	 => std_logic_vector(to_unsigned(90,8) ,
44544	 => std_logic_vector(to_unsigned(86,8) ,
44545	 => std_logic_vector(to_unsigned(95,8) ,
44546	 => std_logic_vector(to_unsigned(101,8) ,
44547	 => std_logic_vector(to_unsigned(93,8) ,
44548	 => std_logic_vector(to_unsigned(84,8) ,
44549	 => std_logic_vector(to_unsigned(81,8) ,
44550	 => std_logic_vector(to_unsigned(86,8) ,
44551	 => std_logic_vector(to_unsigned(78,8) ,
44552	 => std_logic_vector(to_unsigned(72,8) ,
44553	 => std_logic_vector(to_unsigned(70,8) ,
44554	 => std_logic_vector(to_unsigned(70,8) ,
44555	 => std_logic_vector(to_unsigned(84,8) ,
44556	 => std_logic_vector(to_unsigned(90,8) ,
44557	 => std_logic_vector(to_unsigned(101,8) ,
44558	 => std_logic_vector(to_unsigned(112,8) ,
44559	 => std_logic_vector(to_unsigned(112,8) ,
44560	 => std_logic_vector(to_unsigned(86,8) ,
44561	 => std_logic_vector(to_unsigned(82,8) ,
44562	 => std_logic_vector(to_unsigned(80,8) ,
44563	 => std_logic_vector(to_unsigned(93,8) ,
44564	 => std_logic_vector(to_unsigned(111,8) ,
44565	 => std_logic_vector(to_unsigned(112,8) ,
44566	 => std_logic_vector(to_unsigned(95,8) ,
44567	 => std_logic_vector(to_unsigned(85,8) ,
44568	 => std_logic_vector(to_unsigned(86,8) ,
44569	 => std_logic_vector(to_unsigned(30,8) ,
44570	 => std_logic_vector(to_unsigned(3,8) ,
44571	 => std_logic_vector(to_unsigned(5,8) ,
44572	 => std_logic_vector(to_unsigned(18,8) ,
44573	 => std_logic_vector(to_unsigned(15,8) ,
44574	 => std_logic_vector(to_unsigned(20,8) ,
44575	 => std_logic_vector(to_unsigned(36,8) ,
44576	 => std_logic_vector(to_unsigned(58,8) ,
44577	 => std_logic_vector(to_unsigned(25,8) ,
44578	 => std_logic_vector(to_unsigned(5,8) ,
44579	 => std_logic_vector(to_unsigned(8,8) ,
44580	 => std_logic_vector(to_unsigned(11,8) ,
44581	 => std_logic_vector(to_unsigned(21,8) ,
44582	 => std_logic_vector(to_unsigned(57,8) ,
44583	 => std_logic_vector(to_unsigned(79,8) ,
44584	 => std_logic_vector(to_unsigned(97,8) ,
44585	 => std_logic_vector(to_unsigned(101,8) ,
44586	 => std_logic_vector(to_unsigned(73,8) ,
44587	 => std_logic_vector(to_unsigned(56,8) ,
44588	 => std_logic_vector(to_unsigned(57,8) ,
44589	 => std_logic_vector(to_unsigned(65,8) ,
44590	 => std_logic_vector(to_unsigned(63,8) ,
44591	 => std_logic_vector(to_unsigned(65,8) ,
44592	 => std_logic_vector(to_unsigned(87,8) ,
44593	 => std_logic_vector(to_unsigned(81,8) ,
44594	 => std_logic_vector(to_unsigned(62,8) ,
44595	 => std_logic_vector(to_unsigned(65,8) ,
44596	 => std_logic_vector(to_unsigned(67,8) ,
44597	 => std_logic_vector(to_unsigned(69,8) ,
44598	 => std_logic_vector(to_unsigned(82,8) ,
44599	 => std_logic_vector(to_unsigned(85,8) ,
44600	 => std_logic_vector(to_unsigned(87,8) ,
44601	 => std_logic_vector(to_unsigned(82,8) ,
44602	 => std_logic_vector(to_unsigned(91,8) ,
44603	 => std_logic_vector(to_unsigned(47,8) ,
44604	 => std_logic_vector(to_unsigned(5,8) ,
44605	 => std_logic_vector(to_unsigned(6,8) ,
44606	 => std_logic_vector(to_unsigned(6,8) ,
44607	 => std_logic_vector(to_unsigned(6,8) ,
44608	 => std_logic_vector(to_unsigned(5,8) ,
44609	 => std_logic_vector(to_unsigned(14,8) ,
44610	 => std_logic_vector(to_unsigned(95,8) ,
44611	 => std_logic_vector(to_unsigned(118,8) ,
44612	 => std_logic_vector(to_unsigned(127,8) ,
44613	 => std_logic_vector(to_unsigned(112,8) ,
44614	 => std_logic_vector(to_unsigned(100,8) ,
44615	 => std_logic_vector(to_unsigned(101,8) ,
44616	 => std_logic_vector(to_unsigned(105,8) ,
44617	 => std_logic_vector(to_unsigned(78,8) ,
44618	 => std_logic_vector(to_unsigned(88,8) ,
44619	 => std_logic_vector(to_unsigned(97,8) ,
44620	 => std_logic_vector(to_unsigned(86,8) ,
44621	 => std_logic_vector(to_unsigned(73,8) ,
44622	 => std_logic_vector(to_unsigned(69,8) ,
44623	 => std_logic_vector(to_unsigned(69,8) ,
44624	 => std_logic_vector(to_unsigned(62,8) ,
44625	 => std_logic_vector(to_unsigned(58,8) ,
44626	 => std_logic_vector(to_unsigned(68,8) ,
44627	 => std_logic_vector(to_unsigned(64,8) ,
44628	 => std_logic_vector(to_unsigned(65,8) ,
44629	 => std_logic_vector(to_unsigned(67,8) ,
44630	 => std_logic_vector(to_unsigned(68,8) ,
44631	 => std_logic_vector(to_unsigned(82,8) ,
44632	 => std_logic_vector(to_unsigned(81,8) ,
44633	 => std_logic_vector(to_unsigned(90,8) ,
44634	 => std_logic_vector(to_unsigned(79,8) ,
44635	 => std_logic_vector(to_unsigned(115,8) ,
44636	 => std_logic_vector(to_unsigned(157,8) ,
44637	 => std_logic_vector(to_unsigned(144,8) ,
44638	 => std_logic_vector(to_unsigned(63,8) ,
44639	 => std_logic_vector(to_unsigned(8,8) ,
44640	 => std_logic_vector(to_unsigned(3,8) ,
44641	 => std_logic_vector(to_unsigned(3,8) ,
44642	 => std_logic_vector(to_unsigned(15,8) ,
44643	 => std_logic_vector(to_unsigned(88,8) ,
44644	 => std_logic_vector(to_unsigned(128,8) ,
44645	 => std_logic_vector(to_unsigned(124,8) ,
44646	 => std_logic_vector(to_unsigned(56,8) ,
44647	 => std_logic_vector(to_unsigned(29,8) ,
44648	 => std_logic_vector(to_unsigned(41,8) ,
44649	 => std_logic_vector(to_unsigned(66,8) ,
44650	 => std_logic_vector(to_unsigned(86,8) ,
44651	 => std_logic_vector(to_unsigned(93,8) ,
44652	 => std_logic_vector(to_unsigned(77,8) ,
44653	 => std_logic_vector(to_unsigned(76,8) ,
44654	 => std_logic_vector(to_unsigned(79,8) ,
44655	 => std_logic_vector(to_unsigned(52,8) ,
44656	 => std_logic_vector(to_unsigned(16,8) ,
44657	 => std_logic_vector(to_unsigned(1,8) ,
44658	 => std_logic_vector(to_unsigned(4,8) ,
44659	 => std_logic_vector(to_unsigned(6,8) ,
44660	 => std_logic_vector(to_unsigned(4,8) ,
44661	 => std_logic_vector(to_unsigned(0,8) ,
44662	 => std_logic_vector(to_unsigned(11,8) ,
44663	 => std_logic_vector(to_unsigned(93,8) ,
44664	 => std_logic_vector(to_unsigned(20,8) ,
44665	 => std_logic_vector(to_unsigned(6,8) ,
44666	 => std_logic_vector(to_unsigned(12,8) ,
44667	 => std_logic_vector(to_unsigned(23,8) ,
44668	 => std_logic_vector(to_unsigned(31,8) ,
44669	 => std_logic_vector(to_unsigned(7,8) ,
44670	 => std_logic_vector(to_unsigned(21,8) ,
44671	 => std_logic_vector(to_unsigned(105,8) ,
44672	 => std_logic_vector(to_unsigned(84,8) ,
44673	 => std_logic_vector(to_unsigned(76,8) ,
44674	 => std_logic_vector(to_unsigned(100,8) ,
44675	 => std_logic_vector(to_unsigned(93,8) ,
44676	 => std_logic_vector(to_unsigned(77,8) ,
44677	 => std_logic_vector(to_unsigned(97,8) ,
44678	 => std_logic_vector(to_unsigned(111,8) ,
44679	 => std_logic_vector(to_unsigned(103,8) ,
44680	 => std_logic_vector(to_unsigned(118,8) ,
44681	 => std_logic_vector(to_unsigned(128,8) ,
44682	 => std_logic_vector(to_unsigned(142,8) ,
44683	 => std_logic_vector(to_unsigned(119,8) ,
44684	 => std_logic_vector(to_unsigned(72,8) ,
44685	 => std_logic_vector(to_unsigned(78,8) ,
44686	 => std_logic_vector(to_unsigned(32,8) ,
44687	 => std_logic_vector(to_unsigned(13,8) ,
44688	 => std_logic_vector(to_unsigned(51,8) ,
44689	 => std_logic_vector(to_unsigned(42,8) ,
44690	 => std_logic_vector(to_unsigned(21,8) ,
44691	 => std_logic_vector(to_unsigned(5,8) ,
44692	 => std_logic_vector(to_unsigned(19,8) ,
44693	 => std_logic_vector(to_unsigned(27,8) ,
44694	 => std_logic_vector(to_unsigned(1,8) ,
44695	 => std_logic_vector(to_unsigned(1,8) ,
44696	 => std_logic_vector(to_unsigned(2,8) ,
44697	 => std_logic_vector(to_unsigned(10,8) ,
44698	 => std_logic_vector(to_unsigned(1,8) ,
44699	 => std_logic_vector(to_unsigned(31,8) ,
44700	 => std_logic_vector(to_unsigned(112,8) ,
44701	 => std_logic_vector(to_unsigned(80,8) ,
44702	 => std_logic_vector(to_unsigned(76,8) ,
44703	 => std_logic_vector(to_unsigned(68,8) ,
44704	 => std_logic_vector(to_unsigned(56,8) ,
44705	 => std_logic_vector(to_unsigned(46,8) ,
44706	 => std_logic_vector(to_unsigned(34,8) ,
44707	 => std_logic_vector(to_unsigned(29,8) ,
44708	 => std_logic_vector(to_unsigned(21,8) ,
44709	 => std_logic_vector(to_unsigned(16,8) ,
44710	 => std_logic_vector(to_unsigned(11,8) ,
44711	 => std_logic_vector(to_unsigned(3,8) ,
44712	 => std_logic_vector(to_unsigned(2,8) ,
44713	 => std_logic_vector(to_unsigned(5,8) ,
44714	 => std_logic_vector(to_unsigned(18,8) ,
44715	 => std_logic_vector(to_unsigned(4,8) ,
44716	 => std_logic_vector(to_unsigned(1,8) ,
44717	 => std_logic_vector(to_unsigned(0,8) ,
44718	 => std_logic_vector(to_unsigned(0,8) ,
44719	 => std_logic_vector(to_unsigned(1,8) ,
44720	 => std_logic_vector(to_unsigned(1,8) ,
44721	 => std_logic_vector(to_unsigned(3,8) ,
44722	 => std_logic_vector(to_unsigned(12,8) ,
44723	 => std_logic_vector(to_unsigned(4,8) ,
44724	 => std_logic_vector(to_unsigned(1,8) ,
44725	 => std_logic_vector(to_unsigned(1,8) ,
44726	 => std_logic_vector(to_unsigned(0,8) ,
44727	 => std_logic_vector(to_unsigned(1,8) ,
44728	 => std_logic_vector(to_unsigned(7,8) ,
44729	 => std_logic_vector(to_unsigned(6,8) ,
44730	 => std_logic_vector(to_unsigned(5,8) ,
44731	 => std_logic_vector(to_unsigned(3,8) ,
44732	 => std_logic_vector(to_unsigned(3,8) ,
44733	 => std_logic_vector(to_unsigned(4,8) ,
44734	 => std_logic_vector(to_unsigned(3,8) ,
44735	 => std_logic_vector(to_unsigned(3,8) ,
44736	 => std_logic_vector(to_unsigned(3,8) ,
44737	 => std_logic_vector(to_unsigned(1,8) ,
44738	 => std_logic_vector(to_unsigned(0,8) ,
44739	 => std_logic_vector(to_unsigned(1,8) ,
44740	 => std_logic_vector(to_unsigned(1,8) ,
44741	 => std_logic_vector(to_unsigned(1,8) ,
44742	 => std_logic_vector(to_unsigned(0,8) ,
44743	 => std_logic_vector(to_unsigned(2,8) ,
44744	 => std_logic_vector(to_unsigned(17,8) ,
44745	 => std_logic_vector(to_unsigned(20,8) ,
44746	 => std_logic_vector(to_unsigned(15,8) ,
44747	 => std_logic_vector(to_unsigned(6,8) ,
44748	 => std_logic_vector(to_unsigned(1,8) ,
44749	 => std_logic_vector(to_unsigned(16,8) ,
44750	 => std_logic_vector(to_unsigned(40,8) ,
44751	 => std_logic_vector(to_unsigned(15,8) ,
44752	 => std_logic_vector(to_unsigned(9,8) ,
44753	 => std_logic_vector(to_unsigned(3,8) ,
44754	 => std_logic_vector(to_unsigned(5,8) ,
44755	 => std_logic_vector(to_unsigned(10,8) ,
44756	 => std_logic_vector(to_unsigned(19,8) ,
44757	 => std_logic_vector(to_unsigned(5,8) ,
44758	 => std_logic_vector(to_unsigned(1,8) ,
44759	 => std_logic_vector(to_unsigned(0,8) ,
44760	 => std_logic_vector(to_unsigned(0,8) ,
44761	 => std_logic_vector(to_unsigned(1,8) ,
44762	 => std_logic_vector(to_unsigned(2,8) ,
44763	 => std_logic_vector(to_unsigned(5,8) ,
44764	 => std_logic_vector(to_unsigned(6,8) ,
44765	 => std_logic_vector(to_unsigned(7,8) ,
44766	 => std_logic_vector(to_unsigned(8,8) ,
44767	 => std_logic_vector(to_unsigned(9,8) ,
44768	 => std_logic_vector(to_unsigned(11,8) ,
44769	 => std_logic_vector(to_unsigned(5,8) ,
44770	 => std_logic_vector(to_unsigned(0,8) ,
44771	 => std_logic_vector(to_unsigned(1,8) ,
44772	 => std_logic_vector(to_unsigned(1,8) ,
44773	 => std_logic_vector(to_unsigned(1,8) ,
44774	 => std_logic_vector(to_unsigned(1,8) ,
44775	 => std_logic_vector(to_unsigned(1,8) ,
44776	 => std_logic_vector(to_unsigned(1,8) ,
44777	 => std_logic_vector(to_unsigned(1,8) ,
44778	 => std_logic_vector(to_unsigned(2,8) ,
44779	 => std_logic_vector(to_unsigned(1,8) ,
44780	 => std_logic_vector(to_unsigned(1,8) ,
44781	 => std_logic_vector(to_unsigned(1,8) ,
44782	 => std_logic_vector(to_unsigned(1,8) ,
44783	 => std_logic_vector(to_unsigned(1,8) ,
44784	 => std_logic_vector(to_unsigned(1,8) ,
44785	 => std_logic_vector(to_unsigned(2,8) ,
44786	 => std_logic_vector(to_unsigned(2,8) ,
44787	 => std_logic_vector(to_unsigned(2,8) ,
44788	 => std_logic_vector(to_unsigned(1,8) ,
44789	 => std_logic_vector(to_unsigned(1,8) ,
44790	 => std_logic_vector(to_unsigned(2,8) ,
44791	 => std_logic_vector(to_unsigned(1,8) ,
44792	 => std_logic_vector(to_unsigned(2,8) ,
44793	 => std_logic_vector(to_unsigned(2,8) ,
44794	 => std_logic_vector(to_unsigned(2,8) ,
44795	 => std_logic_vector(to_unsigned(2,8) ,
44796	 => std_logic_vector(to_unsigned(1,8) ,
44797	 => std_logic_vector(to_unsigned(2,8) ,
44798	 => std_logic_vector(to_unsigned(2,8) ,
44799	 => std_logic_vector(to_unsigned(2,8) ,
44800	 => std_logic_vector(to_unsigned(2,8) ,
44801	 => std_logic_vector(to_unsigned(63,8) ,
44802	 => std_logic_vector(to_unsigned(60,8) ,
44803	 => std_logic_vector(to_unsigned(68,8) ,
44804	 => std_logic_vector(to_unsigned(65,8) ,
44805	 => std_logic_vector(to_unsigned(64,8) ,
44806	 => std_logic_vector(to_unsigned(61,8) ,
44807	 => std_logic_vector(to_unsigned(63,8) ,
44808	 => std_logic_vector(to_unsigned(56,8) ,
44809	 => std_logic_vector(to_unsigned(32,8) ,
44810	 => std_logic_vector(to_unsigned(34,8) ,
44811	 => std_logic_vector(to_unsigned(37,8) ,
44812	 => std_logic_vector(to_unsigned(42,8) ,
44813	 => std_logic_vector(to_unsigned(46,8) ,
44814	 => std_logic_vector(to_unsigned(71,8) ,
44815	 => std_logic_vector(to_unsigned(115,8) ,
44816	 => std_logic_vector(to_unsigned(115,8) ,
44817	 => std_logic_vector(to_unsigned(116,8) ,
44818	 => std_logic_vector(to_unsigned(121,8) ,
44819	 => std_logic_vector(to_unsigned(121,8) ,
44820	 => std_logic_vector(to_unsigned(124,8) ,
44821	 => std_logic_vector(to_unsigned(121,8) ,
44822	 => std_logic_vector(to_unsigned(121,8) ,
44823	 => std_logic_vector(to_unsigned(131,8) ,
44824	 => std_logic_vector(to_unsigned(134,8) ,
44825	 => std_logic_vector(to_unsigned(121,8) ,
44826	 => std_logic_vector(to_unsigned(125,8) ,
44827	 => std_logic_vector(to_unsigned(133,8) ,
44828	 => std_logic_vector(to_unsigned(119,8) ,
44829	 => std_logic_vector(to_unsigned(122,8) ,
44830	 => std_logic_vector(to_unsigned(144,8) ,
44831	 => std_logic_vector(to_unsigned(146,8) ,
44832	 => std_logic_vector(to_unsigned(144,8) ,
44833	 => std_logic_vector(to_unsigned(157,8) ,
44834	 => std_logic_vector(to_unsigned(124,8) ,
44835	 => std_logic_vector(to_unsigned(124,8) ,
44836	 => std_logic_vector(to_unsigned(154,8) ,
44837	 => std_logic_vector(to_unsigned(152,8) ,
44838	 => std_logic_vector(to_unsigned(154,8) ,
44839	 => std_logic_vector(to_unsigned(147,8) ,
44840	 => std_logic_vector(to_unsigned(147,8) ,
44841	 => std_logic_vector(to_unsigned(127,8) ,
44842	 => std_logic_vector(to_unsigned(114,8) ,
44843	 => std_logic_vector(to_unsigned(114,8) ,
44844	 => std_logic_vector(to_unsigned(99,8) ,
44845	 => std_logic_vector(to_unsigned(88,8) ,
44846	 => std_logic_vector(to_unsigned(78,8) ,
44847	 => std_logic_vector(to_unsigned(71,8) ,
44848	 => std_logic_vector(to_unsigned(74,8) ,
44849	 => std_logic_vector(to_unsigned(81,8) ,
44850	 => std_logic_vector(to_unsigned(104,8) ,
44851	 => std_logic_vector(to_unsigned(115,8) ,
44852	 => std_logic_vector(to_unsigned(130,8) ,
44853	 => std_logic_vector(to_unsigned(142,8) ,
44854	 => std_logic_vector(to_unsigned(142,8) ,
44855	 => std_logic_vector(to_unsigned(133,8) ,
44856	 => std_logic_vector(to_unsigned(136,8) ,
44857	 => std_logic_vector(to_unsigned(127,8) ,
44858	 => std_logic_vector(to_unsigned(107,8) ,
44859	 => std_logic_vector(to_unsigned(111,8) ,
44860	 => std_logic_vector(to_unsigned(115,8) ,
44861	 => std_logic_vector(to_unsigned(112,8) ,
44862	 => std_logic_vector(to_unsigned(91,8) ,
44863	 => std_logic_vector(to_unsigned(85,8) ,
44864	 => std_logic_vector(to_unsigned(85,8) ,
44865	 => std_logic_vector(to_unsigned(86,8) ,
44866	 => std_logic_vector(to_unsigned(96,8) ,
44867	 => std_logic_vector(to_unsigned(91,8) ,
44868	 => std_logic_vector(to_unsigned(81,8) ,
44869	 => std_logic_vector(to_unsigned(80,8) ,
44870	 => std_logic_vector(to_unsigned(79,8) ,
44871	 => std_logic_vector(to_unsigned(73,8) ,
44872	 => std_logic_vector(to_unsigned(70,8) ,
44873	 => std_logic_vector(to_unsigned(65,8) ,
44874	 => std_logic_vector(to_unsigned(63,8) ,
44875	 => std_logic_vector(to_unsigned(78,8) ,
44876	 => std_logic_vector(to_unsigned(105,8) ,
44877	 => std_logic_vector(to_unsigned(101,8) ,
44878	 => std_logic_vector(to_unsigned(100,8) ,
44879	 => std_logic_vector(to_unsigned(104,8) ,
44880	 => std_logic_vector(to_unsigned(93,8) ,
44881	 => std_logic_vector(to_unsigned(86,8) ,
44882	 => std_logic_vector(to_unsigned(91,8) ,
44883	 => std_logic_vector(to_unsigned(105,8) ,
44884	 => std_logic_vector(to_unsigned(99,8) ,
44885	 => std_logic_vector(to_unsigned(91,8) ,
44886	 => std_logic_vector(to_unsigned(91,8) ,
44887	 => std_logic_vector(to_unsigned(80,8) ,
44888	 => std_logic_vector(to_unsigned(78,8) ,
44889	 => std_logic_vector(to_unsigned(74,8) ,
44890	 => std_logic_vector(to_unsigned(46,8) ,
44891	 => std_logic_vector(to_unsigned(41,8) ,
44892	 => std_logic_vector(to_unsigned(37,8) ,
44893	 => std_logic_vector(to_unsigned(46,8) ,
44894	 => std_logic_vector(to_unsigned(58,8) ,
44895	 => std_logic_vector(to_unsigned(68,8) ,
44896	 => std_logic_vector(to_unsigned(85,8) ,
44897	 => std_logic_vector(to_unsigned(62,8) ,
44898	 => std_logic_vector(to_unsigned(47,8) ,
44899	 => std_logic_vector(to_unsigned(51,8) ,
44900	 => std_logic_vector(to_unsigned(71,8) ,
44901	 => std_logic_vector(to_unsigned(88,8) ,
44902	 => std_logic_vector(to_unsigned(88,8) ,
44903	 => std_logic_vector(to_unsigned(91,8) ,
44904	 => std_logic_vector(to_unsigned(111,8) ,
44905	 => std_logic_vector(to_unsigned(124,8) ,
44906	 => std_logic_vector(to_unsigned(82,8) ,
44907	 => std_logic_vector(to_unsigned(60,8) ,
44908	 => std_logic_vector(to_unsigned(62,8) ,
44909	 => std_logic_vector(to_unsigned(67,8) ,
44910	 => std_logic_vector(to_unsigned(90,8) ,
44911	 => std_logic_vector(to_unsigned(82,8) ,
44912	 => std_logic_vector(to_unsigned(92,8) ,
44913	 => std_logic_vector(to_unsigned(88,8) ,
44914	 => std_logic_vector(to_unsigned(55,8) ,
44915	 => std_logic_vector(to_unsigned(62,8) ,
44916	 => std_logic_vector(to_unsigned(59,8) ,
44917	 => std_logic_vector(to_unsigned(58,8) ,
44918	 => std_logic_vector(to_unsigned(81,8) ,
44919	 => std_logic_vector(to_unsigned(71,8) ,
44920	 => std_logic_vector(to_unsigned(76,8) ,
44921	 => std_logic_vector(to_unsigned(76,8) ,
44922	 => std_logic_vector(to_unsigned(86,8) ,
44923	 => std_logic_vector(to_unsigned(19,8) ,
44924	 => std_logic_vector(to_unsigned(2,8) ,
44925	 => std_logic_vector(to_unsigned(5,8) ,
44926	 => std_logic_vector(to_unsigned(4,8) ,
44927	 => std_logic_vector(to_unsigned(7,8) ,
44928	 => std_logic_vector(to_unsigned(6,8) ,
44929	 => std_logic_vector(to_unsigned(9,8) ,
44930	 => std_logic_vector(to_unsigned(99,8) ,
44931	 => std_logic_vector(to_unsigned(130,8) ,
44932	 => std_logic_vector(to_unsigned(136,8) ,
44933	 => std_logic_vector(to_unsigned(122,8) ,
44934	 => std_logic_vector(to_unsigned(115,8) ,
44935	 => std_logic_vector(to_unsigned(119,8) ,
44936	 => std_logic_vector(to_unsigned(101,8) ,
44937	 => std_logic_vector(to_unsigned(72,8) ,
44938	 => std_logic_vector(to_unsigned(79,8) ,
44939	 => std_logic_vector(to_unsigned(91,8) ,
44940	 => std_logic_vector(to_unsigned(87,8) ,
44941	 => std_logic_vector(to_unsigned(73,8) ,
44942	 => std_logic_vector(to_unsigned(68,8) ,
44943	 => std_logic_vector(to_unsigned(66,8) ,
44944	 => std_logic_vector(to_unsigned(60,8) ,
44945	 => std_logic_vector(to_unsigned(52,8) ,
44946	 => std_logic_vector(to_unsigned(54,8) ,
44947	 => std_logic_vector(to_unsigned(52,8) ,
44948	 => std_logic_vector(to_unsigned(55,8) ,
44949	 => std_logic_vector(to_unsigned(53,8) ,
44950	 => std_logic_vector(to_unsigned(46,8) ,
44951	 => std_logic_vector(to_unsigned(70,8) ,
44952	 => std_logic_vector(to_unsigned(69,8) ,
44953	 => std_logic_vector(to_unsigned(61,8) ,
44954	 => std_logic_vector(to_unsigned(61,8) ,
44955	 => std_logic_vector(to_unsigned(76,8) ,
44956	 => std_logic_vector(to_unsigned(112,8) ,
44957	 => std_logic_vector(to_unsigned(114,8) ,
44958	 => std_logic_vector(to_unsigned(103,8) ,
44959	 => std_logic_vector(to_unsigned(84,8) ,
44960	 => std_logic_vector(to_unsigned(55,8) ,
44961	 => std_logic_vector(to_unsigned(54,8) ,
44962	 => std_logic_vector(to_unsigned(86,8) ,
44963	 => std_logic_vector(to_unsigned(107,8) ,
44964	 => std_logic_vector(to_unsigned(115,8) ,
44965	 => std_logic_vector(to_unsigned(131,8) ,
44966	 => std_logic_vector(to_unsigned(68,8) ,
44967	 => std_logic_vector(to_unsigned(20,8) ,
44968	 => std_logic_vector(to_unsigned(29,8) ,
44969	 => std_logic_vector(to_unsigned(41,8) ,
44970	 => std_logic_vector(to_unsigned(63,8) ,
44971	 => std_logic_vector(to_unsigned(56,8) ,
44972	 => std_logic_vector(to_unsigned(28,8) ,
44973	 => std_logic_vector(to_unsigned(32,8) ,
44974	 => std_logic_vector(to_unsigned(56,8) ,
44975	 => std_logic_vector(to_unsigned(62,8) ,
44976	 => std_logic_vector(to_unsigned(19,8) ,
44977	 => std_logic_vector(to_unsigned(0,8) ,
44978	 => std_logic_vector(to_unsigned(1,8) ,
44979	 => std_logic_vector(to_unsigned(2,8) ,
44980	 => std_logic_vector(to_unsigned(1,8) ,
44981	 => std_logic_vector(to_unsigned(6,8) ,
44982	 => std_logic_vector(to_unsigned(65,8) ,
44983	 => std_logic_vector(to_unsigned(84,8) ,
44984	 => std_logic_vector(to_unsigned(17,8) ,
44985	 => std_logic_vector(to_unsigned(12,8) ,
44986	 => std_logic_vector(to_unsigned(18,8) ,
44987	 => std_logic_vector(to_unsigned(23,8) ,
44988	 => std_logic_vector(to_unsigned(12,8) ,
44989	 => std_logic_vector(to_unsigned(2,8) ,
44990	 => std_logic_vector(to_unsigned(37,8) ,
44991	 => std_logic_vector(to_unsigned(112,8) ,
44992	 => std_logic_vector(to_unsigned(86,8) ,
44993	 => std_logic_vector(to_unsigned(82,8) ,
44994	 => std_logic_vector(to_unsigned(99,8) ,
44995	 => std_logic_vector(to_unsigned(86,8) ,
44996	 => std_logic_vector(to_unsigned(65,8) ,
44997	 => std_logic_vector(to_unsigned(86,8) ,
44998	 => std_logic_vector(to_unsigned(97,8) ,
44999	 => std_logic_vector(to_unsigned(65,8) ,
45000	 => std_logic_vector(to_unsigned(79,8) ,
45001	 => std_logic_vector(to_unsigned(124,8) ,
45002	 => std_logic_vector(to_unsigned(141,8) ,
45003	 => std_logic_vector(to_unsigned(95,8) ,
45004	 => std_logic_vector(to_unsigned(61,8) ,
45005	 => std_logic_vector(to_unsigned(68,8) ,
45006	 => std_logic_vector(to_unsigned(22,8) ,
45007	 => std_logic_vector(to_unsigned(15,8) ,
45008	 => std_logic_vector(to_unsigned(41,8) ,
45009	 => std_logic_vector(to_unsigned(50,8) ,
45010	 => std_logic_vector(to_unsigned(32,8) ,
45011	 => std_logic_vector(to_unsigned(8,8) ,
45012	 => std_logic_vector(to_unsigned(8,8) ,
45013	 => std_logic_vector(to_unsigned(6,8) ,
45014	 => std_logic_vector(to_unsigned(4,8) ,
45015	 => std_logic_vector(to_unsigned(4,8) ,
45016	 => std_logic_vector(to_unsigned(2,8) ,
45017	 => std_logic_vector(to_unsigned(4,8) ,
45018	 => std_logic_vector(to_unsigned(2,8) ,
45019	 => std_logic_vector(to_unsigned(62,8) ,
45020	 => std_logic_vector(to_unsigned(109,8) ,
45021	 => std_logic_vector(to_unsigned(95,8) ,
45022	 => std_logic_vector(to_unsigned(104,8) ,
45023	 => std_logic_vector(to_unsigned(93,8) ,
45024	 => std_logic_vector(to_unsigned(101,8) ,
45025	 => std_logic_vector(to_unsigned(99,8) ,
45026	 => std_logic_vector(to_unsigned(93,8) ,
45027	 => std_logic_vector(to_unsigned(101,8) ,
45028	 => std_logic_vector(to_unsigned(103,8) ,
45029	 => std_logic_vector(to_unsigned(101,8) ,
45030	 => std_logic_vector(to_unsigned(87,8) ,
45031	 => std_logic_vector(to_unsigned(13,8) ,
45032	 => std_logic_vector(to_unsigned(1,8) ,
45033	 => std_logic_vector(to_unsigned(2,8) ,
45034	 => std_logic_vector(to_unsigned(16,8) ,
45035	 => std_logic_vector(to_unsigned(6,8) ,
45036	 => std_logic_vector(to_unsigned(2,8) ,
45037	 => std_logic_vector(to_unsigned(5,8) ,
45038	 => std_logic_vector(to_unsigned(2,8) ,
45039	 => std_logic_vector(to_unsigned(2,8) ,
45040	 => std_logic_vector(to_unsigned(2,8) ,
45041	 => std_logic_vector(to_unsigned(6,8) ,
45042	 => std_logic_vector(to_unsigned(15,8) ,
45043	 => std_logic_vector(to_unsigned(3,8) ,
45044	 => std_logic_vector(to_unsigned(0,8) ,
45045	 => std_logic_vector(to_unsigned(0,8) ,
45046	 => std_logic_vector(to_unsigned(0,8) ,
45047	 => std_logic_vector(to_unsigned(1,8) ,
45048	 => std_logic_vector(to_unsigned(7,8) ,
45049	 => std_logic_vector(to_unsigned(5,8) ,
45050	 => std_logic_vector(to_unsigned(1,8) ,
45051	 => std_logic_vector(to_unsigned(1,8) ,
45052	 => std_logic_vector(to_unsigned(1,8) ,
45053	 => std_logic_vector(to_unsigned(1,8) ,
45054	 => std_logic_vector(to_unsigned(1,8) ,
45055	 => std_logic_vector(to_unsigned(1,8) ,
45056	 => std_logic_vector(to_unsigned(1,8) ,
45057	 => std_logic_vector(to_unsigned(1,8) ,
45058	 => std_logic_vector(to_unsigned(1,8) ,
45059	 => std_logic_vector(to_unsigned(1,8) ,
45060	 => std_logic_vector(to_unsigned(1,8) ,
45061	 => std_logic_vector(to_unsigned(0,8) ,
45062	 => std_logic_vector(to_unsigned(0,8) ,
45063	 => std_logic_vector(to_unsigned(0,8) ,
45064	 => std_logic_vector(to_unsigned(1,8) ,
45065	 => std_logic_vector(to_unsigned(1,8) ,
45066	 => std_logic_vector(to_unsigned(1,8) ,
45067	 => std_logic_vector(to_unsigned(3,8) ,
45068	 => std_logic_vector(to_unsigned(6,8) ,
45069	 => std_logic_vector(to_unsigned(6,8) ,
45070	 => std_logic_vector(to_unsigned(31,8) ,
45071	 => std_logic_vector(to_unsigned(20,8) ,
45072	 => std_logic_vector(to_unsigned(10,8) ,
45073	 => std_logic_vector(to_unsigned(4,8) ,
45074	 => std_logic_vector(to_unsigned(5,8) ,
45075	 => std_logic_vector(to_unsigned(7,8) ,
45076	 => std_logic_vector(to_unsigned(15,8) ,
45077	 => std_logic_vector(to_unsigned(5,8) ,
45078	 => std_logic_vector(to_unsigned(0,8) ,
45079	 => std_logic_vector(to_unsigned(0,8) ,
45080	 => std_logic_vector(to_unsigned(0,8) ,
45081	 => std_logic_vector(to_unsigned(0,8) ,
45082	 => std_logic_vector(to_unsigned(2,8) ,
45083	 => std_logic_vector(to_unsigned(4,8) ,
45084	 => std_logic_vector(to_unsigned(5,8) ,
45085	 => std_logic_vector(to_unsigned(7,8) ,
45086	 => std_logic_vector(to_unsigned(8,8) ,
45087	 => std_logic_vector(to_unsigned(10,8) ,
45088	 => std_logic_vector(to_unsigned(12,8) ,
45089	 => std_logic_vector(to_unsigned(2,8) ,
45090	 => std_logic_vector(to_unsigned(0,8) ,
45091	 => std_logic_vector(to_unsigned(1,8) ,
45092	 => std_logic_vector(to_unsigned(1,8) ,
45093	 => std_logic_vector(to_unsigned(1,8) ,
45094	 => std_logic_vector(to_unsigned(1,8) ,
45095	 => std_logic_vector(to_unsigned(1,8) ,
45096	 => std_logic_vector(to_unsigned(1,8) ,
45097	 => std_logic_vector(to_unsigned(1,8) ,
45098	 => std_logic_vector(to_unsigned(2,8) ,
45099	 => std_logic_vector(to_unsigned(2,8) ,
45100	 => std_logic_vector(to_unsigned(1,8) ,
45101	 => std_logic_vector(to_unsigned(2,8) ,
45102	 => std_logic_vector(to_unsigned(1,8) ,
45103	 => std_logic_vector(to_unsigned(1,8) ,
45104	 => std_logic_vector(to_unsigned(2,8) ,
45105	 => std_logic_vector(to_unsigned(2,8) ,
45106	 => std_logic_vector(to_unsigned(2,8) ,
45107	 => std_logic_vector(to_unsigned(2,8) ,
45108	 => std_logic_vector(to_unsigned(2,8) ,
45109	 => std_logic_vector(to_unsigned(1,8) ,
45110	 => std_logic_vector(to_unsigned(2,8) ,
45111	 => std_logic_vector(to_unsigned(1,8) ,
45112	 => std_logic_vector(to_unsigned(2,8) ,
45113	 => std_logic_vector(to_unsigned(3,8) ,
45114	 => std_logic_vector(to_unsigned(2,8) ,
45115	 => std_logic_vector(to_unsigned(2,8) ,
45116	 => std_logic_vector(to_unsigned(2,8) ,
45117	 => std_logic_vector(to_unsigned(2,8) ,
45118	 => std_logic_vector(to_unsigned(3,8) ,
45119	 => std_logic_vector(to_unsigned(2,8) ,
45120	 => std_logic_vector(to_unsigned(2,8) ,
45121	 => std_logic_vector(to_unsigned(63,8) ,
45122	 => std_logic_vector(to_unsigned(64,8) ,
45123	 => std_logic_vector(to_unsigned(65,8) ,
45124	 => std_logic_vector(to_unsigned(60,8) ,
45125	 => std_logic_vector(to_unsigned(61,8) ,
45126	 => std_logic_vector(to_unsigned(67,8) ,
45127	 => std_logic_vector(to_unsigned(69,8) ,
45128	 => std_logic_vector(to_unsigned(56,8) ,
45129	 => std_logic_vector(to_unsigned(34,8) ,
45130	 => std_logic_vector(to_unsigned(35,8) ,
45131	 => std_logic_vector(to_unsigned(38,8) ,
45132	 => std_logic_vector(to_unsigned(40,8) ,
45133	 => std_logic_vector(to_unsigned(41,8) ,
45134	 => std_logic_vector(to_unsigned(62,8) ,
45135	 => std_logic_vector(to_unsigned(122,8) ,
45136	 => std_logic_vector(to_unsigned(122,8) ,
45137	 => std_logic_vector(to_unsigned(112,8) ,
45138	 => std_logic_vector(to_unsigned(109,8) ,
45139	 => std_logic_vector(to_unsigned(112,8) ,
45140	 => std_logic_vector(to_unsigned(121,8) ,
45141	 => std_logic_vector(to_unsigned(121,8) ,
45142	 => std_logic_vector(to_unsigned(128,8) ,
45143	 => std_logic_vector(to_unsigned(127,8) ,
45144	 => std_logic_vector(to_unsigned(130,8) ,
45145	 => std_logic_vector(to_unsigned(133,8) ,
45146	 => std_logic_vector(to_unsigned(139,8) ,
45147	 => std_logic_vector(to_unsigned(138,8) ,
45148	 => std_logic_vector(to_unsigned(128,8) ,
45149	 => std_logic_vector(to_unsigned(138,8) ,
45150	 => std_logic_vector(to_unsigned(144,8) ,
45151	 => std_logic_vector(to_unsigned(133,8) ,
45152	 => std_logic_vector(to_unsigned(141,8) ,
45153	 => std_logic_vector(to_unsigned(152,8) ,
45154	 => std_logic_vector(to_unsigned(134,8) ,
45155	 => std_logic_vector(to_unsigned(130,8) ,
45156	 => std_logic_vector(to_unsigned(154,8) ,
45157	 => std_logic_vector(to_unsigned(152,8) ,
45158	 => std_logic_vector(to_unsigned(147,8) ,
45159	 => std_logic_vector(to_unsigned(149,8) ,
45160	 => std_logic_vector(to_unsigned(154,8) ,
45161	 => std_logic_vector(to_unsigned(115,8) ,
45162	 => std_logic_vector(to_unsigned(71,8) ,
45163	 => std_logic_vector(to_unsigned(85,8) ,
45164	 => std_logic_vector(to_unsigned(85,8) ,
45165	 => std_logic_vector(to_unsigned(80,8) ,
45166	 => std_logic_vector(to_unsigned(87,8) ,
45167	 => std_logic_vector(to_unsigned(79,8) ,
45168	 => std_logic_vector(to_unsigned(87,8) ,
45169	 => std_logic_vector(to_unsigned(85,8) ,
45170	 => std_logic_vector(to_unsigned(92,8) ,
45171	 => std_logic_vector(to_unsigned(109,8) ,
45172	 => std_logic_vector(to_unsigned(133,8) ,
45173	 => std_logic_vector(to_unsigned(144,8) ,
45174	 => std_logic_vector(to_unsigned(136,8) ,
45175	 => std_logic_vector(to_unsigned(112,8) ,
45176	 => std_logic_vector(to_unsigned(107,8) ,
45177	 => std_logic_vector(to_unsigned(115,8) ,
45178	 => std_logic_vector(to_unsigned(115,8) ,
45179	 => std_logic_vector(to_unsigned(119,8) ,
45180	 => std_logic_vector(to_unsigned(144,8) ,
45181	 => std_logic_vector(to_unsigned(147,8) ,
45182	 => std_logic_vector(to_unsigned(86,8) ,
45183	 => std_logic_vector(to_unsigned(77,8) ,
45184	 => std_logic_vector(to_unsigned(84,8) ,
45185	 => std_logic_vector(to_unsigned(82,8) ,
45186	 => std_logic_vector(to_unsigned(87,8) ,
45187	 => std_logic_vector(to_unsigned(81,8) ,
45188	 => std_logic_vector(to_unsigned(79,8) ,
45189	 => std_logic_vector(to_unsigned(81,8) ,
45190	 => std_logic_vector(to_unsigned(81,8) ,
45191	 => std_logic_vector(to_unsigned(73,8) ,
45192	 => std_logic_vector(to_unsigned(66,8) ,
45193	 => std_logic_vector(to_unsigned(60,8) ,
45194	 => std_logic_vector(to_unsigned(62,8) ,
45195	 => std_logic_vector(to_unsigned(71,8) ,
45196	 => std_logic_vector(to_unsigned(93,8) ,
45197	 => std_logic_vector(to_unsigned(100,8) ,
45198	 => std_logic_vector(to_unsigned(93,8) ,
45199	 => std_logic_vector(to_unsigned(101,8) ,
45200	 => std_logic_vector(to_unsigned(115,8) ,
45201	 => std_logic_vector(to_unsigned(97,8) ,
45202	 => std_logic_vector(to_unsigned(85,8) ,
45203	 => std_logic_vector(to_unsigned(87,8) ,
45204	 => std_logic_vector(to_unsigned(87,8) ,
45205	 => std_logic_vector(to_unsigned(87,8) ,
45206	 => std_logic_vector(to_unsigned(96,8) ,
45207	 => std_logic_vector(to_unsigned(78,8) ,
45208	 => std_logic_vector(to_unsigned(66,8) ,
45209	 => std_logic_vector(to_unsigned(69,8) ,
45210	 => std_logic_vector(to_unsigned(82,8) ,
45211	 => std_logic_vector(to_unsigned(86,8) ,
45212	 => std_logic_vector(to_unsigned(73,8) ,
45213	 => std_logic_vector(to_unsigned(80,8) ,
45214	 => std_logic_vector(to_unsigned(84,8) ,
45215	 => std_logic_vector(to_unsigned(78,8) ,
45216	 => std_logic_vector(to_unsigned(72,8) ,
45217	 => std_logic_vector(to_unsigned(66,8) ,
45218	 => std_logic_vector(to_unsigned(77,8) ,
45219	 => std_logic_vector(to_unsigned(88,8) ,
45220	 => std_logic_vector(to_unsigned(80,8) ,
45221	 => std_logic_vector(to_unsigned(78,8) ,
45222	 => std_logic_vector(to_unsigned(72,8) ,
45223	 => std_logic_vector(to_unsigned(72,8) ,
45224	 => std_logic_vector(to_unsigned(101,8) ,
45225	 => std_logic_vector(to_unsigned(85,8) ,
45226	 => std_logic_vector(to_unsigned(62,8) ,
45227	 => std_logic_vector(to_unsigned(79,8) ,
45228	 => std_logic_vector(to_unsigned(71,8) ,
45229	 => std_logic_vector(to_unsigned(73,8) ,
45230	 => std_logic_vector(to_unsigned(95,8) ,
45231	 => std_logic_vector(to_unsigned(91,8) ,
45232	 => std_logic_vector(to_unsigned(88,8) ,
45233	 => std_logic_vector(to_unsigned(78,8) ,
45234	 => std_logic_vector(to_unsigned(54,8) ,
45235	 => std_logic_vector(to_unsigned(62,8) ,
45236	 => std_logic_vector(to_unsigned(84,8) ,
45237	 => std_logic_vector(to_unsigned(80,8) ,
45238	 => std_logic_vector(to_unsigned(81,8) ,
45239	 => std_logic_vector(to_unsigned(76,8) ,
45240	 => std_logic_vector(to_unsigned(72,8) ,
45241	 => std_logic_vector(to_unsigned(82,8) ,
45242	 => std_logic_vector(to_unsigned(79,8) ,
45243	 => std_logic_vector(to_unsigned(16,8) ,
45244	 => std_logic_vector(to_unsigned(7,8) ,
45245	 => std_logic_vector(to_unsigned(7,8) ,
45246	 => std_logic_vector(to_unsigned(6,8) ,
45247	 => std_logic_vector(to_unsigned(11,8) ,
45248	 => std_logic_vector(to_unsigned(3,8) ,
45249	 => std_logic_vector(to_unsigned(25,8) ,
45250	 => std_logic_vector(to_unsigned(128,8) ,
45251	 => std_logic_vector(to_unsigned(108,8) ,
45252	 => std_logic_vector(to_unsigned(139,8) ,
45253	 => std_logic_vector(to_unsigned(141,8) ,
45254	 => std_logic_vector(to_unsigned(136,8) ,
45255	 => std_logic_vector(to_unsigned(122,8) ,
45256	 => std_logic_vector(to_unsigned(92,8) ,
45257	 => std_logic_vector(to_unsigned(70,8) ,
45258	 => std_logic_vector(to_unsigned(81,8) ,
45259	 => std_logic_vector(to_unsigned(99,8) ,
45260	 => std_logic_vector(to_unsigned(86,8) ,
45261	 => std_logic_vector(to_unsigned(68,8) ,
45262	 => std_logic_vector(to_unsigned(73,8) ,
45263	 => std_logic_vector(to_unsigned(64,8) ,
45264	 => std_logic_vector(to_unsigned(57,8) ,
45265	 => std_logic_vector(to_unsigned(52,8) ,
45266	 => std_logic_vector(to_unsigned(50,8) ,
45267	 => std_logic_vector(to_unsigned(57,8) ,
45268	 => std_logic_vector(to_unsigned(60,8) ,
45269	 => std_logic_vector(to_unsigned(59,8) ,
45270	 => std_logic_vector(to_unsigned(59,8) ,
45271	 => std_logic_vector(to_unsigned(81,8) ,
45272	 => std_logic_vector(to_unsigned(65,8) ,
45273	 => std_logic_vector(to_unsigned(51,8) ,
45274	 => std_logic_vector(to_unsigned(31,8) ,
45275	 => std_logic_vector(to_unsigned(25,8) ,
45276	 => std_logic_vector(to_unsigned(54,8) ,
45277	 => std_logic_vector(to_unsigned(92,8) ,
45278	 => std_logic_vector(to_unsigned(71,8) ,
45279	 => std_logic_vector(to_unsigned(81,8) ,
45280	 => std_logic_vector(to_unsigned(95,8) ,
45281	 => std_logic_vector(to_unsigned(100,8) ,
45282	 => std_logic_vector(to_unsigned(71,8) ,
45283	 => std_logic_vector(to_unsigned(82,8) ,
45284	 => std_logic_vector(to_unsigned(77,8) ,
45285	 => std_logic_vector(to_unsigned(62,8) ,
45286	 => std_logic_vector(to_unsigned(60,8) ,
45287	 => std_logic_vector(to_unsigned(20,8) ,
45288	 => std_logic_vector(to_unsigned(37,8) ,
45289	 => std_logic_vector(to_unsigned(65,8) ,
45290	 => std_logic_vector(to_unsigned(79,8) ,
45291	 => std_logic_vector(to_unsigned(53,8) ,
45292	 => std_logic_vector(to_unsigned(14,8) ,
45293	 => std_logic_vector(to_unsigned(19,8) ,
45294	 => std_logic_vector(to_unsigned(48,8) ,
45295	 => std_logic_vector(to_unsigned(62,8) ,
45296	 => std_logic_vector(to_unsigned(42,8) ,
45297	 => std_logic_vector(to_unsigned(7,8) ,
45298	 => std_logic_vector(to_unsigned(3,8) ,
45299	 => std_logic_vector(to_unsigned(4,8) ,
45300	 => std_logic_vector(to_unsigned(15,8) ,
45301	 => std_logic_vector(to_unsigned(47,8) ,
45302	 => std_logic_vector(to_unsigned(82,8) ,
45303	 => std_logic_vector(to_unsigned(48,8) ,
45304	 => std_logic_vector(to_unsigned(8,8) ,
45305	 => std_logic_vector(to_unsigned(20,8) ,
45306	 => std_logic_vector(to_unsigned(22,8) ,
45307	 => std_logic_vector(to_unsigned(10,8) ,
45308	 => std_logic_vector(to_unsigned(3,8) ,
45309	 => std_logic_vector(to_unsigned(7,8) ,
45310	 => std_logic_vector(to_unsigned(62,8) ,
45311	 => std_logic_vector(to_unsigned(108,8) ,
45312	 => std_logic_vector(to_unsigned(82,8) ,
45313	 => std_logic_vector(to_unsigned(71,8) ,
45314	 => std_logic_vector(to_unsigned(91,8) ,
45315	 => std_logic_vector(to_unsigned(97,8) ,
45316	 => std_logic_vector(to_unsigned(97,8) ,
45317	 => std_logic_vector(to_unsigned(115,8) ,
45318	 => std_logic_vector(to_unsigned(101,8) ,
45319	 => std_logic_vector(to_unsigned(91,8) ,
45320	 => std_logic_vector(to_unsigned(103,8) ,
45321	 => std_logic_vector(to_unsigned(125,8) ,
45322	 => std_logic_vector(to_unsigned(108,8) ,
45323	 => std_logic_vector(to_unsigned(68,8) ,
45324	 => std_logic_vector(to_unsigned(69,8) ,
45325	 => std_logic_vector(to_unsigned(62,8) ,
45326	 => std_logic_vector(to_unsigned(16,8) ,
45327	 => std_logic_vector(to_unsigned(15,8) ,
45328	 => std_logic_vector(to_unsigned(28,8) ,
45329	 => std_logic_vector(to_unsigned(46,8) ,
45330	 => std_logic_vector(to_unsigned(49,8) ,
45331	 => std_logic_vector(to_unsigned(11,8) ,
45332	 => std_logic_vector(to_unsigned(2,8) ,
45333	 => std_logic_vector(to_unsigned(8,8) ,
45334	 => std_logic_vector(to_unsigned(17,8) ,
45335	 => std_logic_vector(to_unsigned(12,8) ,
45336	 => std_logic_vector(to_unsigned(6,8) ,
45337	 => std_logic_vector(to_unsigned(2,8) ,
45338	 => std_logic_vector(to_unsigned(9,8) ,
45339	 => std_logic_vector(to_unsigned(96,8) ,
45340	 => std_logic_vector(to_unsigned(99,8) ,
45341	 => std_logic_vector(to_unsigned(88,8) ,
45342	 => std_logic_vector(to_unsigned(95,8) ,
45343	 => std_logic_vector(to_unsigned(87,8) ,
45344	 => std_logic_vector(to_unsigned(84,8) ,
45345	 => std_logic_vector(to_unsigned(79,8) ,
45346	 => std_logic_vector(to_unsigned(91,8) ,
45347	 => std_logic_vector(to_unsigned(93,8) ,
45348	 => std_logic_vector(to_unsigned(81,8) ,
45349	 => std_logic_vector(to_unsigned(93,8) ,
45350	 => std_logic_vector(to_unsigned(80,8) ,
45351	 => std_logic_vector(to_unsigned(8,8) ,
45352	 => std_logic_vector(to_unsigned(3,8) ,
45353	 => std_logic_vector(to_unsigned(5,8) ,
45354	 => std_logic_vector(to_unsigned(11,8) ,
45355	 => std_logic_vector(to_unsigned(8,8) ,
45356	 => std_logic_vector(to_unsigned(5,8) ,
45357	 => std_logic_vector(to_unsigned(8,8) ,
45358	 => std_logic_vector(to_unsigned(3,8) ,
45359	 => std_logic_vector(to_unsigned(2,8) ,
45360	 => std_logic_vector(to_unsigned(5,8) ,
45361	 => std_logic_vector(to_unsigned(8,8) ,
45362	 => std_logic_vector(to_unsigned(7,8) ,
45363	 => std_logic_vector(to_unsigned(1,8) ,
45364	 => std_logic_vector(to_unsigned(7,8) ,
45365	 => std_logic_vector(to_unsigned(34,8) ,
45366	 => std_logic_vector(to_unsigned(29,8) ,
45367	 => std_logic_vector(to_unsigned(16,8) ,
45368	 => std_logic_vector(to_unsigned(7,8) ,
45369	 => std_logic_vector(to_unsigned(5,8) ,
45370	 => std_logic_vector(to_unsigned(9,8) ,
45371	 => std_logic_vector(to_unsigned(8,8) ,
45372	 => std_logic_vector(to_unsigned(3,8) ,
45373	 => std_logic_vector(to_unsigned(3,8) ,
45374	 => std_logic_vector(to_unsigned(1,8) ,
45375	 => std_logic_vector(to_unsigned(0,8) ,
45376	 => std_logic_vector(to_unsigned(0,8) ,
45377	 => std_logic_vector(to_unsigned(2,8) ,
45378	 => std_logic_vector(to_unsigned(2,8) ,
45379	 => std_logic_vector(to_unsigned(1,8) ,
45380	 => std_logic_vector(to_unsigned(1,8) ,
45381	 => std_logic_vector(to_unsigned(0,8) ,
45382	 => std_logic_vector(to_unsigned(0,8) ,
45383	 => std_logic_vector(to_unsigned(0,8) ,
45384	 => std_logic_vector(to_unsigned(0,8) ,
45385	 => std_logic_vector(to_unsigned(0,8) ,
45386	 => std_logic_vector(to_unsigned(1,8) ,
45387	 => std_logic_vector(to_unsigned(9,8) ,
45388	 => std_logic_vector(to_unsigned(10,8) ,
45389	 => std_logic_vector(to_unsigned(4,8) ,
45390	 => std_logic_vector(to_unsigned(4,8) ,
45391	 => std_logic_vector(to_unsigned(3,8) ,
45392	 => std_logic_vector(to_unsigned(7,8) ,
45393	 => std_logic_vector(to_unsigned(8,8) ,
45394	 => std_logic_vector(to_unsigned(3,8) ,
45395	 => std_logic_vector(to_unsigned(7,8) ,
45396	 => std_logic_vector(to_unsigned(15,8) ,
45397	 => std_logic_vector(to_unsigned(7,8) ,
45398	 => std_logic_vector(to_unsigned(0,8) ,
45399	 => std_logic_vector(to_unsigned(1,8) ,
45400	 => std_logic_vector(to_unsigned(1,8) ,
45401	 => std_logic_vector(to_unsigned(0,8) ,
45402	 => std_logic_vector(to_unsigned(2,8) ,
45403	 => std_logic_vector(to_unsigned(3,8) ,
45404	 => std_logic_vector(to_unsigned(3,8) ,
45405	 => std_logic_vector(to_unsigned(6,8) ,
45406	 => std_logic_vector(to_unsigned(7,8) ,
45407	 => std_logic_vector(to_unsigned(10,8) ,
45408	 => std_logic_vector(to_unsigned(14,8) ,
45409	 => std_logic_vector(to_unsigned(2,8) ,
45410	 => std_logic_vector(to_unsigned(1,8) ,
45411	 => std_logic_vector(to_unsigned(1,8) ,
45412	 => std_logic_vector(to_unsigned(1,8) ,
45413	 => std_logic_vector(to_unsigned(1,8) ,
45414	 => std_logic_vector(to_unsigned(2,8) ,
45415	 => std_logic_vector(to_unsigned(2,8) ,
45416	 => std_logic_vector(to_unsigned(1,8) ,
45417	 => std_logic_vector(to_unsigned(2,8) ,
45418	 => std_logic_vector(to_unsigned(1,8) ,
45419	 => std_logic_vector(to_unsigned(2,8) ,
45420	 => std_logic_vector(to_unsigned(2,8) ,
45421	 => std_logic_vector(to_unsigned(1,8) ,
45422	 => std_logic_vector(to_unsigned(2,8) ,
45423	 => std_logic_vector(to_unsigned(3,8) ,
45424	 => std_logic_vector(to_unsigned(2,8) ,
45425	 => std_logic_vector(to_unsigned(2,8) ,
45426	 => std_logic_vector(to_unsigned(2,8) ,
45427	 => std_logic_vector(to_unsigned(2,8) ,
45428	 => std_logic_vector(to_unsigned(2,8) ,
45429	 => std_logic_vector(to_unsigned(3,8) ,
45430	 => std_logic_vector(to_unsigned(2,8) ,
45431	 => std_logic_vector(to_unsigned(2,8) ,
45432	 => std_logic_vector(to_unsigned(2,8) ,
45433	 => std_logic_vector(to_unsigned(3,8) ,
45434	 => std_logic_vector(to_unsigned(3,8) ,
45435	 => std_logic_vector(to_unsigned(3,8) ,
45436	 => std_logic_vector(to_unsigned(3,8) ,
45437	 => std_logic_vector(to_unsigned(4,8) ,
45438	 => std_logic_vector(to_unsigned(3,8) ,
45439	 => std_logic_vector(to_unsigned(2,8) ,
45440	 => std_logic_vector(to_unsigned(3,8) ,
45441	 => std_logic_vector(to_unsigned(58,8) ,
45442	 => std_logic_vector(to_unsigned(51,8) ,
45443	 => std_logic_vector(to_unsigned(64,8) ,
45444	 => std_logic_vector(to_unsigned(62,8) ,
45445	 => std_logic_vector(to_unsigned(62,8) ,
45446	 => std_logic_vector(to_unsigned(66,8) ,
45447	 => std_logic_vector(to_unsigned(59,8) ,
45448	 => std_logic_vector(to_unsigned(51,8) ,
45449	 => std_logic_vector(to_unsigned(27,8) ,
45450	 => std_logic_vector(to_unsigned(34,8) ,
45451	 => std_logic_vector(to_unsigned(34,8) ,
45452	 => std_logic_vector(to_unsigned(35,8) ,
45453	 => std_logic_vector(to_unsigned(41,8) ,
45454	 => std_logic_vector(to_unsigned(46,8) ,
45455	 => std_logic_vector(to_unsigned(103,8) ,
45456	 => std_logic_vector(to_unsigned(122,8) ,
45457	 => std_logic_vector(to_unsigned(119,8) ,
45458	 => std_logic_vector(to_unsigned(111,8) ,
45459	 => std_logic_vector(to_unsigned(109,8) ,
45460	 => std_logic_vector(to_unsigned(105,8) ,
45461	 => std_logic_vector(to_unsigned(105,8) ,
45462	 => std_logic_vector(to_unsigned(115,8) ,
45463	 => std_logic_vector(to_unsigned(116,8) ,
45464	 => std_logic_vector(to_unsigned(127,8) ,
45465	 => std_logic_vector(to_unsigned(131,8) ,
45466	 => std_logic_vector(to_unsigned(146,8) ,
45467	 => std_logic_vector(to_unsigned(147,8) ,
45468	 => std_logic_vector(to_unsigned(144,8) ,
45469	 => std_logic_vector(to_unsigned(146,8) ,
45470	 => std_logic_vector(to_unsigned(146,8) ,
45471	 => std_logic_vector(to_unsigned(146,8) ,
45472	 => std_logic_vector(to_unsigned(146,8) ,
45473	 => std_logic_vector(to_unsigned(152,8) ,
45474	 => std_logic_vector(to_unsigned(154,8) ,
45475	 => std_logic_vector(to_unsigned(146,8) ,
45476	 => std_logic_vector(to_unsigned(149,8) ,
45477	 => std_logic_vector(to_unsigned(157,8) ,
45478	 => std_logic_vector(to_unsigned(152,8) ,
45479	 => std_logic_vector(to_unsigned(154,8) ,
45480	 => std_logic_vector(to_unsigned(156,8) ,
45481	 => std_logic_vector(to_unsigned(95,8) ,
45482	 => std_logic_vector(to_unsigned(52,8) ,
45483	 => std_logic_vector(to_unsigned(72,8) ,
45484	 => std_logic_vector(to_unsigned(74,8) ,
45485	 => std_logic_vector(to_unsigned(60,8) ,
45486	 => std_logic_vector(to_unsigned(71,8) ,
45487	 => std_logic_vector(to_unsigned(67,8) ,
45488	 => std_logic_vector(to_unsigned(73,8) ,
45489	 => std_logic_vector(to_unsigned(80,8) ,
45490	 => std_logic_vector(to_unsigned(78,8) ,
45491	 => std_logic_vector(to_unsigned(70,8) ,
45492	 => std_logic_vector(to_unsigned(86,8) ,
45493	 => std_logic_vector(to_unsigned(131,8) ,
45494	 => std_logic_vector(to_unsigned(146,8) ,
45495	 => std_logic_vector(to_unsigned(109,8) ,
45496	 => std_logic_vector(to_unsigned(101,8) ,
45497	 => std_logic_vector(to_unsigned(125,8) ,
45498	 => std_logic_vector(to_unsigned(138,8) ,
45499	 => std_logic_vector(to_unsigned(115,8) ,
45500	 => std_logic_vector(to_unsigned(118,8) ,
45501	 => std_logic_vector(to_unsigned(114,8) ,
45502	 => std_logic_vector(to_unsigned(84,8) ,
45503	 => std_logic_vector(to_unsigned(85,8) ,
45504	 => std_logic_vector(to_unsigned(91,8) ,
45505	 => std_logic_vector(to_unsigned(80,8) ,
45506	 => std_logic_vector(to_unsigned(78,8) ,
45507	 => std_logic_vector(to_unsigned(73,8) ,
45508	 => std_logic_vector(to_unsigned(73,8) ,
45509	 => std_logic_vector(to_unsigned(77,8) ,
45510	 => std_logic_vector(to_unsigned(76,8) ,
45511	 => std_logic_vector(to_unsigned(68,8) ,
45512	 => std_logic_vector(to_unsigned(63,8) ,
45513	 => std_logic_vector(to_unsigned(60,8) ,
45514	 => std_logic_vector(to_unsigned(59,8) ,
45515	 => std_logic_vector(to_unsigned(72,8) ,
45516	 => std_logic_vector(to_unsigned(92,8) ,
45517	 => std_logic_vector(to_unsigned(100,8) ,
45518	 => std_logic_vector(to_unsigned(105,8) ,
45519	 => std_logic_vector(to_unsigned(109,8) ,
45520	 => std_logic_vector(to_unsigned(93,8) ,
45521	 => std_logic_vector(to_unsigned(77,8) ,
45522	 => std_logic_vector(to_unsigned(77,8) ,
45523	 => std_logic_vector(to_unsigned(81,8) ,
45524	 => std_logic_vector(to_unsigned(92,8) ,
45525	 => std_logic_vector(to_unsigned(91,8) ,
45526	 => std_logic_vector(to_unsigned(84,8) ,
45527	 => std_logic_vector(to_unsigned(58,8) ,
45528	 => std_logic_vector(to_unsigned(62,8) ,
45529	 => std_logic_vector(to_unsigned(56,8) ,
45530	 => std_logic_vector(to_unsigned(48,8) ,
45531	 => std_logic_vector(to_unsigned(57,8) ,
45532	 => std_logic_vector(to_unsigned(72,8) ,
45533	 => std_logic_vector(to_unsigned(74,8) ,
45534	 => std_logic_vector(to_unsigned(64,8) ,
45535	 => std_logic_vector(to_unsigned(59,8) ,
45536	 => std_logic_vector(to_unsigned(69,8) ,
45537	 => std_logic_vector(to_unsigned(79,8) ,
45538	 => std_logic_vector(to_unsigned(78,8) ,
45539	 => std_logic_vector(to_unsigned(90,8) ,
45540	 => std_logic_vector(to_unsigned(76,8) ,
45541	 => std_logic_vector(to_unsigned(73,8) ,
45542	 => std_logic_vector(to_unsigned(71,8) ,
45543	 => std_logic_vector(to_unsigned(60,8) ,
45544	 => std_logic_vector(to_unsigned(84,8) ,
45545	 => std_logic_vector(to_unsigned(71,8) ,
45546	 => std_logic_vector(to_unsigned(69,8) ,
45547	 => std_logic_vector(to_unsigned(97,8) ,
45548	 => std_logic_vector(to_unsigned(87,8) ,
45549	 => std_logic_vector(to_unsigned(90,8) ,
45550	 => std_logic_vector(to_unsigned(88,8) ,
45551	 => std_logic_vector(to_unsigned(91,8) ,
45552	 => std_logic_vector(to_unsigned(90,8) ,
45553	 => std_logic_vector(to_unsigned(72,8) ,
45554	 => std_logic_vector(to_unsigned(77,8) ,
45555	 => std_logic_vector(to_unsigned(65,8) ,
45556	 => std_logic_vector(to_unsigned(66,8) ,
45557	 => std_logic_vector(to_unsigned(69,8) ,
45558	 => std_logic_vector(to_unsigned(64,8) ,
45559	 => std_logic_vector(to_unsigned(69,8) ,
45560	 => std_logic_vector(to_unsigned(74,8) ,
45561	 => std_logic_vector(to_unsigned(72,8) ,
45562	 => std_logic_vector(to_unsigned(68,8) ,
45563	 => std_logic_vector(to_unsigned(11,8) ,
45564	 => std_logic_vector(to_unsigned(5,8) ,
45565	 => std_logic_vector(to_unsigned(8,8) ,
45566	 => std_logic_vector(to_unsigned(4,8) ,
45567	 => std_logic_vector(to_unsigned(4,8) ,
45568	 => std_logic_vector(to_unsigned(7,8) ,
45569	 => std_logic_vector(to_unsigned(90,8) ,
45570	 => std_logic_vector(to_unsigned(122,8) ,
45571	 => std_logic_vector(to_unsigned(86,8) ,
45572	 => std_logic_vector(to_unsigned(130,8) ,
45573	 => std_logic_vector(to_unsigned(124,8) ,
45574	 => std_logic_vector(to_unsigned(121,8) ,
45575	 => std_logic_vector(to_unsigned(118,8) ,
45576	 => std_logic_vector(to_unsigned(86,8) ,
45577	 => std_logic_vector(to_unsigned(60,8) ,
45578	 => std_logic_vector(to_unsigned(71,8) ,
45579	 => std_logic_vector(to_unsigned(73,8) ,
45580	 => std_logic_vector(to_unsigned(71,8) ,
45581	 => std_logic_vector(to_unsigned(54,8) ,
45582	 => std_logic_vector(to_unsigned(54,8) ,
45583	 => std_logic_vector(to_unsigned(61,8) ,
45584	 => std_logic_vector(to_unsigned(69,8) ,
45585	 => std_logic_vector(to_unsigned(51,8) ,
45586	 => std_logic_vector(to_unsigned(49,8) ,
45587	 => std_logic_vector(to_unsigned(48,8) ,
45588	 => std_logic_vector(to_unsigned(54,8) ,
45589	 => std_logic_vector(to_unsigned(60,8) ,
45590	 => std_logic_vector(to_unsigned(51,8) ,
45591	 => std_logic_vector(to_unsigned(54,8) ,
45592	 => std_logic_vector(to_unsigned(49,8) ,
45593	 => std_logic_vector(to_unsigned(45,8) ,
45594	 => std_logic_vector(to_unsigned(24,8) ,
45595	 => std_logic_vector(to_unsigned(20,8) ,
45596	 => std_logic_vector(to_unsigned(36,8) ,
45597	 => std_logic_vector(to_unsigned(86,8) ,
45598	 => std_logic_vector(to_unsigned(77,8) ,
45599	 => std_logic_vector(to_unsigned(73,8) ,
45600	 => std_logic_vector(to_unsigned(81,8) ,
45601	 => std_logic_vector(to_unsigned(77,8) ,
45602	 => std_logic_vector(to_unsigned(53,8) ,
45603	 => std_logic_vector(to_unsigned(58,8) ,
45604	 => std_logic_vector(to_unsigned(35,8) ,
45605	 => std_logic_vector(to_unsigned(20,8) ,
45606	 => std_logic_vector(to_unsigned(32,8) ,
45607	 => std_logic_vector(to_unsigned(35,8) ,
45608	 => std_logic_vector(to_unsigned(59,8) ,
45609	 => std_logic_vector(to_unsigned(70,8) ,
45610	 => std_logic_vector(to_unsigned(80,8) ,
45611	 => std_logic_vector(to_unsigned(74,8) ,
45612	 => std_logic_vector(to_unsigned(26,8) ,
45613	 => std_logic_vector(to_unsigned(27,8) ,
45614	 => std_logic_vector(to_unsigned(53,8) ,
45615	 => std_logic_vector(to_unsigned(45,8) ,
45616	 => std_logic_vector(to_unsigned(39,8) ,
45617	 => std_logic_vector(to_unsigned(40,8) ,
45618	 => std_logic_vector(to_unsigned(45,8) ,
45619	 => std_logic_vector(to_unsigned(43,8) ,
45620	 => std_logic_vector(to_unsigned(58,8) ,
45621	 => std_logic_vector(to_unsigned(51,8) ,
45622	 => std_logic_vector(to_unsigned(57,8) ,
45623	 => std_logic_vector(to_unsigned(57,8) ,
45624	 => std_logic_vector(to_unsigned(4,8) ,
45625	 => std_logic_vector(to_unsigned(3,8) ,
45626	 => std_logic_vector(to_unsigned(4,8) ,
45627	 => std_logic_vector(to_unsigned(2,8) ,
45628	 => std_logic_vector(to_unsigned(8,8) ,
45629	 => std_logic_vector(to_unsigned(26,8) ,
45630	 => std_logic_vector(to_unsigned(60,8) ,
45631	 => std_logic_vector(to_unsigned(95,8) ,
45632	 => std_logic_vector(to_unsigned(69,8) ,
45633	 => std_logic_vector(to_unsigned(61,8) ,
45634	 => std_logic_vector(to_unsigned(73,8) ,
45635	 => std_logic_vector(to_unsigned(71,8) ,
45636	 => std_logic_vector(to_unsigned(66,8) ,
45637	 => std_logic_vector(to_unsigned(82,8) ,
45638	 => std_logic_vector(to_unsigned(76,8) ,
45639	 => std_logic_vector(to_unsigned(55,8) ,
45640	 => std_logic_vector(to_unsigned(70,8) ,
45641	 => std_logic_vector(to_unsigned(112,8) ,
45642	 => std_logic_vector(to_unsigned(121,8) ,
45643	 => std_logic_vector(to_unsigned(85,8) ,
45644	 => std_logic_vector(to_unsigned(87,8) ,
45645	 => std_logic_vector(to_unsigned(63,8) ,
45646	 => std_logic_vector(to_unsigned(14,8) ,
45647	 => std_logic_vector(to_unsigned(22,8) ,
45648	 => std_logic_vector(to_unsigned(29,8) ,
45649	 => std_logic_vector(to_unsigned(26,8) ,
45650	 => std_logic_vector(to_unsigned(28,8) ,
45651	 => std_logic_vector(to_unsigned(4,8) ,
45652	 => std_logic_vector(to_unsigned(3,8) ,
45653	 => std_logic_vector(to_unsigned(8,8) ,
45654	 => std_logic_vector(to_unsigned(12,8) ,
45655	 => std_logic_vector(to_unsigned(12,8) ,
45656	 => std_logic_vector(to_unsigned(9,8) ,
45657	 => std_logic_vector(to_unsigned(2,8) ,
45658	 => std_logic_vector(to_unsigned(8,8) ,
45659	 => std_logic_vector(to_unsigned(85,8) ,
45660	 => std_logic_vector(to_unsigned(97,8) ,
45661	 => std_logic_vector(to_unsigned(90,8) ,
45662	 => std_logic_vector(to_unsigned(100,8) ,
45663	 => std_logic_vector(to_unsigned(101,8) ,
45664	 => std_logic_vector(to_unsigned(97,8) ,
45665	 => std_logic_vector(to_unsigned(97,8) ,
45666	 => std_logic_vector(to_unsigned(101,8) ,
45667	 => std_logic_vector(to_unsigned(101,8) ,
45668	 => std_logic_vector(to_unsigned(90,8) ,
45669	 => std_logic_vector(to_unsigned(97,8) ,
45670	 => std_logic_vector(to_unsigned(72,8) ,
45671	 => std_logic_vector(to_unsigned(5,8) ,
45672	 => std_logic_vector(to_unsigned(7,8) ,
45673	 => std_logic_vector(to_unsigned(19,8) ,
45674	 => std_logic_vector(to_unsigned(11,8) ,
45675	 => std_logic_vector(to_unsigned(6,8) ,
45676	 => std_logic_vector(to_unsigned(3,8) ,
45677	 => std_logic_vector(to_unsigned(2,8) ,
45678	 => std_logic_vector(to_unsigned(4,8) ,
45679	 => std_logic_vector(to_unsigned(6,8) ,
45680	 => std_logic_vector(to_unsigned(4,8) ,
45681	 => std_logic_vector(to_unsigned(5,8) ,
45682	 => std_logic_vector(to_unsigned(3,8) ,
45683	 => std_logic_vector(to_unsigned(1,8) ,
45684	 => std_logic_vector(to_unsigned(60,8) ,
45685	 => std_logic_vector(to_unsigned(136,8) ,
45686	 => std_logic_vector(to_unsigned(130,8) ,
45687	 => std_logic_vector(to_unsigned(59,8) ,
45688	 => std_logic_vector(to_unsigned(4,8) ,
45689	 => std_logic_vector(to_unsigned(8,8) ,
45690	 => std_logic_vector(to_unsigned(97,8) ,
45691	 => std_logic_vector(to_unsigned(103,8) ,
45692	 => std_logic_vector(to_unsigned(54,8) ,
45693	 => std_logic_vector(to_unsigned(80,8) ,
45694	 => std_logic_vector(to_unsigned(33,8) ,
45695	 => std_logic_vector(to_unsigned(34,8) ,
45696	 => std_logic_vector(to_unsigned(16,8) ,
45697	 => std_logic_vector(to_unsigned(2,8) ,
45698	 => std_logic_vector(to_unsigned(2,8) ,
45699	 => std_logic_vector(to_unsigned(1,8) ,
45700	 => std_logic_vector(to_unsigned(2,8) ,
45701	 => std_logic_vector(to_unsigned(1,8) ,
45702	 => std_logic_vector(to_unsigned(0,8) ,
45703	 => std_logic_vector(to_unsigned(0,8) ,
45704	 => std_logic_vector(to_unsigned(0,8) ,
45705	 => std_logic_vector(to_unsigned(0,8) ,
45706	 => std_logic_vector(to_unsigned(0,8) ,
45707	 => std_logic_vector(to_unsigned(1,8) ,
45708	 => std_logic_vector(to_unsigned(1,8) ,
45709	 => std_logic_vector(to_unsigned(1,8) ,
45710	 => std_logic_vector(to_unsigned(0,8) ,
45711	 => std_logic_vector(to_unsigned(2,8) ,
45712	 => std_logic_vector(to_unsigned(6,8) ,
45713	 => std_logic_vector(to_unsigned(6,8) ,
45714	 => std_logic_vector(to_unsigned(2,8) ,
45715	 => std_logic_vector(to_unsigned(4,8) ,
45716	 => std_logic_vector(to_unsigned(10,8) ,
45717	 => std_logic_vector(to_unsigned(7,8) ,
45718	 => std_logic_vector(to_unsigned(0,8) ,
45719	 => std_logic_vector(to_unsigned(1,8) ,
45720	 => std_logic_vector(to_unsigned(1,8) ,
45721	 => std_logic_vector(to_unsigned(0,8) ,
45722	 => std_logic_vector(to_unsigned(2,8) ,
45723	 => std_logic_vector(to_unsigned(3,8) ,
45724	 => std_logic_vector(to_unsigned(4,8) ,
45725	 => std_logic_vector(to_unsigned(4,8) ,
45726	 => std_logic_vector(to_unsigned(5,8) ,
45727	 => std_logic_vector(to_unsigned(9,8) ,
45728	 => std_logic_vector(to_unsigned(14,8) ,
45729	 => std_logic_vector(to_unsigned(3,8) ,
45730	 => std_logic_vector(to_unsigned(1,8) ,
45731	 => std_logic_vector(to_unsigned(2,8) ,
45732	 => std_logic_vector(to_unsigned(1,8) ,
45733	 => std_logic_vector(to_unsigned(2,8) ,
45734	 => std_logic_vector(to_unsigned(2,8) ,
45735	 => std_logic_vector(to_unsigned(2,8) ,
45736	 => std_logic_vector(to_unsigned(2,8) ,
45737	 => std_logic_vector(to_unsigned(2,8) ,
45738	 => std_logic_vector(to_unsigned(2,8) ,
45739	 => std_logic_vector(to_unsigned(3,8) ,
45740	 => std_logic_vector(to_unsigned(3,8) ,
45741	 => std_logic_vector(to_unsigned(2,8) ,
45742	 => std_logic_vector(to_unsigned(2,8) ,
45743	 => std_logic_vector(to_unsigned(2,8) ,
45744	 => std_logic_vector(to_unsigned(2,8) ,
45745	 => std_logic_vector(to_unsigned(1,8) ,
45746	 => std_logic_vector(to_unsigned(2,8) ,
45747	 => std_logic_vector(to_unsigned(3,8) ,
45748	 => std_logic_vector(to_unsigned(2,8) ,
45749	 => std_logic_vector(to_unsigned(2,8) ,
45750	 => std_logic_vector(to_unsigned(2,8) ,
45751	 => std_logic_vector(to_unsigned(2,8) ,
45752	 => std_logic_vector(to_unsigned(3,8) ,
45753	 => std_logic_vector(to_unsigned(2,8) ,
45754	 => std_logic_vector(to_unsigned(3,8) ,
45755	 => std_logic_vector(to_unsigned(4,8) ,
45756	 => std_logic_vector(to_unsigned(3,8) ,
45757	 => std_logic_vector(to_unsigned(3,8) ,
45758	 => std_logic_vector(to_unsigned(2,8) ,
45759	 => std_logic_vector(to_unsigned(2,8) ,
45760	 => std_logic_vector(to_unsigned(2,8) ,
45761	 => std_logic_vector(to_unsigned(72,8) ,
45762	 => std_logic_vector(to_unsigned(66,8) ,
45763	 => std_logic_vector(to_unsigned(56,8) ,
45764	 => std_logic_vector(to_unsigned(55,8) ,
45765	 => std_logic_vector(to_unsigned(51,8) ,
45766	 => std_logic_vector(to_unsigned(66,8) ,
45767	 => std_logic_vector(to_unsigned(62,8) ,
45768	 => std_logic_vector(to_unsigned(45,8) ,
45769	 => std_logic_vector(to_unsigned(32,8) ,
45770	 => std_logic_vector(to_unsigned(34,8) ,
45771	 => std_logic_vector(to_unsigned(30,8) ,
45772	 => std_logic_vector(to_unsigned(34,8) ,
45773	 => std_logic_vector(to_unsigned(36,8) ,
45774	 => std_logic_vector(to_unsigned(51,8) ,
45775	 => std_logic_vector(to_unsigned(103,8) ,
45776	 => std_logic_vector(to_unsigned(111,8) ,
45777	 => std_logic_vector(to_unsigned(114,8) ,
45778	 => std_logic_vector(to_unsigned(115,8) ,
45779	 => std_logic_vector(to_unsigned(108,8) ,
45780	 => std_logic_vector(to_unsigned(114,8) ,
45781	 => std_logic_vector(to_unsigned(112,8) ,
45782	 => std_logic_vector(to_unsigned(115,8) ,
45783	 => std_logic_vector(to_unsigned(115,8) ,
45784	 => std_logic_vector(to_unsigned(124,8) ,
45785	 => std_logic_vector(to_unsigned(128,8) ,
45786	 => std_logic_vector(to_unsigned(138,8) ,
45787	 => std_logic_vector(to_unsigned(146,8) ,
45788	 => std_logic_vector(to_unsigned(136,8) ,
45789	 => std_logic_vector(to_unsigned(139,8) ,
45790	 => std_logic_vector(to_unsigned(144,8) ,
45791	 => std_logic_vector(to_unsigned(138,8) ,
45792	 => std_logic_vector(to_unsigned(138,8) ,
45793	 => std_logic_vector(to_unsigned(154,8) ,
45794	 => std_logic_vector(to_unsigned(151,8) ,
45795	 => std_logic_vector(to_unsigned(144,8) ,
45796	 => std_logic_vector(to_unsigned(152,8) ,
45797	 => std_logic_vector(to_unsigned(159,8) ,
45798	 => std_logic_vector(to_unsigned(152,8) ,
45799	 => std_logic_vector(to_unsigned(151,8) ,
45800	 => std_logic_vector(to_unsigned(156,8) ,
45801	 => std_logic_vector(to_unsigned(116,8) ,
45802	 => std_logic_vector(to_unsigned(85,8) ,
45803	 => std_logic_vector(to_unsigned(77,8) ,
45804	 => std_logic_vector(to_unsigned(73,8) ,
45805	 => std_logic_vector(to_unsigned(65,8) ,
45806	 => std_logic_vector(to_unsigned(64,8) ,
45807	 => std_logic_vector(to_unsigned(63,8) ,
45808	 => std_logic_vector(to_unsigned(70,8) ,
45809	 => std_logic_vector(to_unsigned(72,8) ,
45810	 => std_logic_vector(to_unsigned(77,8) ,
45811	 => std_logic_vector(to_unsigned(69,8) ,
45812	 => std_logic_vector(to_unsigned(73,8) ,
45813	 => std_logic_vector(to_unsigned(70,8) ,
45814	 => std_logic_vector(to_unsigned(81,8) ,
45815	 => std_logic_vector(to_unsigned(101,8) ,
45816	 => std_logic_vector(to_unsigned(109,8) ,
45817	 => std_logic_vector(to_unsigned(122,8) ,
45818	 => std_logic_vector(to_unsigned(116,8) ,
45819	 => std_logic_vector(to_unsigned(97,8) ,
45820	 => std_logic_vector(to_unsigned(93,8) ,
45821	 => std_logic_vector(to_unsigned(97,8) ,
45822	 => std_logic_vector(to_unsigned(78,8) ,
45823	 => std_logic_vector(to_unsigned(82,8) ,
45824	 => std_logic_vector(to_unsigned(86,8) ,
45825	 => std_logic_vector(to_unsigned(77,8) ,
45826	 => std_logic_vector(to_unsigned(71,8) ,
45827	 => std_logic_vector(to_unsigned(71,8) ,
45828	 => std_logic_vector(to_unsigned(74,8) ,
45829	 => std_logic_vector(to_unsigned(80,8) ,
45830	 => std_logic_vector(to_unsigned(73,8) ,
45831	 => std_logic_vector(to_unsigned(62,8) ,
45832	 => std_logic_vector(to_unsigned(59,8) ,
45833	 => std_logic_vector(to_unsigned(62,8) ,
45834	 => std_logic_vector(to_unsigned(55,8) ,
45835	 => std_logic_vector(to_unsigned(63,8) ,
45836	 => std_logic_vector(to_unsigned(93,8) ,
45837	 => std_logic_vector(to_unsigned(101,8) ,
45838	 => std_logic_vector(to_unsigned(91,8) ,
45839	 => std_logic_vector(to_unsigned(100,8) ,
45840	 => std_logic_vector(to_unsigned(79,8) ,
45841	 => std_logic_vector(to_unsigned(66,8) ,
45842	 => std_logic_vector(to_unsigned(82,8) ,
45843	 => std_logic_vector(to_unsigned(87,8) ,
45844	 => std_logic_vector(to_unsigned(74,8) ,
45845	 => std_logic_vector(to_unsigned(69,8) ,
45846	 => std_logic_vector(to_unsigned(68,8) ,
45847	 => std_logic_vector(to_unsigned(50,8) ,
45848	 => std_logic_vector(to_unsigned(59,8) ,
45849	 => std_logic_vector(to_unsigned(54,8) ,
45850	 => std_logic_vector(to_unsigned(45,8) ,
45851	 => std_logic_vector(to_unsigned(49,8) ,
45852	 => std_logic_vector(to_unsigned(57,8) ,
45853	 => std_logic_vector(to_unsigned(61,8) ,
45854	 => std_logic_vector(to_unsigned(60,8) ,
45855	 => std_logic_vector(to_unsigned(59,8) ,
45856	 => std_logic_vector(to_unsigned(77,8) ,
45857	 => std_logic_vector(to_unsigned(88,8) ,
45858	 => std_logic_vector(to_unsigned(71,8) ,
45859	 => std_logic_vector(to_unsigned(92,8) ,
45860	 => std_logic_vector(to_unsigned(96,8) ,
45861	 => std_logic_vector(to_unsigned(86,8) ,
45862	 => std_logic_vector(to_unsigned(78,8) ,
45863	 => std_logic_vector(to_unsigned(91,8) ,
45864	 => std_logic_vector(to_unsigned(92,8) ,
45865	 => std_logic_vector(to_unsigned(77,8) ,
45866	 => std_logic_vector(to_unsigned(84,8) ,
45867	 => std_logic_vector(to_unsigned(95,8) ,
45868	 => std_logic_vector(to_unsigned(82,8) ,
45869	 => std_logic_vector(to_unsigned(86,8) ,
45870	 => std_logic_vector(to_unsigned(82,8) ,
45871	 => std_logic_vector(to_unsigned(82,8) ,
45872	 => std_logic_vector(to_unsigned(92,8) ,
45873	 => std_logic_vector(to_unsigned(68,8) ,
45874	 => std_logic_vector(to_unsigned(69,8) ,
45875	 => std_logic_vector(to_unsigned(58,8) ,
45876	 => std_logic_vector(to_unsigned(45,8) ,
45877	 => std_logic_vector(to_unsigned(54,8) ,
45878	 => std_logic_vector(to_unsigned(61,8) ,
45879	 => std_logic_vector(to_unsigned(63,8) ,
45880	 => std_logic_vector(to_unsigned(71,8) ,
45881	 => std_logic_vector(to_unsigned(72,8) ,
45882	 => std_logic_vector(to_unsigned(81,8) ,
45883	 => std_logic_vector(to_unsigned(33,8) ,
45884	 => std_logic_vector(to_unsigned(11,8) ,
45885	 => std_logic_vector(to_unsigned(13,8) ,
45886	 => std_logic_vector(to_unsigned(11,8) ,
45887	 => std_logic_vector(to_unsigned(16,8) ,
45888	 => std_logic_vector(to_unsigned(78,8) ,
45889	 => std_logic_vector(to_unsigned(112,8) ,
45890	 => std_logic_vector(to_unsigned(87,8) ,
45891	 => std_logic_vector(to_unsigned(99,8) ,
45892	 => std_logic_vector(to_unsigned(103,8) ,
45893	 => std_logic_vector(to_unsigned(96,8) ,
45894	 => std_logic_vector(to_unsigned(97,8) ,
45895	 => std_logic_vector(to_unsigned(104,8) ,
45896	 => std_logic_vector(to_unsigned(73,8) ,
45897	 => std_logic_vector(to_unsigned(53,8) ,
45898	 => std_logic_vector(to_unsigned(60,8) ,
45899	 => std_logic_vector(to_unsigned(45,8) ,
45900	 => std_logic_vector(to_unsigned(57,8) ,
45901	 => std_logic_vector(to_unsigned(51,8) ,
45902	 => std_logic_vector(to_unsigned(49,8) ,
45903	 => std_logic_vector(to_unsigned(85,8) ,
45904	 => std_logic_vector(to_unsigned(70,8) ,
45905	 => std_logic_vector(to_unsigned(39,8) ,
45906	 => std_logic_vector(to_unsigned(46,8) ,
45907	 => std_logic_vector(to_unsigned(38,8) ,
45908	 => std_logic_vector(to_unsigned(32,8) ,
45909	 => std_logic_vector(to_unsigned(43,8) ,
45910	 => std_logic_vector(to_unsigned(54,8) ,
45911	 => std_logic_vector(to_unsigned(47,8) ,
45912	 => std_logic_vector(to_unsigned(33,8) ,
45913	 => std_logic_vector(to_unsigned(24,8) ,
45914	 => std_logic_vector(to_unsigned(18,8) ,
45915	 => std_logic_vector(to_unsigned(19,8) ,
45916	 => std_logic_vector(to_unsigned(23,8) ,
45917	 => std_logic_vector(to_unsigned(40,8) ,
45918	 => std_logic_vector(to_unsigned(49,8) ,
45919	 => std_logic_vector(to_unsigned(58,8) ,
45920	 => std_logic_vector(to_unsigned(59,8) ,
45921	 => std_logic_vector(to_unsigned(52,8) ,
45922	 => std_logic_vector(to_unsigned(39,8) ,
45923	 => std_logic_vector(to_unsigned(58,8) ,
45924	 => std_logic_vector(to_unsigned(54,8) ,
45925	 => std_logic_vector(to_unsigned(16,8) ,
45926	 => std_logic_vector(to_unsigned(18,8) ,
45927	 => std_logic_vector(to_unsigned(22,8) ,
45928	 => std_logic_vector(to_unsigned(27,8) ,
45929	 => std_logic_vector(to_unsigned(57,8) ,
45930	 => std_logic_vector(to_unsigned(70,8) ,
45931	 => std_logic_vector(to_unsigned(76,8) ,
45932	 => std_logic_vector(to_unsigned(40,8) ,
45933	 => std_logic_vector(to_unsigned(57,8) ,
45934	 => std_logic_vector(to_unsigned(66,8) ,
45935	 => std_logic_vector(to_unsigned(25,8) ,
45936	 => std_logic_vector(to_unsigned(19,8) ,
45937	 => std_logic_vector(to_unsigned(30,8) ,
45938	 => std_logic_vector(to_unsigned(29,8) ,
45939	 => std_logic_vector(to_unsigned(40,8) ,
45940	 => std_logic_vector(to_unsigned(35,8) ,
45941	 => std_logic_vector(to_unsigned(28,8) ,
45942	 => std_logic_vector(to_unsigned(48,8) ,
45943	 => std_logic_vector(to_unsigned(61,8) ,
45944	 => std_logic_vector(to_unsigned(28,8) ,
45945	 => std_logic_vector(to_unsigned(8,8) ,
45946	 => std_logic_vector(to_unsigned(6,8) ,
45947	 => std_logic_vector(to_unsigned(13,8) ,
45948	 => std_logic_vector(to_unsigned(23,8) ,
45949	 => std_logic_vector(to_unsigned(18,8) ,
45950	 => std_logic_vector(to_unsigned(41,8) ,
45951	 => std_logic_vector(to_unsigned(92,8) ,
45952	 => std_logic_vector(to_unsigned(82,8) ,
45953	 => std_logic_vector(to_unsigned(88,8) ,
45954	 => std_logic_vector(to_unsigned(90,8) ,
45955	 => std_logic_vector(to_unsigned(85,8) ,
45956	 => std_logic_vector(to_unsigned(79,8) ,
45957	 => std_logic_vector(to_unsigned(84,8) ,
45958	 => std_logic_vector(to_unsigned(84,8) ,
45959	 => std_logic_vector(to_unsigned(71,8) ,
45960	 => std_logic_vector(to_unsigned(70,8) ,
45961	 => std_logic_vector(to_unsigned(107,8) ,
45962	 => std_logic_vector(to_unsigned(109,8) ,
45963	 => std_logic_vector(to_unsigned(84,8) ,
45964	 => std_logic_vector(to_unsigned(93,8) ,
45965	 => std_logic_vector(to_unsigned(51,8) ,
45966	 => std_logic_vector(to_unsigned(6,8) ,
45967	 => std_logic_vector(to_unsigned(24,8) ,
45968	 => std_logic_vector(to_unsigned(30,8) ,
45969	 => std_logic_vector(to_unsigned(20,8) ,
45970	 => std_logic_vector(to_unsigned(8,8) ,
45971	 => std_logic_vector(to_unsigned(2,8) ,
45972	 => std_logic_vector(to_unsigned(9,8) ,
45973	 => std_logic_vector(to_unsigned(5,8) ,
45974	 => std_logic_vector(to_unsigned(9,8) ,
45975	 => std_logic_vector(to_unsigned(12,8) ,
45976	 => std_logic_vector(to_unsigned(6,8) ,
45977	 => std_logic_vector(to_unsigned(1,8) ,
45978	 => std_logic_vector(to_unsigned(8,8) ,
45979	 => std_logic_vector(to_unsigned(90,8) ,
45980	 => std_logic_vector(to_unsigned(87,8) ,
45981	 => std_logic_vector(to_unsigned(84,8) ,
45982	 => std_logic_vector(to_unsigned(100,8) ,
45983	 => std_logic_vector(to_unsigned(99,8) ,
45984	 => std_logic_vector(to_unsigned(104,8) ,
45985	 => std_logic_vector(to_unsigned(104,8) ,
45986	 => std_logic_vector(to_unsigned(92,8) ,
45987	 => std_logic_vector(to_unsigned(95,8) ,
45988	 => std_logic_vector(to_unsigned(101,8) ,
45989	 => std_logic_vector(to_unsigned(99,8) ,
45990	 => std_logic_vector(to_unsigned(71,8) ,
45991	 => std_logic_vector(to_unsigned(5,8) ,
45992	 => std_logic_vector(to_unsigned(6,8) ,
45993	 => std_logic_vector(to_unsigned(16,8) ,
45994	 => std_logic_vector(to_unsigned(10,8) ,
45995	 => std_logic_vector(to_unsigned(8,8) ,
45996	 => std_logic_vector(to_unsigned(2,8) ,
45997	 => std_logic_vector(to_unsigned(2,8) ,
45998	 => std_logic_vector(to_unsigned(6,8) ,
45999	 => std_logic_vector(to_unsigned(5,8) ,
46000	 => std_logic_vector(to_unsigned(2,8) ,
46001	 => std_logic_vector(to_unsigned(3,8) ,
46002	 => std_logic_vector(to_unsigned(1,8) ,
46003	 => std_logic_vector(to_unsigned(7,8) ,
46004	 => std_logic_vector(to_unsigned(111,8) ,
46005	 => std_logic_vector(to_unsigned(111,8) ,
46006	 => std_logic_vector(to_unsigned(107,8) ,
46007	 => std_logic_vector(to_unsigned(46,8) ,
46008	 => std_logic_vector(to_unsigned(4,8) ,
46009	 => std_logic_vector(to_unsigned(7,8) ,
46010	 => std_logic_vector(to_unsigned(91,8) ,
46011	 => std_logic_vector(to_unsigned(149,8) ,
46012	 => std_logic_vector(to_unsigned(130,8) ,
46013	 => std_logic_vector(to_unsigned(164,8) ,
46014	 => std_logic_vector(to_unsigned(118,8) ,
46015	 => std_logic_vector(to_unsigned(173,8) ,
46016	 => std_logic_vector(to_unsigned(99,8) ,
46017	 => std_logic_vector(to_unsigned(4,8) ,
46018	 => std_logic_vector(to_unsigned(2,8) ,
46019	 => std_logic_vector(to_unsigned(1,8) ,
46020	 => std_logic_vector(to_unsigned(2,8) ,
46021	 => std_logic_vector(to_unsigned(1,8) ,
46022	 => std_logic_vector(to_unsigned(0,8) ,
46023	 => std_logic_vector(to_unsigned(12,8) ,
46024	 => std_logic_vector(to_unsigned(48,8) ,
46025	 => std_logic_vector(to_unsigned(26,8) ,
46026	 => std_logic_vector(to_unsigned(13,8) ,
46027	 => std_logic_vector(to_unsigned(14,8) ,
46028	 => std_logic_vector(to_unsigned(9,8) ,
46029	 => std_logic_vector(to_unsigned(3,8) ,
46030	 => std_logic_vector(to_unsigned(1,8) ,
46031	 => std_logic_vector(to_unsigned(5,8) ,
46032	 => std_logic_vector(to_unsigned(9,8) ,
46033	 => std_logic_vector(to_unsigned(5,8) ,
46034	 => std_logic_vector(to_unsigned(1,8) ,
46035	 => std_logic_vector(to_unsigned(1,8) ,
46036	 => std_logic_vector(to_unsigned(6,8) ,
46037	 => std_logic_vector(to_unsigned(7,8) ,
46038	 => std_logic_vector(to_unsigned(1,8) ,
46039	 => std_logic_vector(to_unsigned(0,8) ,
46040	 => std_logic_vector(to_unsigned(0,8) ,
46041	 => std_logic_vector(to_unsigned(0,8) ,
46042	 => std_logic_vector(to_unsigned(2,8) ,
46043	 => std_logic_vector(to_unsigned(3,8) ,
46044	 => std_logic_vector(to_unsigned(3,8) ,
46045	 => std_logic_vector(to_unsigned(6,8) ,
46046	 => std_logic_vector(to_unsigned(6,8) ,
46047	 => std_logic_vector(to_unsigned(5,8) ,
46048	 => std_logic_vector(to_unsigned(8,8) ,
46049	 => std_logic_vector(to_unsigned(2,8) ,
46050	 => std_logic_vector(to_unsigned(1,8) ,
46051	 => std_logic_vector(to_unsigned(1,8) ,
46052	 => std_logic_vector(to_unsigned(2,8) ,
46053	 => std_logic_vector(to_unsigned(3,8) ,
46054	 => std_logic_vector(to_unsigned(3,8) ,
46055	 => std_logic_vector(to_unsigned(4,8) ,
46056	 => std_logic_vector(to_unsigned(3,8) ,
46057	 => std_logic_vector(to_unsigned(4,8) ,
46058	 => std_logic_vector(to_unsigned(4,8) ,
46059	 => std_logic_vector(to_unsigned(3,8) ,
46060	 => std_logic_vector(to_unsigned(3,8) ,
46061	 => std_logic_vector(to_unsigned(3,8) ,
46062	 => std_logic_vector(to_unsigned(2,8) ,
46063	 => std_logic_vector(to_unsigned(1,8) ,
46064	 => std_logic_vector(to_unsigned(1,8) ,
46065	 => std_logic_vector(to_unsigned(2,8) ,
46066	 => std_logic_vector(to_unsigned(2,8) ,
46067	 => std_logic_vector(to_unsigned(2,8) ,
46068	 => std_logic_vector(to_unsigned(2,8) ,
46069	 => std_logic_vector(to_unsigned(2,8) ,
46070	 => std_logic_vector(to_unsigned(2,8) ,
46071	 => std_logic_vector(to_unsigned(2,8) ,
46072	 => std_logic_vector(to_unsigned(3,8) ,
46073	 => std_logic_vector(to_unsigned(3,8) ,
46074	 => std_logic_vector(to_unsigned(2,8) ,
46075	 => std_logic_vector(to_unsigned(3,8) ,
46076	 => std_logic_vector(to_unsigned(2,8) ,
46077	 => std_logic_vector(to_unsigned(2,8) ,
46078	 => std_logic_vector(to_unsigned(2,8) ,
46079	 => std_logic_vector(to_unsigned(3,8) ,
46080	 => std_logic_vector(to_unsigned(3,8) ,
46081	 => std_logic_vector(to_unsigned(56,8) ,
46082	 => std_logic_vector(to_unsigned(62,8) ,
46083	 => std_logic_vector(to_unsigned(50,8) ,
46084	 => std_logic_vector(to_unsigned(50,8) ,
46085	 => std_logic_vector(to_unsigned(47,8) ,
46086	 => std_logic_vector(to_unsigned(52,8) ,
46087	 => std_logic_vector(to_unsigned(51,8) ,
46088	 => std_logic_vector(to_unsigned(45,8) ,
46089	 => std_logic_vector(to_unsigned(30,8) ,
46090	 => std_logic_vector(to_unsigned(28,8) ,
46091	 => std_logic_vector(to_unsigned(27,8) ,
46092	 => std_logic_vector(to_unsigned(30,8) ,
46093	 => std_logic_vector(to_unsigned(32,8) ,
46094	 => std_logic_vector(to_unsigned(49,8) ,
46095	 => std_logic_vector(to_unsigned(97,8) ,
46096	 => std_logic_vector(to_unsigned(114,8) ,
46097	 => std_logic_vector(to_unsigned(109,8) ,
46098	 => std_logic_vector(to_unsigned(101,8) ,
46099	 => std_logic_vector(to_unsigned(88,8) ,
46100	 => std_logic_vector(to_unsigned(111,8) ,
46101	 => std_logic_vector(to_unsigned(107,8) ,
46102	 => std_logic_vector(to_unsigned(111,8) ,
46103	 => std_logic_vector(to_unsigned(118,8) ,
46104	 => std_logic_vector(to_unsigned(118,8) ,
46105	 => std_logic_vector(to_unsigned(118,8) ,
46106	 => std_logic_vector(to_unsigned(125,8) ,
46107	 => std_logic_vector(to_unsigned(141,8) ,
46108	 => std_logic_vector(to_unsigned(136,8) ,
46109	 => std_logic_vector(to_unsigned(134,8) ,
46110	 => std_logic_vector(to_unsigned(131,8) ,
46111	 => std_logic_vector(to_unsigned(133,8) ,
46112	 => std_logic_vector(to_unsigned(142,8) ,
46113	 => std_logic_vector(to_unsigned(157,8) ,
46114	 => std_logic_vector(to_unsigned(154,8) ,
46115	 => std_logic_vector(to_unsigned(151,8) ,
46116	 => std_logic_vector(to_unsigned(159,8) ,
46117	 => std_logic_vector(to_unsigned(161,8) ,
46118	 => std_logic_vector(to_unsigned(154,8) ,
46119	 => std_logic_vector(to_unsigned(154,8) ,
46120	 => std_logic_vector(to_unsigned(157,8) ,
46121	 => std_logic_vector(to_unsigned(133,8) ,
46122	 => std_logic_vector(to_unsigned(88,8) ,
46123	 => std_logic_vector(to_unsigned(61,8) ,
46124	 => std_logic_vector(to_unsigned(70,8) ,
46125	 => std_logic_vector(to_unsigned(68,8) ,
46126	 => std_logic_vector(to_unsigned(58,8) ,
46127	 => std_logic_vector(to_unsigned(69,8) ,
46128	 => std_logic_vector(to_unsigned(76,8) ,
46129	 => std_logic_vector(to_unsigned(70,8) ,
46130	 => std_logic_vector(to_unsigned(82,8) ,
46131	 => std_logic_vector(to_unsigned(107,8) ,
46132	 => std_logic_vector(to_unsigned(91,8) ,
46133	 => std_logic_vector(to_unsigned(62,8) ,
46134	 => std_logic_vector(to_unsigned(78,8) ,
46135	 => std_logic_vector(to_unsigned(111,8) ,
46136	 => std_logic_vector(to_unsigned(104,8) ,
46137	 => std_logic_vector(to_unsigned(104,8) ,
46138	 => std_logic_vector(to_unsigned(107,8) ,
46139	 => std_logic_vector(to_unsigned(91,8) ,
46140	 => std_logic_vector(to_unsigned(87,8) ,
46141	 => std_logic_vector(to_unsigned(97,8) ,
46142	 => std_logic_vector(to_unsigned(74,8) ,
46143	 => std_logic_vector(to_unsigned(67,8) ,
46144	 => std_logic_vector(to_unsigned(60,8) ,
46145	 => std_logic_vector(to_unsigned(68,8) ,
46146	 => std_logic_vector(to_unsigned(71,8) ,
46147	 => std_logic_vector(to_unsigned(70,8) ,
46148	 => std_logic_vector(to_unsigned(70,8) ,
46149	 => std_logic_vector(to_unsigned(70,8) ,
46150	 => std_logic_vector(to_unsigned(76,8) ,
46151	 => std_logic_vector(to_unsigned(64,8) ,
46152	 => std_logic_vector(to_unsigned(51,8) ,
46153	 => std_logic_vector(to_unsigned(52,8) ,
46154	 => std_logic_vector(to_unsigned(49,8) ,
46155	 => std_logic_vector(to_unsigned(54,8) ,
46156	 => std_logic_vector(to_unsigned(85,8) ,
46157	 => std_logic_vector(to_unsigned(96,8) ,
46158	 => std_logic_vector(to_unsigned(80,8) ,
46159	 => std_logic_vector(to_unsigned(88,8) ,
46160	 => std_logic_vector(to_unsigned(92,8) ,
46161	 => std_logic_vector(to_unsigned(85,8) ,
46162	 => std_logic_vector(to_unsigned(77,8) ,
46163	 => std_logic_vector(to_unsigned(65,8) ,
46164	 => std_logic_vector(to_unsigned(79,8) ,
46165	 => std_logic_vector(to_unsigned(86,8) ,
46166	 => std_logic_vector(to_unsigned(65,8) ,
46167	 => std_logic_vector(to_unsigned(43,8) ,
46168	 => std_logic_vector(to_unsigned(53,8) ,
46169	 => std_logic_vector(to_unsigned(57,8) ,
46170	 => std_logic_vector(to_unsigned(48,8) ,
46171	 => std_logic_vector(to_unsigned(51,8) ,
46172	 => std_logic_vector(to_unsigned(56,8) ,
46173	 => std_logic_vector(to_unsigned(54,8) ,
46174	 => std_logic_vector(to_unsigned(57,8) ,
46175	 => std_logic_vector(to_unsigned(71,8) ,
46176	 => std_logic_vector(to_unsigned(80,8) ,
46177	 => std_logic_vector(to_unsigned(84,8) ,
46178	 => std_logic_vector(to_unsigned(77,8) ,
46179	 => std_logic_vector(to_unsigned(90,8) ,
46180	 => std_logic_vector(to_unsigned(97,8) ,
46181	 => std_logic_vector(to_unsigned(88,8) ,
46182	 => std_logic_vector(to_unsigned(69,8) ,
46183	 => std_logic_vector(to_unsigned(80,8) ,
46184	 => std_logic_vector(to_unsigned(85,8) ,
46185	 => std_logic_vector(to_unsigned(74,8) ,
46186	 => std_logic_vector(to_unsigned(77,8) ,
46187	 => std_logic_vector(to_unsigned(86,8) ,
46188	 => std_logic_vector(to_unsigned(73,8) ,
46189	 => std_logic_vector(to_unsigned(84,8) ,
46190	 => std_logic_vector(to_unsigned(84,8) ,
46191	 => std_logic_vector(to_unsigned(85,8) ,
46192	 => std_logic_vector(to_unsigned(85,8) ,
46193	 => std_logic_vector(to_unsigned(82,8) ,
46194	 => std_logic_vector(to_unsigned(91,8) ,
46195	 => std_logic_vector(to_unsigned(63,8) ,
46196	 => std_logic_vector(to_unsigned(53,8) ,
46197	 => std_logic_vector(to_unsigned(56,8) ,
46198	 => std_logic_vector(to_unsigned(57,8) ,
46199	 => std_logic_vector(to_unsigned(63,8) ,
46200	 => std_logic_vector(to_unsigned(58,8) ,
46201	 => std_logic_vector(to_unsigned(71,8) ,
46202	 => std_logic_vector(to_unsigned(76,8) ,
46203	 => std_logic_vector(to_unsigned(69,8) ,
46204	 => std_logic_vector(to_unsigned(64,8) ,
46205	 => std_logic_vector(to_unsigned(82,8) ,
46206	 => std_logic_vector(to_unsigned(90,8) ,
46207	 => std_logic_vector(to_unsigned(96,8) ,
46208	 => std_logic_vector(to_unsigned(115,8) ,
46209	 => std_logic_vector(to_unsigned(84,8) ,
46210	 => std_logic_vector(to_unsigned(87,8) ,
46211	 => std_logic_vector(to_unsigned(118,8) ,
46212	 => std_logic_vector(to_unsigned(112,8) ,
46213	 => std_logic_vector(to_unsigned(114,8) ,
46214	 => std_logic_vector(to_unsigned(97,8) ,
46215	 => std_logic_vector(to_unsigned(79,8) ,
46216	 => std_logic_vector(to_unsigned(60,8) ,
46217	 => std_logic_vector(to_unsigned(52,8) ,
46218	 => std_logic_vector(to_unsigned(59,8) ,
46219	 => std_logic_vector(to_unsigned(54,8) ,
46220	 => std_logic_vector(to_unsigned(65,8) ,
46221	 => std_logic_vector(to_unsigned(68,8) ,
46222	 => std_logic_vector(to_unsigned(61,8) ,
46223	 => std_logic_vector(to_unsigned(86,8) ,
46224	 => std_logic_vector(to_unsigned(85,8) ,
46225	 => std_logic_vector(to_unsigned(50,8) ,
46226	 => std_logic_vector(to_unsigned(42,8) ,
46227	 => std_logic_vector(to_unsigned(40,8) ,
46228	 => std_logic_vector(to_unsigned(44,8) ,
46229	 => std_logic_vector(to_unsigned(77,8) ,
46230	 => std_logic_vector(to_unsigned(121,8) ,
46231	 => std_logic_vector(to_unsigned(77,8) ,
46232	 => std_logic_vector(to_unsigned(41,8) ,
46233	 => std_logic_vector(to_unsigned(32,8) ,
46234	 => std_logic_vector(to_unsigned(15,8) ,
46235	 => std_logic_vector(to_unsigned(17,8) ,
46236	 => std_logic_vector(to_unsigned(29,8) ,
46237	 => std_logic_vector(to_unsigned(45,8) ,
46238	 => std_logic_vector(to_unsigned(46,8) ,
46239	 => std_logic_vector(to_unsigned(35,8) ,
46240	 => std_logic_vector(to_unsigned(39,8) ,
46241	 => std_logic_vector(to_unsigned(42,8) ,
46242	 => std_logic_vector(to_unsigned(37,8) ,
46243	 => std_logic_vector(to_unsigned(51,8) ,
46244	 => std_logic_vector(to_unsigned(36,8) ,
46245	 => std_logic_vector(to_unsigned(15,8) ,
46246	 => std_logic_vector(to_unsigned(13,8) ,
46247	 => std_logic_vector(to_unsigned(12,8) ,
46248	 => std_logic_vector(to_unsigned(20,8) ,
46249	 => std_logic_vector(to_unsigned(51,8) ,
46250	 => std_logic_vector(to_unsigned(59,8) ,
46251	 => std_logic_vector(to_unsigned(80,8) ,
46252	 => std_logic_vector(to_unsigned(44,8) ,
46253	 => std_logic_vector(to_unsigned(47,8) ,
46254	 => std_logic_vector(to_unsigned(61,8) ,
46255	 => std_logic_vector(to_unsigned(29,8) ,
46256	 => std_logic_vector(to_unsigned(27,8) ,
46257	 => std_logic_vector(to_unsigned(35,8) ,
46258	 => std_logic_vector(to_unsigned(34,8) ,
46259	 => std_logic_vector(to_unsigned(33,8) ,
46260	 => std_logic_vector(to_unsigned(27,8) ,
46261	 => std_logic_vector(to_unsigned(20,8) ,
46262	 => std_logic_vector(to_unsigned(37,8) ,
46263	 => std_logic_vector(to_unsigned(55,8) ,
46264	 => std_logic_vector(to_unsigned(48,8) ,
46265	 => std_logic_vector(to_unsigned(26,8) ,
46266	 => std_logic_vector(to_unsigned(22,8) ,
46267	 => std_logic_vector(to_unsigned(19,8) ,
46268	 => std_logic_vector(to_unsigned(13,8) ,
46269	 => std_logic_vector(to_unsigned(12,8) ,
46270	 => std_logic_vector(to_unsigned(43,8) ,
46271	 => std_logic_vector(to_unsigned(80,8) ,
46272	 => std_logic_vector(to_unsigned(53,8) ,
46273	 => std_logic_vector(to_unsigned(62,8) ,
46274	 => std_logic_vector(to_unsigned(72,8) ,
46275	 => std_logic_vector(to_unsigned(58,8) ,
46276	 => std_logic_vector(to_unsigned(57,8) ,
46277	 => std_logic_vector(to_unsigned(72,8) ,
46278	 => std_logic_vector(to_unsigned(82,8) ,
46279	 => std_logic_vector(to_unsigned(78,8) ,
46280	 => std_logic_vector(to_unsigned(82,8) ,
46281	 => std_logic_vector(to_unsigned(100,8) ,
46282	 => std_logic_vector(to_unsigned(95,8) ,
46283	 => std_logic_vector(to_unsigned(71,8) ,
46284	 => std_logic_vector(to_unsigned(85,8) ,
46285	 => std_logic_vector(to_unsigned(40,8) ,
46286	 => std_logic_vector(to_unsigned(8,8) ,
46287	 => std_logic_vector(to_unsigned(21,8) ,
46288	 => std_logic_vector(to_unsigned(37,8) ,
46289	 => std_logic_vector(to_unsigned(20,8) ,
46290	 => std_logic_vector(to_unsigned(3,8) ,
46291	 => std_logic_vector(to_unsigned(7,8) ,
46292	 => std_logic_vector(to_unsigned(24,8) ,
46293	 => std_logic_vector(to_unsigned(5,8) ,
46294	 => std_logic_vector(to_unsigned(9,8) ,
46295	 => std_logic_vector(to_unsigned(9,8) ,
46296	 => std_logic_vector(to_unsigned(4,8) ,
46297	 => std_logic_vector(to_unsigned(1,8) ,
46298	 => std_logic_vector(to_unsigned(23,8) ,
46299	 => std_logic_vector(to_unsigned(104,8) ,
46300	 => std_logic_vector(to_unsigned(85,8) ,
46301	 => std_logic_vector(to_unsigned(81,8) ,
46302	 => std_logic_vector(to_unsigned(87,8) ,
46303	 => std_logic_vector(to_unsigned(87,8) ,
46304	 => std_logic_vector(to_unsigned(87,8) ,
46305	 => std_logic_vector(to_unsigned(86,8) ,
46306	 => std_logic_vector(to_unsigned(84,8) ,
46307	 => std_logic_vector(to_unsigned(88,8) ,
46308	 => std_logic_vector(to_unsigned(104,8) ,
46309	 => std_logic_vector(to_unsigned(101,8) ,
46310	 => std_logic_vector(to_unsigned(49,8) ,
46311	 => std_logic_vector(to_unsigned(3,8) ,
46312	 => std_logic_vector(to_unsigned(7,8) ,
46313	 => std_logic_vector(to_unsigned(10,8) ,
46314	 => std_logic_vector(to_unsigned(7,8) ,
46315	 => std_logic_vector(to_unsigned(8,8) ,
46316	 => std_logic_vector(to_unsigned(1,8) ,
46317	 => std_logic_vector(to_unsigned(2,8) ,
46318	 => std_logic_vector(to_unsigned(4,8) ,
46319	 => std_logic_vector(to_unsigned(6,8) ,
46320	 => std_logic_vector(to_unsigned(6,8) ,
46321	 => std_logic_vector(to_unsigned(5,8) ,
46322	 => std_logic_vector(to_unsigned(1,8) ,
46323	 => std_logic_vector(to_unsigned(8,8) ,
46324	 => std_logic_vector(to_unsigned(111,8) ,
46325	 => std_logic_vector(to_unsigned(103,8) ,
46326	 => std_logic_vector(to_unsigned(101,8) ,
46327	 => std_logic_vector(to_unsigned(63,8) ,
46328	 => std_logic_vector(to_unsigned(6,8) ,
46329	 => std_logic_vector(to_unsigned(4,8) ,
46330	 => std_logic_vector(to_unsigned(74,8) ,
46331	 => std_logic_vector(to_unsigned(161,8) ,
46332	 => std_logic_vector(to_unsigned(142,8) ,
46333	 => std_logic_vector(to_unsigned(151,8) ,
46334	 => std_logic_vector(to_unsigned(142,8) ,
46335	 => std_logic_vector(to_unsigned(164,8) ,
46336	 => std_logic_vector(to_unsigned(86,8) ,
46337	 => std_logic_vector(to_unsigned(4,8) ,
46338	 => std_logic_vector(to_unsigned(3,8) ,
46339	 => std_logic_vector(to_unsigned(4,8) ,
46340	 => std_logic_vector(to_unsigned(2,8) ,
46341	 => std_logic_vector(to_unsigned(1,8) ,
46342	 => std_logic_vector(to_unsigned(0,8) ,
46343	 => std_logic_vector(to_unsigned(37,8) ,
46344	 => std_logic_vector(to_unsigned(186,8) ,
46345	 => std_logic_vector(to_unsigned(149,8) ,
46346	 => std_logic_vector(to_unsigned(141,8) ,
46347	 => std_logic_vector(to_unsigned(166,8) ,
46348	 => std_logic_vector(to_unsigned(173,8) ,
46349	 => std_logic_vector(to_unsigned(53,8) ,
46350	 => std_logic_vector(to_unsigned(1,8) ,
46351	 => std_logic_vector(to_unsigned(5,8) ,
46352	 => std_logic_vector(to_unsigned(11,8) ,
46353	 => std_logic_vector(to_unsigned(6,8) ,
46354	 => std_logic_vector(to_unsigned(1,8) ,
46355	 => std_logic_vector(to_unsigned(1,8) ,
46356	 => std_logic_vector(to_unsigned(2,8) ,
46357	 => std_logic_vector(to_unsigned(5,8) ,
46358	 => std_logic_vector(to_unsigned(4,8) ,
46359	 => std_logic_vector(to_unsigned(1,8) ,
46360	 => std_logic_vector(to_unsigned(1,8) ,
46361	 => std_logic_vector(to_unsigned(1,8) ,
46362	 => std_logic_vector(to_unsigned(1,8) ,
46363	 => std_logic_vector(to_unsigned(2,8) ,
46364	 => std_logic_vector(to_unsigned(2,8) ,
46365	 => std_logic_vector(to_unsigned(4,8) ,
46366	 => std_logic_vector(to_unsigned(7,8) ,
46367	 => std_logic_vector(to_unsigned(8,8) ,
46368	 => std_logic_vector(to_unsigned(5,8) ,
46369	 => std_logic_vector(to_unsigned(2,8) ,
46370	 => std_logic_vector(to_unsigned(2,8) ,
46371	 => std_logic_vector(to_unsigned(2,8) ,
46372	 => std_logic_vector(to_unsigned(1,8) ,
46373	 => std_logic_vector(to_unsigned(2,8) ,
46374	 => std_logic_vector(to_unsigned(2,8) ,
46375	 => std_logic_vector(to_unsigned(2,8) ,
46376	 => std_logic_vector(to_unsigned(4,8) ,
46377	 => std_logic_vector(to_unsigned(4,8) ,
46378	 => std_logic_vector(to_unsigned(3,8) ,
46379	 => std_logic_vector(to_unsigned(4,8) ,
46380	 => std_logic_vector(to_unsigned(3,8) ,
46381	 => std_logic_vector(to_unsigned(4,8) ,
46382	 => std_logic_vector(to_unsigned(3,8) ,
46383	 => std_logic_vector(to_unsigned(4,8) ,
46384	 => std_logic_vector(to_unsigned(5,8) ,
46385	 => std_logic_vector(to_unsigned(5,8) ,
46386	 => std_logic_vector(to_unsigned(4,8) ,
46387	 => std_logic_vector(to_unsigned(4,8) ,
46388	 => std_logic_vector(to_unsigned(4,8) ,
46389	 => std_logic_vector(to_unsigned(3,8) ,
46390	 => std_logic_vector(to_unsigned(3,8) ,
46391	 => std_logic_vector(to_unsigned(3,8) ,
46392	 => std_logic_vector(to_unsigned(3,8) ,
46393	 => std_logic_vector(to_unsigned(3,8) ,
46394	 => std_logic_vector(to_unsigned(2,8) ,
46395	 => std_logic_vector(to_unsigned(3,8) ,
46396	 => std_logic_vector(to_unsigned(2,8) ,
46397	 => std_logic_vector(to_unsigned(3,8) ,
46398	 => std_logic_vector(to_unsigned(3,8) ,
46399	 => std_logic_vector(to_unsigned(2,8) ,
46400	 => std_logic_vector(to_unsigned(2,8) ,
46401	 => std_logic_vector(to_unsigned(54,8) ,
46402	 => std_logic_vector(to_unsigned(53,8) ,
46403	 => std_logic_vector(to_unsigned(49,8) ,
46404	 => std_logic_vector(to_unsigned(47,8) ,
46405	 => std_logic_vector(to_unsigned(50,8) ,
46406	 => std_logic_vector(to_unsigned(55,8) ,
46407	 => std_logic_vector(to_unsigned(51,8) ,
46408	 => std_logic_vector(to_unsigned(53,8) ,
46409	 => std_logic_vector(to_unsigned(32,8) ,
46410	 => std_logic_vector(to_unsigned(29,8) ,
46411	 => std_logic_vector(to_unsigned(29,8) ,
46412	 => std_logic_vector(to_unsigned(26,8) ,
46413	 => std_logic_vector(to_unsigned(32,8) ,
46414	 => std_logic_vector(to_unsigned(36,8) ,
46415	 => std_logic_vector(to_unsigned(86,8) ,
46416	 => std_logic_vector(to_unsigned(116,8) ,
46417	 => std_logic_vector(to_unsigned(101,8) ,
46418	 => std_logic_vector(to_unsigned(103,8) ,
46419	 => std_logic_vector(to_unsigned(95,8) ,
46420	 => std_logic_vector(to_unsigned(109,8) ,
46421	 => std_logic_vector(to_unsigned(115,8) ,
46422	 => std_logic_vector(to_unsigned(108,8) ,
46423	 => std_logic_vector(to_unsigned(107,8) ,
46424	 => std_logic_vector(to_unsigned(107,8) ,
46425	 => std_logic_vector(to_unsigned(114,8) ,
46426	 => std_logic_vector(to_unsigned(118,8) ,
46427	 => std_logic_vector(to_unsigned(114,8) ,
46428	 => std_logic_vector(to_unsigned(118,8) ,
46429	 => std_logic_vector(to_unsigned(119,8) ,
46430	 => std_logic_vector(to_unsigned(114,8) ,
46431	 => std_logic_vector(to_unsigned(131,8) ,
46432	 => std_logic_vector(to_unsigned(146,8) ,
46433	 => std_logic_vector(to_unsigned(156,8) ,
46434	 => std_logic_vector(to_unsigned(156,8) ,
46435	 => std_logic_vector(to_unsigned(154,8) ,
46436	 => std_logic_vector(to_unsigned(159,8) ,
46437	 => std_logic_vector(to_unsigned(159,8) ,
46438	 => std_logic_vector(to_unsigned(159,8) ,
46439	 => std_logic_vector(to_unsigned(152,8) ,
46440	 => std_logic_vector(to_unsigned(156,8) ,
46441	 => std_logic_vector(to_unsigned(139,8) ,
46442	 => std_logic_vector(to_unsigned(90,8) ,
46443	 => std_logic_vector(to_unsigned(69,8) ,
46444	 => std_logic_vector(to_unsigned(65,8) ,
46445	 => std_logic_vector(to_unsigned(55,8) ,
46446	 => std_logic_vector(to_unsigned(63,8) ,
46447	 => std_logic_vector(to_unsigned(77,8) ,
46448	 => std_logic_vector(to_unsigned(81,8) ,
46449	 => std_logic_vector(to_unsigned(88,8) ,
46450	 => std_logic_vector(to_unsigned(105,8) ,
46451	 => std_logic_vector(to_unsigned(107,8) ,
46452	 => std_logic_vector(to_unsigned(76,8) ,
46453	 => std_logic_vector(to_unsigned(63,8) ,
46454	 => std_logic_vector(to_unsigned(76,8) ,
46455	 => std_logic_vector(to_unsigned(78,8) ,
46456	 => std_logic_vector(to_unsigned(97,8) ,
46457	 => std_logic_vector(to_unsigned(109,8) ,
46458	 => std_logic_vector(to_unsigned(112,8) ,
46459	 => std_logic_vector(to_unsigned(96,8) ,
46460	 => std_logic_vector(to_unsigned(85,8) ,
46461	 => std_logic_vector(to_unsigned(95,8) ,
46462	 => std_logic_vector(to_unsigned(69,8) ,
46463	 => std_logic_vector(to_unsigned(64,8) ,
46464	 => std_logic_vector(to_unsigned(58,8) ,
46465	 => std_logic_vector(to_unsigned(59,8) ,
46466	 => std_logic_vector(to_unsigned(64,8) ,
46467	 => std_logic_vector(to_unsigned(59,8) ,
46468	 => std_logic_vector(to_unsigned(56,8) ,
46469	 => std_logic_vector(to_unsigned(60,8) ,
46470	 => std_logic_vector(to_unsigned(58,8) ,
46471	 => std_logic_vector(to_unsigned(57,8) ,
46472	 => std_logic_vector(to_unsigned(53,8) ,
46473	 => std_logic_vector(to_unsigned(51,8) ,
46474	 => std_logic_vector(to_unsigned(49,8) ,
46475	 => std_logic_vector(to_unsigned(49,8) ,
46476	 => std_logic_vector(to_unsigned(79,8) ,
46477	 => std_logic_vector(to_unsigned(95,8) ,
46478	 => std_logic_vector(to_unsigned(90,8) ,
46479	 => std_logic_vector(to_unsigned(86,8) ,
46480	 => std_logic_vector(to_unsigned(84,8) ,
46481	 => std_logic_vector(to_unsigned(80,8) ,
46482	 => std_logic_vector(to_unsigned(79,8) ,
46483	 => std_logic_vector(to_unsigned(72,8) ,
46484	 => std_logic_vector(to_unsigned(91,8) ,
46485	 => std_logic_vector(to_unsigned(90,8) ,
46486	 => std_logic_vector(to_unsigned(59,8) ,
46487	 => std_logic_vector(to_unsigned(39,8) ,
46488	 => std_logic_vector(to_unsigned(50,8) ,
46489	 => std_logic_vector(to_unsigned(51,8) ,
46490	 => std_logic_vector(to_unsigned(42,8) ,
46491	 => std_logic_vector(to_unsigned(45,8) ,
46492	 => std_logic_vector(to_unsigned(58,8) ,
46493	 => std_logic_vector(to_unsigned(57,8) ,
46494	 => std_logic_vector(to_unsigned(54,8) ,
46495	 => std_logic_vector(to_unsigned(74,8) ,
46496	 => std_logic_vector(to_unsigned(74,8) ,
46497	 => std_logic_vector(to_unsigned(69,8) ,
46498	 => std_logic_vector(to_unsigned(77,8) ,
46499	 => std_logic_vector(to_unsigned(79,8) ,
46500	 => std_logic_vector(to_unsigned(77,8) ,
46501	 => std_logic_vector(to_unsigned(69,8) ,
46502	 => std_logic_vector(to_unsigned(68,8) ,
46503	 => std_logic_vector(to_unsigned(74,8) ,
46504	 => std_logic_vector(to_unsigned(79,8) ,
46505	 => std_logic_vector(to_unsigned(81,8) ,
46506	 => std_logic_vector(to_unsigned(80,8) ,
46507	 => std_logic_vector(to_unsigned(70,8) ,
46508	 => std_logic_vector(to_unsigned(71,8) ,
46509	 => std_logic_vector(to_unsigned(73,8) ,
46510	 => std_logic_vector(to_unsigned(68,8) ,
46511	 => std_logic_vector(to_unsigned(56,8) ,
46512	 => std_logic_vector(to_unsigned(54,8) ,
46513	 => std_logic_vector(to_unsigned(74,8) ,
46514	 => std_logic_vector(to_unsigned(114,8) ,
46515	 => std_logic_vector(to_unsigned(88,8) ,
46516	 => std_logic_vector(to_unsigned(60,8) ,
46517	 => std_logic_vector(to_unsigned(69,8) ,
46518	 => std_logic_vector(to_unsigned(62,8) ,
46519	 => std_logic_vector(to_unsigned(61,8) ,
46520	 => std_logic_vector(to_unsigned(57,8) ,
46521	 => std_logic_vector(to_unsigned(57,8) ,
46522	 => std_logic_vector(to_unsigned(59,8) ,
46523	 => std_logic_vector(to_unsigned(62,8) ,
46524	 => std_logic_vector(to_unsigned(63,8) ,
46525	 => std_logic_vector(to_unsigned(87,8) ,
46526	 => std_logic_vector(to_unsigned(97,8) ,
46527	 => std_logic_vector(to_unsigned(95,8) ,
46528	 => std_logic_vector(to_unsigned(96,8) ,
46529	 => std_logic_vector(to_unsigned(91,8) ,
46530	 => std_logic_vector(to_unsigned(91,8) ,
46531	 => std_logic_vector(to_unsigned(103,8) ,
46532	 => std_logic_vector(to_unsigned(111,8) ,
46533	 => std_logic_vector(to_unsigned(107,8) ,
46534	 => std_logic_vector(to_unsigned(92,8) ,
46535	 => std_logic_vector(to_unsigned(81,8) ,
46536	 => std_logic_vector(to_unsigned(59,8) ,
46537	 => std_logic_vector(to_unsigned(45,8) ,
46538	 => std_logic_vector(to_unsigned(40,8) ,
46539	 => std_logic_vector(to_unsigned(49,8) ,
46540	 => std_logic_vector(to_unsigned(61,8) ,
46541	 => std_logic_vector(to_unsigned(71,8) ,
46542	 => std_logic_vector(to_unsigned(72,8) ,
46543	 => std_logic_vector(to_unsigned(76,8) ,
46544	 => std_logic_vector(to_unsigned(95,8) ,
46545	 => std_logic_vector(to_unsigned(64,8) ,
46546	 => std_logic_vector(to_unsigned(42,8) ,
46547	 => std_logic_vector(to_unsigned(69,8) ,
46548	 => std_logic_vector(to_unsigned(101,8) ,
46549	 => std_logic_vector(to_unsigned(115,8) ,
46550	 => std_logic_vector(to_unsigned(108,8) ,
46551	 => std_logic_vector(to_unsigned(90,8) ,
46552	 => std_logic_vector(to_unsigned(70,8) ,
46553	 => std_logic_vector(to_unsigned(38,8) ,
46554	 => std_logic_vector(to_unsigned(32,8) ,
46555	 => std_logic_vector(to_unsigned(23,8) ,
46556	 => std_logic_vector(to_unsigned(32,8) ,
46557	 => std_logic_vector(to_unsigned(54,8) ,
46558	 => std_logic_vector(to_unsigned(57,8) ,
46559	 => std_logic_vector(to_unsigned(66,8) ,
46560	 => std_logic_vector(to_unsigned(76,8) ,
46561	 => std_logic_vector(to_unsigned(37,8) ,
46562	 => std_logic_vector(to_unsigned(46,8) ,
46563	 => std_logic_vector(to_unsigned(68,8) ,
46564	 => std_logic_vector(to_unsigned(27,8) ,
46565	 => std_logic_vector(to_unsigned(17,8) ,
46566	 => std_logic_vector(to_unsigned(15,8) ,
46567	 => std_logic_vector(to_unsigned(23,8) ,
46568	 => std_logic_vector(to_unsigned(22,8) ,
46569	 => std_logic_vector(to_unsigned(16,8) ,
46570	 => std_logic_vector(to_unsigned(25,8) ,
46571	 => std_logic_vector(to_unsigned(41,8) ,
46572	 => std_logic_vector(to_unsigned(27,8) ,
46573	 => std_logic_vector(to_unsigned(33,8) ,
46574	 => std_logic_vector(to_unsigned(38,8) ,
46575	 => std_logic_vector(to_unsigned(26,8) ,
46576	 => std_logic_vector(to_unsigned(23,8) ,
46577	 => std_logic_vector(to_unsigned(23,8) ,
46578	 => std_logic_vector(to_unsigned(30,8) ,
46579	 => std_logic_vector(to_unsigned(36,8) ,
46580	 => std_logic_vector(to_unsigned(40,8) ,
46581	 => std_logic_vector(to_unsigned(43,8) ,
46582	 => std_logic_vector(to_unsigned(48,8) ,
46583	 => std_logic_vector(to_unsigned(59,8) ,
46584	 => std_logic_vector(to_unsigned(37,8) ,
46585	 => std_logic_vector(to_unsigned(27,8) ,
46586	 => std_logic_vector(to_unsigned(18,8) ,
46587	 => std_logic_vector(to_unsigned(15,8) ,
46588	 => std_logic_vector(to_unsigned(13,8) ,
46589	 => std_logic_vector(to_unsigned(11,8) ,
46590	 => std_logic_vector(to_unsigned(35,8) ,
46591	 => std_logic_vector(to_unsigned(79,8) ,
46592	 => std_logic_vector(to_unsigned(65,8) ,
46593	 => std_logic_vector(to_unsigned(65,8) ,
46594	 => std_logic_vector(to_unsigned(61,8) ,
46595	 => std_logic_vector(to_unsigned(60,8) ,
46596	 => std_logic_vector(to_unsigned(52,8) ,
46597	 => std_logic_vector(to_unsigned(64,8) ,
46598	 => std_logic_vector(to_unsigned(70,8) ,
46599	 => std_logic_vector(to_unsigned(53,8) ,
46600	 => std_logic_vector(to_unsigned(65,8) ,
46601	 => std_logic_vector(to_unsigned(101,8) ,
46602	 => std_logic_vector(to_unsigned(103,8) ,
46603	 => std_logic_vector(to_unsigned(59,8) ,
46604	 => std_logic_vector(to_unsigned(62,8) ,
46605	 => std_logic_vector(to_unsigned(30,8) ,
46606	 => std_logic_vector(to_unsigned(6,8) ,
46607	 => std_logic_vector(to_unsigned(17,8) ,
46608	 => std_logic_vector(to_unsigned(30,8) ,
46609	 => std_logic_vector(to_unsigned(8,8) ,
46610	 => std_logic_vector(to_unsigned(1,8) ,
46611	 => std_logic_vector(to_unsigned(25,8) ,
46612	 => std_logic_vector(to_unsigned(29,8) ,
46613	 => std_logic_vector(to_unsigned(2,8) ,
46614	 => std_logic_vector(to_unsigned(6,8) ,
46615	 => std_logic_vector(to_unsigned(6,8) ,
46616	 => std_logic_vector(to_unsigned(3,8) ,
46617	 => std_logic_vector(to_unsigned(5,8) ,
46618	 => std_logic_vector(to_unsigned(59,8) ,
46619	 => std_logic_vector(to_unsigned(108,8) ,
46620	 => std_logic_vector(to_unsigned(101,8) ,
46621	 => std_logic_vector(to_unsigned(82,8) ,
46622	 => std_logic_vector(to_unsigned(78,8) ,
46623	 => std_logic_vector(to_unsigned(76,8) ,
46624	 => std_logic_vector(to_unsigned(74,8) ,
46625	 => std_logic_vector(to_unsigned(79,8) ,
46626	 => std_logic_vector(to_unsigned(81,8) ,
46627	 => std_logic_vector(to_unsigned(78,8) ,
46628	 => std_logic_vector(to_unsigned(86,8) ,
46629	 => std_logic_vector(to_unsigned(87,8) ,
46630	 => std_logic_vector(to_unsigned(21,8) ,
46631	 => std_logic_vector(to_unsigned(4,8) ,
46632	 => std_logic_vector(to_unsigned(8,8) ,
46633	 => std_logic_vector(to_unsigned(12,8) ,
46634	 => std_logic_vector(to_unsigned(13,8) ,
46635	 => std_logic_vector(to_unsigned(3,8) ,
46636	 => std_logic_vector(to_unsigned(1,8) ,
46637	 => std_logic_vector(to_unsigned(5,8) ,
46638	 => std_logic_vector(to_unsigned(4,8) ,
46639	 => std_logic_vector(to_unsigned(4,8) ,
46640	 => std_logic_vector(to_unsigned(5,8) ,
46641	 => std_logic_vector(to_unsigned(3,8) ,
46642	 => std_logic_vector(to_unsigned(0,8) ,
46643	 => std_logic_vector(to_unsigned(18,8) ,
46644	 => std_logic_vector(to_unsigned(115,8) ,
46645	 => std_logic_vector(to_unsigned(104,8) ,
46646	 => std_logic_vector(to_unsigned(116,8) ,
46647	 => std_logic_vector(to_unsigned(91,8) ,
46648	 => std_logic_vector(to_unsigned(9,8) ,
46649	 => std_logic_vector(to_unsigned(5,8) ,
46650	 => std_logic_vector(to_unsigned(66,8) ,
46651	 => std_logic_vector(to_unsigned(141,8) ,
46652	 => std_logic_vector(to_unsigned(122,8) ,
46653	 => std_logic_vector(to_unsigned(124,8) ,
46654	 => std_logic_vector(to_unsigned(122,8) ,
46655	 => std_logic_vector(to_unsigned(149,8) ,
46656	 => std_logic_vector(to_unsigned(54,8) ,
46657	 => std_logic_vector(to_unsigned(2,8) ,
46658	 => std_logic_vector(to_unsigned(5,8) ,
46659	 => std_logic_vector(to_unsigned(7,8) ,
46660	 => std_logic_vector(to_unsigned(4,8) ,
46661	 => std_logic_vector(to_unsigned(2,8) ,
46662	 => std_logic_vector(to_unsigned(0,8) ,
46663	 => std_logic_vector(to_unsigned(30,8) ,
46664	 => std_logic_vector(to_unsigned(163,8) ,
46665	 => std_logic_vector(to_unsigned(144,8) ,
46666	 => std_logic_vector(to_unsigned(154,8) ,
46667	 => std_logic_vector(to_unsigned(168,8) ,
46668	 => std_logic_vector(to_unsigned(173,8) ,
46669	 => std_logic_vector(to_unsigned(24,8) ,
46670	 => std_logic_vector(to_unsigned(2,8) ,
46671	 => std_logic_vector(to_unsigned(6,8) ,
46672	 => std_logic_vector(to_unsigned(11,8) ,
46673	 => std_logic_vector(to_unsigned(7,8) ,
46674	 => std_logic_vector(to_unsigned(2,8) ,
46675	 => std_logic_vector(to_unsigned(1,8) ,
46676	 => std_logic_vector(to_unsigned(1,8) ,
46677	 => std_logic_vector(to_unsigned(3,8) ,
46678	 => std_logic_vector(to_unsigned(25,8) ,
46679	 => std_logic_vector(to_unsigned(50,8) ,
46680	 => std_logic_vector(to_unsigned(31,8) ,
46681	 => std_logic_vector(to_unsigned(38,8) ,
46682	 => std_logic_vector(to_unsigned(13,8) ,
46683	 => std_logic_vector(to_unsigned(2,8) ,
46684	 => std_logic_vector(to_unsigned(4,8) ,
46685	 => std_logic_vector(to_unsigned(4,8) ,
46686	 => std_logic_vector(to_unsigned(4,8) ,
46687	 => std_logic_vector(to_unsigned(4,8) ,
46688	 => std_logic_vector(to_unsigned(3,8) ,
46689	 => std_logic_vector(to_unsigned(1,8) ,
46690	 => std_logic_vector(to_unsigned(2,8) ,
46691	 => std_logic_vector(to_unsigned(2,8) ,
46692	 => std_logic_vector(to_unsigned(1,8) ,
46693	 => std_logic_vector(to_unsigned(1,8) ,
46694	 => std_logic_vector(to_unsigned(1,8) ,
46695	 => std_logic_vector(to_unsigned(1,8) ,
46696	 => std_logic_vector(to_unsigned(1,8) ,
46697	 => std_logic_vector(to_unsigned(1,8) ,
46698	 => std_logic_vector(to_unsigned(2,8) ,
46699	 => std_logic_vector(to_unsigned(4,8) ,
46700	 => std_logic_vector(to_unsigned(4,8) ,
46701	 => std_logic_vector(to_unsigned(4,8) ,
46702	 => std_logic_vector(to_unsigned(3,8) ,
46703	 => std_logic_vector(to_unsigned(2,8) ,
46704	 => std_logic_vector(to_unsigned(5,8) ,
46705	 => std_logic_vector(to_unsigned(6,8) ,
46706	 => std_logic_vector(to_unsigned(5,8) ,
46707	 => std_logic_vector(to_unsigned(5,8) ,
46708	 => std_logic_vector(to_unsigned(4,8) ,
46709	 => std_logic_vector(to_unsigned(5,8) ,
46710	 => std_logic_vector(to_unsigned(5,8) ,
46711	 => std_logic_vector(to_unsigned(5,8) ,
46712	 => std_logic_vector(to_unsigned(5,8) ,
46713	 => std_logic_vector(to_unsigned(5,8) ,
46714	 => std_logic_vector(to_unsigned(6,8) ,
46715	 => std_logic_vector(to_unsigned(7,8) ,
46716	 => std_logic_vector(to_unsigned(6,8) ,
46717	 => std_logic_vector(to_unsigned(4,8) ,
46718	 => std_logic_vector(to_unsigned(5,8) ,
46719	 => std_logic_vector(to_unsigned(4,8) ,
46720	 => std_logic_vector(to_unsigned(3,8) ,
46721	 => std_logic_vector(to_unsigned(49,8) ,
46722	 => std_logic_vector(to_unsigned(51,8) ,
46723	 => std_logic_vector(to_unsigned(54,8) ,
46724	 => std_logic_vector(to_unsigned(58,8) ,
46725	 => std_logic_vector(to_unsigned(55,8) ,
46726	 => std_logic_vector(to_unsigned(56,8) ,
46727	 => std_logic_vector(to_unsigned(46,8) ,
46728	 => std_logic_vector(to_unsigned(48,8) ,
46729	 => std_logic_vector(to_unsigned(38,8) ,
46730	 => std_logic_vector(to_unsigned(30,8) ,
46731	 => std_logic_vector(to_unsigned(28,8) ,
46732	 => std_logic_vector(to_unsigned(25,8) ,
46733	 => std_logic_vector(to_unsigned(27,8) ,
46734	 => std_logic_vector(to_unsigned(32,8) ,
46735	 => std_logic_vector(to_unsigned(78,8) ,
46736	 => std_logic_vector(to_unsigned(101,8) ,
46737	 => std_logic_vector(to_unsigned(99,8) ,
46738	 => std_logic_vector(to_unsigned(103,8) ,
46739	 => std_logic_vector(to_unsigned(92,8) ,
46740	 => std_logic_vector(to_unsigned(99,8) ,
46741	 => std_logic_vector(to_unsigned(111,8) ,
46742	 => std_logic_vector(to_unsigned(109,8) ,
46743	 => std_logic_vector(to_unsigned(100,8) ,
46744	 => std_logic_vector(to_unsigned(112,8) ,
46745	 => std_logic_vector(to_unsigned(121,8) ,
46746	 => std_logic_vector(to_unsigned(130,8) ,
46747	 => std_logic_vector(to_unsigned(127,8) ,
46748	 => std_logic_vector(to_unsigned(109,8) ,
46749	 => std_logic_vector(to_unsigned(115,8) ,
46750	 => std_logic_vector(to_unsigned(119,8) ,
46751	 => std_logic_vector(to_unsigned(131,8) ,
46752	 => std_logic_vector(to_unsigned(136,8) ,
46753	 => std_logic_vector(to_unsigned(151,8) ,
46754	 => std_logic_vector(to_unsigned(156,8) ,
46755	 => std_logic_vector(to_unsigned(156,8) ,
46756	 => std_logic_vector(to_unsigned(157,8) ,
46757	 => std_logic_vector(to_unsigned(159,8) ,
46758	 => std_logic_vector(to_unsigned(156,8) ,
46759	 => std_logic_vector(to_unsigned(156,8) ,
46760	 => std_logic_vector(to_unsigned(156,8) ,
46761	 => std_logic_vector(to_unsigned(146,8) ,
46762	 => std_logic_vector(to_unsigned(100,8) ,
46763	 => std_logic_vector(to_unsigned(70,8) ,
46764	 => std_logic_vector(to_unsigned(65,8) ,
46765	 => std_logic_vector(to_unsigned(61,8) ,
46766	 => std_logic_vector(to_unsigned(66,8) ,
46767	 => std_logic_vector(to_unsigned(73,8) ,
46768	 => std_logic_vector(to_unsigned(81,8) ,
46769	 => std_logic_vector(to_unsigned(93,8) ,
46770	 => std_logic_vector(to_unsigned(97,8) ,
46771	 => std_logic_vector(to_unsigned(82,8) ,
46772	 => std_logic_vector(to_unsigned(60,8) ,
46773	 => std_logic_vector(to_unsigned(73,8) ,
46774	 => std_logic_vector(to_unsigned(99,8) ,
46775	 => std_logic_vector(to_unsigned(92,8) ,
46776	 => std_logic_vector(to_unsigned(99,8) ,
46777	 => std_logic_vector(to_unsigned(96,8) ,
46778	 => std_logic_vector(to_unsigned(97,8) ,
46779	 => std_logic_vector(to_unsigned(104,8) ,
46780	 => std_logic_vector(to_unsigned(86,8) ,
46781	 => std_logic_vector(to_unsigned(86,8) ,
46782	 => std_logic_vector(to_unsigned(64,8) ,
46783	 => std_logic_vector(to_unsigned(55,8) ,
46784	 => std_logic_vector(to_unsigned(51,8) ,
46785	 => std_logic_vector(to_unsigned(57,8) ,
46786	 => std_logic_vector(to_unsigned(63,8) ,
46787	 => std_logic_vector(to_unsigned(53,8) ,
46788	 => std_logic_vector(to_unsigned(55,8) ,
46789	 => std_logic_vector(to_unsigned(53,8) ,
46790	 => std_logic_vector(to_unsigned(48,8) ,
46791	 => std_logic_vector(to_unsigned(56,8) ,
46792	 => std_logic_vector(to_unsigned(59,8) ,
46793	 => std_logic_vector(to_unsigned(50,8) ,
46794	 => std_logic_vector(to_unsigned(48,8) ,
46795	 => std_logic_vector(to_unsigned(47,8) ,
46796	 => std_logic_vector(to_unsigned(73,8) ,
46797	 => std_logic_vector(to_unsigned(93,8) ,
46798	 => std_logic_vector(to_unsigned(81,8) ,
46799	 => std_logic_vector(to_unsigned(77,8) ,
46800	 => std_logic_vector(to_unsigned(81,8) ,
46801	 => std_logic_vector(to_unsigned(73,8) ,
46802	 => std_logic_vector(to_unsigned(74,8) ,
46803	 => std_logic_vector(to_unsigned(70,8) ,
46804	 => std_logic_vector(to_unsigned(90,8) ,
46805	 => std_logic_vector(to_unsigned(72,8) ,
46806	 => std_logic_vector(to_unsigned(53,8) ,
46807	 => std_logic_vector(to_unsigned(51,8) ,
46808	 => std_logic_vector(to_unsigned(51,8) ,
46809	 => std_logic_vector(to_unsigned(44,8) ,
46810	 => std_logic_vector(to_unsigned(45,8) ,
46811	 => std_logic_vector(to_unsigned(48,8) ,
46812	 => std_logic_vector(to_unsigned(59,8) ,
46813	 => std_logic_vector(to_unsigned(62,8) ,
46814	 => std_logic_vector(to_unsigned(52,8) ,
46815	 => std_logic_vector(to_unsigned(67,8) ,
46816	 => std_logic_vector(to_unsigned(69,8) ,
46817	 => std_logic_vector(to_unsigned(60,8) ,
46818	 => std_logic_vector(to_unsigned(62,8) ,
46819	 => std_logic_vector(to_unsigned(71,8) ,
46820	 => std_logic_vector(to_unsigned(71,8) ,
46821	 => std_logic_vector(to_unsigned(66,8) ,
46822	 => std_logic_vector(to_unsigned(71,8) ,
46823	 => std_logic_vector(to_unsigned(71,8) ,
46824	 => std_logic_vector(to_unsigned(97,8) ,
46825	 => std_logic_vector(to_unsigned(103,8) ,
46826	 => std_logic_vector(to_unsigned(93,8) ,
46827	 => std_logic_vector(to_unsigned(88,8) ,
46828	 => std_logic_vector(to_unsigned(88,8) ,
46829	 => std_logic_vector(to_unsigned(84,8) ,
46830	 => std_logic_vector(to_unsigned(68,8) ,
46831	 => std_logic_vector(to_unsigned(63,8) ,
46832	 => std_logic_vector(to_unsigned(93,8) ,
46833	 => std_logic_vector(to_unsigned(95,8) ,
46834	 => std_logic_vector(to_unsigned(95,8) ,
46835	 => std_logic_vector(to_unsigned(88,8) ,
46836	 => std_logic_vector(to_unsigned(63,8) ,
46837	 => std_logic_vector(to_unsigned(68,8) ,
46838	 => std_logic_vector(to_unsigned(69,8) ,
46839	 => std_logic_vector(to_unsigned(69,8) ,
46840	 => std_logic_vector(to_unsigned(57,8) ,
46841	 => std_logic_vector(to_unsigned(58,8) ,
46842	 => std_logic_vector(to_unsigned(53,8) ,
46843	 => std_logic_vector(to_unsigned(57,8) ,
46844	 => std_logic_vector(to_unsigned(64,8) ,
46845	 => std_logic_vector(to_unsigned(81,8) ,
46846	 => std_logic_vector(to_unsigned(78,8) ,
46847	 => std_logic_vector(to_unsigned(93,8) ,
46848	 => std_logic_vector(to_unsigned(97,8) ,
46849	 => std_logic_vector(to_unsigned(77,8) ,
46850	 => std_logic_vector(to_unsigned(77,8) ,
46851	 => std_logic_vector(to_unsigned(103,8) ,
46852	 => std_logic_vector(to_unsigned(93,8) ,
46853	 => std_logic_vector(to_unsigned(86,8) ,
46854	 => std_logic_vector(to_unsigned(86,8) ,
46855	 => std_logic_vector(to_unsigned(79,8) ,
46856	 => std_logic_vector(to_unsigned(58,8) ,
46857	 => std_logic_vector(to_unsigned(41,8) ,
46858	 => std_logic_vector(to_unsigned(37,8) ,
46859	 => std_logic_vector(to_unsigned(46,8) ,
46860	 => std_logic_vector(to_unsigned(64,8) ,
46861	 => std_logic_vector(to_unsigned(79,8) ,
46862	 => std_logic_vector(to_unsigned(78,8) ,
46863	 => std_logic_vector(to_unsigned(80,8) ,
46864	 => std_logic_vector(to_unsigned(88,8) ,
46865	 => std_logic_vector(to_unsigned(65,8) ,
46866	 => std_logic_vector(to_unsigned(34,8) ,
46867	 => std_logic_vector(to_unsigned(51,8) ,
46868	 => std_logic_vector(to_unsigned(53,8) ,
46869	 => std_logic_vector(to_unsigned(65,8) ,
46870	 => std_logic_vector(to_unsigned(61,8) ,
46871	 => std_logic_vector(to_unsigned(37,8) ,
46872	 => std_logic_vector(to_unsigned(25,8) ,
46873	 => std_logic_vector(to_unsigned(20,8) ,
46874	 => std_logic_vector(to_unsigned(24,8) ,
46875	 => std_logic_vector(to_unsigned(17,8) ,
46876	 => std_logic_vector(to_unsigned(13,8) ,
46877	 => std_logic_vector(to_unsigned(13,8) ,
46878	 => std_logic_vector(to_unsigned(8,8) ,
46879	 => std_logic_vector(to_unsigned(13,8) ,
46880	 => std_logic_vector(to_unsigned(22,8) ,
46881	 => std_logic_vector(to_unsigned(11,8) ,
46882	 => std_logic_vector(to_unsigned(20,8) ,
46883	 => std_logic_vector(to_unsigned(43,8) ,
46884	 => std_logic_vector(to_unsigned(37,8) ,
46885	 => std_logic_vector(to_unsigned(26,8) ,
46886	 => std_logic_vector(to_unsigned(20,8) ,
46887	 => std_logic_vector(to_unsigned(21,8) ,
46888	 => std_logic_vector(to_unsigned(13,8) ,
46889	 => std_logic_vector(to_unsigned(15,8) ,
46890	 => std_logic_vector(to_unsigned(18,8) ,
46891	 => std_logic_vector(to_unsigned(16,8) ,
46892	 => std_logic_vector(to_unsigned(18,8) ,
46893	 => std_logic_vector(to_unsigned(15,8) ,
46894	 => std_logic_vector(to_unsigned(18,8) ,
46895	 => std_logic_vector(to_unsigned(39,8) ,
46896	 => std_logic_vector(to_unsigned(36,8) ,
46897	 => std_logic_vector(to_unsigned(27,8) ,
46898	 => std_logic_vector(to_unsigned(26,8) ,
46899	 => std_logic_vector(to_unsigned(25,8) ,
46900	 => std_logic_vector(to_unsigned(24,8) ,
46901	 => std_logic_vector(to_unsigned(24,8) ,
46902	 => std_logic_vector(to_unsigned(29,8) ,
46903	 => std_logic_vector(to_unsigned(38,8) ,
46904	 => std_logic_vector(to_unsigned(35,8) ,
46905	 => std_logic_vector(to_unsigned(20,8) ,
46906	 => std_logic_vector(to_unsigned(15,8) ,
46907	 => std_logic_vector(to_unsigned(16,8) ,
46908	 => std_logic_vector(to_unsigned(13,8) ,
46909	 => std_logic_vector(to_unsigned(12,8) ,
46910	 => std_logic_vector(to_unsigned(30,8) ,
46911	 => std_logic_vector(to_unsigned(69,8) ,
46912	 => std_logic_vector(to_unsigned(51,8) ,
46913	 => std_logic_vector(to_unsigned(45,8) ,
46914	 => std_logic_vector(to_unsigned(58,8) ,
46915	 => std_logic_vector(to_unsigned(69,8) ,
46916	 => std_logic_vector(to_unsigned(64,8) ,
46917	 => std_logic_vector(to_unsigned(64,8) ,
46918	 => std_logic_vector(to_unsigned(79,8) ,
46919	 => std_logic_vector(to_unsigned(78,8) ,
46920	 => std_logic_vector(to_unsigned(65,8) ,
46921	 => std_logic_vector(to_unsigned(76,8) ,
46922	 => std_logic_vector(to_unsigned(66,8) ,
46923	 => std_logic_vector(to_unsigned(45,8) ,
46924	 => std_logic_vector(to_unsigned(50,8) ,
46925	 => std_logic_vector(to_unsigned(31,8) ,
46926	 => std_logic_vector(to_unsigned(4,8) ,
46927	 => std_logic_vector(to_unsigned(4,8) ,
46928	 => std_logic_vector(to_unsigned(3,8) ,
46929	 => std_logic_vector(to_unsigned(2,8) ,
46930	 => std_logic_vector(to_unsigned(8,8) ,
46931	 => std_logic_vector(to_unsigned(47,8) ,
46932	 => std_logic_vector(to_unsigned(32,8) ,
46933	 => std_logic_vector(to_unsigned(3,8) ,
46934	 => std_logic_vector(to_unsigned(2,8) ,
46935	 => std_logic_vector(to_unsigned(2,8) ,
46936	 => std_logic_vector(to_unsigned(2,8) ,
46937	 => std_logic_vector(to_unsigned(24,8) ,
46938	 => std_logic_vector(to_unsigned(74,8) ,
46939	 => std_logic_vector(to_unsigned(90,8) ,
46940	 => std_logic_vector(to_unsigned(88,8) ,
46941	 => std_logic_vector(to_unsigned(68,8) ,
46942	 => std_logic_vector(to_unsigned(69,8) ,
46943	 => std_logic_vector(to_unsigned(71,8) ,
46944	 => std_logic_vector(to_unsigned(78,8) ,
46945	 => std_logic_vector(to_unsigned(92,8) ,
46946	 => std_logic_vector(to_unsigned(82,8) ,
46947	 => std_logic_vector(to_unsigned(73,8) ,
46948	 => std_logic_vector(to_unsigned(79,8) ,
46949	 => std_logic_vector(to_unsigned(73,8) ,
46950	 => std_logic_vector(to_unsigned(11,8) ,
46951	 => std_logic_vector(to_unsigned(4,8) ,
46952	 => std_logic_vector(to_unsigned(7,8) ,
46953	 => std_logic_vector(to_unsigned(9,8) ,
46954	 => std_logic_vector(to_unsigned(5,8) ,
46955	 => std_logic_vector(to_unsigned(4,8) ,
46956	 => std_logic_vector(to_unsigned(5,8) ,
46957	 => std_logic_vector(to_unsigned(1,8) ,
46958	 => std_logic_vector(to_unsigned(2,8) ,
46959	 => std_logic_vector(to_unsigned(4,8) ,
46960	 => std_logic_vector(to_unsigned(3,8) ,
46961	 => std_logic_vector(to_unsigned(1,8) ,
46962	 => std_logic_vector(to_unsigned(4,8) ,
46963	 => std_logic_vector(to_unsigned(70,8) ,
46964	 => std_logic_vector(to_unsigned(115,8) ,
46965	 => std_logic_vector(to_unsigned(100,8) ,
46966	 => std_logic_vector(to_unsigned(119,8) ,
46967	 => std_logic_vector(to_unsigned(109,8) ,
46968	 => std_logic_vector(to_unsigned(19,8) ,
46969	 => std_logic_vector(to_unsigned(1,8) ,
46970	 => std_logic_vector(to_unsigned(18,8) ,
46971	 => std_logic_vector(to_unsigned(136,8) ,
46972	 => std_logic_vector(to_unsigned(157,8) ,
46973	 => std_logic_vector(to_unsigned(127,8) ,
46974	 => std_logic_vector(to_unsigned(118,8) ,
46975	 => std_logic_vector(to_unsigned(142,8) ,
46976	 => std_logic_vector(to_unsigned(32,8) ,
46977	 => std_logic_vector(to_unsigned(2,8) ,
46978	 => std_logic_vector(to_unsigned(4,8) ,
46979	 => std_logic_vector(to_unsigned(4,8) ,
46980	 => std_logic_vector(to_unsigned(3,8) ,
46981	 => std_logic_vector(to_unsigned(2,8) ,
46982	 => std_logic_vector(to_unsigned(0,8) ,
46983	 => std_logic_vector(to_unsigned(15,8) ,
46984	 => std_logic_vector(to_unsigned(149,8) ,
46985	 => std_logic_vector(to_unsigned(138,8) ,
46986	 => std_logic_vector(to_unsigned(144,8) ,
46987	 => std_logic_vector(to_unsigned(177,8) ,
46988	 => std_logic_vector(to_unsigned(91,8) ,
46989	 => std_logic_vector(to_unsigned(5,8) ,
46990	 => std_logic_vector(to_unsigned(5,8) ,
46991	 => std_logic_vector(to_unsigned(2,8) ,
46992	 => std_logic_vector(to_unsigned(8,8) ,
46993	 => std_logic_vector(to_unsigned(6,8) ,
46994	 => std_logic_vector(to_unsigned(2,8) ,
46995	 => std_logic_vector(to_unsigned(1,8) ,
46996	 => std_logic_vector(to_unsigned(2,8) ,
46997	 => std_logic_vector(to_unsigned(2,8) ,
46998	 => std_logic_vector(to_unsigned(17,8) ,
46999	 => std_logic_vector(to_unsigned(92,8) ,
47000	 => std_logic_vector(to_unsigned(81,8) ,
47001	 => std_logic_vector(to_unsigned(108,8) ,
47002	 => std_logic_vector(to_unsigned(51,8) ,
47003	 => std_logic_vector(to_unsigned(1,8) ,
47004	 => std_logic_vector(to_unsigned(2,8) ,
47005	 => std_logic_vector(to_unsigned(4,8) ,
47006	 => std_logic_vector(to_unsigned(2,8) ,
47007	 => std_logic_vector(to_unsigned(2,8) ,
47008	 => std_logic_vector(to_unsigned(2,8) ,
47009	 => std_logic_vector(to_unsigned(18,8) ,
47010	 => std_logic_vector(to_unsigned(28,8) ,
47011	 => std_logic_vector(to_unsigned(22,8) ,
47012	 => std_logic_vector(to_unsigned(21,8) ,
47013	 => std_logic_vector(to_unsigned(19,8) ,
47014	 => std_logic_vector(to_unsigned(16,8) ,
47015	 => std_logic_vector(to_unsigned(8,8) ,
47016	 => std_logic_vector(to_unsigned(3,8) ,
47017	 => std_logic_vector(to_unsigned(3,8) ,
47018	 => std_logic_vector(to_unsigned(3,8) ,
47019	 => std_logic_vector(to_unsigned(3,8) ,
47020	 => std_logic_vector(to_unsigned(3,8) ,
47021	 => std_logic_vector(to_unsigned(2,8) ,
47022	 => std_logic_vector(to_unsigned(3,8) ,
47023	 => std_logic_vector(to_unsigned(2,8) ,
47024	 => std_logic_vector(to_unsigned(2,8) ,
47025	 => std_logic_vector(to_unsigned(2,8) ,
47026	 => std_logic_vector(to_unsigned(2,8) ,
47027	 => std_logic_vector(to_unsigned(3,8) ,
47028	 => std_logic_vector(to_unsigned(3,8) ,
47029	 => std_logic_vector(to_unsigned(2,8) ,
47030	 => std_logic_vector(to_unsigned(3,8) ,
47031	 => std_logic_vector(to_unsigned(5,8) ,
47032	 => std_logic_vector(to_unsigned(6,8) ,
47033	 => std_logic_vector(to_unsigned(5,8) ,
47034	 => std_logic_vector(to_unsigned(5,8) ,
47035	 => std_logic_vector(to_unsigned(6,8) ,
47036	 => std_logic_vector(to_unsigned(6,8) ,
47037	 => std_logic_vector(to_unsigned(7,8) ,
47038	 => std_logic_vector(to_unsigned(7,8) ,
47039	 => std_logic_vector(to_unsigned(7,8) ,
47040	 => std_logic_vector(to_unsigned(7,8) ,
47041	 => std_logic_vector(to_unsigned(68,8) ,
47042	 => std_logic_vector(to_unsigned(67,8) ,
47043	 => std_logic_vector(to_unsigned(62,8) ,
47044	 => std_logic_vector(to_unsigned(58,8) ,
47045	 => std_logic_vector(to_unsigned(44,8) ,
47046	 => std_logic_vector(to_unsigned(46,8) ,
47047	 => std_logic_vector(to_unsigned(49,8) ,
47048	 => std_logic_vector(to_unsigned(49,8) ,
47049	 => std_logic_vector(to_unsigned(41,8) ,
47050	 => std_logic_vector(to_unsigned(29,8) ,
47051	 => std_logic_vector(to_unsigned(30,8) ,
47052	 => std_logic_vector(to_unsigned(32,8) ,
47053	 => std_logic_vector(to_unsigned(26,8) ,
47054	 => std_logic_vector(to_unsigned(32,8) ,
47055	 => std_logic_vector(to_unsigned(69,8) ,
47056	 => std_logic_vector(to_unsigned(100,8) ,
47057	 => std_logic_vector(to_unsigned(100,8) ,
47058	 => std_logic_vector(to_unsigned(99,8) ,
47059	 => std_logic_vector(to_unsigned(99,8) ,
47060	 => std_logic_vector(to_unsigned(107,8) ,
47061	 => std_logic_vector(to_unsigned(104,8) ,
47062	 => std_logic_vector(to_unsigned(99,8) ,
47063	 => std_logic_vector(to_unsigned(99,8) ,
47064	 => std_logic_vector(to_unsigned(114,8) ,
47065	 => std_logic_vector(to_unsigned(108,8) ,
47066	 => std_logic_vector(to_unsigned(115,8) ,
47067	 => std_logic_vector(to_unsigned(124,8) ,
47068	 => std_logic_vector(to_unsigned(115,8) ,
47069	 => std_logic_vector(to_unsigned(111,8) ,
47070	 => std_logic_vector(to_unsigned(107,8) ,
47071	 => std_logic_vector(to_unsigned(125,8) ,
47072	 => std_logic_vector(to_unsigned(142,8) ,
47073	 => std_logic_vector(to_unsigned(156,8) ,
47074	 => std_logic_vector(to_unsigned(154,8) ,
47075	 => std_logic_vector(to_unsigned(149,8) ,
47076	 => std_logic_vector(to_unsigned(149,8) ,
47077	 => std_logic_vector(to_unsigned(156,8) ,
47078	 => std_logic_vector(to_unsigned(154,8) ,
47079	 => std_logic_vector(to_unsigned(161,8) ,
47080	 => std_logic_vector(to_unsigned(157,8) ,
47081	 => std_logic_vector(to_unsigned(149,8) ,
47082	 => std_logic_vector(to_unsigned(104,8) ,
47083	 => std_logic_vector(to_unsigned(66,8) ,
47084	 => std_logic_vector(to_unsigned(68,8) ,
47085	 => std_logic_vector(to_unsigned(71,8) ,
47086	 => std_logic_vector(to_unsigned(64,8) ,
47087	 => std_logic_vector(to_unsigned(67,8) ,
47088	 => std_logic_vector(to_unsigned(69,8) ,
47089	 => std_logic_vector(to_unsigned(86,8) ,
47090	 => std_logic_vector(to_unsigned(100,8) ,
47091	 => std_logic_vector(to_unsigned(84,8) ,
47092	 => std_logic_vector(to_unsigned(59,8) ,
47093	 => std_logic_vector(to_unsigned(63,8) ,
47094	 => std_logic_vector(to_unsigned(97,8) ,
47095	 => std_logic_vector(to_unsigned(96,8) ,
47096	 => std_logic_vector(to_unsigned(92,8) ,
47097	 => std_logic_vector(to_unsigned(96,8) ,
47098	 => std_logic_vector(to_unsigned(85,8) ,
47099	 => std_logic_vector(to_unsigned(80,8) ,
47100	 => std_logic_vector(to_unsigned(80,8) ,
47101	 => std_logic_vector(to_unsigned(85,8) ,
47102	 => std_logic_vector(to_unsigned(59,8) ,
47103	 => std_logic_vector(to_unsigned(55,8) ,
47104	 => std_logic_vector(to_unsigned(58,8) ,
47105	 => std_logic_vector(to_unsigned(53,8) ,
47106	 => std_logic_vector(to_unsigned(60,8) ,
47107	 => std_logic_vector(to_unsigned(64,8) ,
47108	 => std_logic_vector(to_unsigned(62,8) ,
47109	 => std_logic_vector(to_unsigned(54,8) ,
47110	 => std_logic_vector(to_unsigned(49,8) ,
47111	 => std_logic_vector(to_unsigned(53,8) ,
47112	 => std_logic_vector(to_unsigned(53,8) ,
47113	 => std_logic_vector(to_unsigned(49,8) ,
47114	 => std_logic_vector(to_unsigned(45,8) ,
47115	 => std_logic_vector(to_unsigned(46,8) ,
47116	 => std_logic_vector(to_unsigned(76,8) ,
47117	 => std_logic_vector(to_unsigned(90,8) ,
47118	 => std_logic_vector(to_unsigned(82,8) ,
47119	 => std_logic_vector(to_unsigned(87,8) ,
47120	 => std_logic_vector(to_unsigned(80,8) ,
47121	 => std_logic_vector(to_unsigned(62,8) ,
47122	 => std_logic_vector(to_unsigned(72,8) ,
47123	 => std_logic_vector(to_unsigned(68,8) ,
47124	 => std_logic_vector(to_unsigned(82,8) ,
47125	 => std_logic_vector(to_unsigned(79,8) ,
47126	 => std_logic_vector(to_unsigned(63,8) ,
47127	 => std_logic_vector(to_unsigned(62,8) ,
47128	 => std_logic_vector(to_unsigned(53,8) ,
47129	 => std_logic_vector(to_unsigned(48,8) ,
47130	 => std_logic_vector(to_unsigned(50,8) ,
47131	 => std_logic_vector(to_unsigned(44,8) ,
47132	 => std_logic_vector(to_unsigned(54,8) ,
47133	 => std_logic_vector(to_unsigned(62,8) ,
47134	 => std_logic_vector(to_unsigned(50,8) ,
47135	 => std_logic_vector(to_unsigned(50,8) ,
47136	 => std_logic_vector(to_unsigned(53,8) ,
47137	 => std_logic_vector(to_unsigned(63,8) ,
47138	 => std_logic_vector(to_unsigned(60,8) ,
47139	 => std_logic_vector(to_unsigned(55,8) ,
47140	 => std_logic_vector(to_unsigned(56,8) ,
47141	 => std_logic_vector(to_unsigned(66,8) ,
47142	 => std_logic_vector(to_unsigned(69,8) ,
47143	 => std_logic_vector(to_unsigned(72,8) ,
47144	 => std_logic_vector(to_unsigned(108,8) ,
47145	 => std_logic_vector(to_unsigned(96,8) ,
47146	 => std_logic_vector(to_unsigned(87,8) ,
47147	 => std_logic_vector(to_unsigned(93,8) ,
47148	 => std_logic_vector(to_unsigned(101,8) ,
47149	 => std_logic_vector(to_unsigned(96,8) ,
47150	 => std_logic_vector(to_unsigned(104,8) ,
47151	 => std_logic_vector(to_unsigned(122,8) ,
47152	 => std_logic_vector(to_unsigned(104,8) ,
47153	 => std_logic_vector(to_unsigned(77,8) ,
47154	 => std_logic_vector(to_unsigned(85,8) ,
47155	 => std_logic_vector(to_unsigned(88,8) ,
47156	 => std_logic_vector(to_unsigned(54,8) ,
47157	 => std_logic_vector(to_unsigned(52,8) ,
47158	 => std_logic_vector(to_unsigned(59,8) ,
47159	 => std_logic_vector(to_unsigned(56,8) ,
47160	 => std_logic_vector(to_unsigned(55,8) ,
47161	 => std_logic_vector(to_unsigned(65,8) ,
47162	 => std_logic_vector(to_unsigned(62,8) ,
47163	 => std_logic_vector(to_unsigned(51,8) ,
47164	 => std_logic_vector(to_unsigned(56,8) ,
47165	 => std_logic_vector(to_unsigned(77,8) ,
47166	 => std_logic_vector(to_unsigned(82,8) ,
47167	 => std_logic_vector(to_unsigned(91,8) ,
47168	 => std_logic_vector(to_unsigned(90,8) ,
47169	 => std_logic_vector(to_unsigned(71,8) ,
47170	 => std_logic_vector(to_unsigned(70,8) ,
47171	 => std_logic_vector(to_unsigned(92,8) ,
47172	 => std_logic_vector(to_unsigned(88,8) ,
47173	 => std_logic_vector(to_unsigned(74,8) ,
47174	 => std_logic_vector(to_unsigned(79,8) ,
47175	 => std_logic_vector(to_unsigned(72,8) ,
47176	 => std_logic_vector(to_unsigned(52,8) ,
47177	 => std_logic_vector(to_unsigned(32,8) ,
47178	 => std_logic_vector(to_unsigned(30,8) ,
47179	 => std_logic_vector(to_unsigned(38,8) ,
47180	 => std_logic_vector(to_unsigned(72,8) ,
47181	 => std_logic_vector(to_unsigned(86,8) ,
47182	 => std_logic_vector(to_unsigned(81,8) ,
47183	 => std_logic_vector(to_unsigned(57,8) ,
47184	 => std_logic_vector(to_unsigned(67,8) ,
47185	 => std_logic_vector(to_unsigned(76,8) ,
47186	 => std_logic_vector(to_unsigned(23,8) ,
47187	 => std_logic_vector(to_unsigned(8,8) ,
47188	 => std_logic_vector(to_unsigned(7,8) ,
47189	 => std_logic_vector(to_unsigned(9,8) ,
47190	 => std_logic_vector(to_unsigned(11,8) ,
47191	 => std_logic_vector(to_unsigned(14,8) ,
47192	 => std_logic_vector(to_unsigned(11,8) ,
47193	 => std_logic_vector(to_unsigned(12,8) ,
47194	 => std_logic_vector(to_unsigned(24,8) ,
47195	 => std_logic_vector(to_unsigned(23,8) ,
47196	 => std_logic_vector(to_unsigned(15,8) ,
47197	 => std_logic_vector(to_unsigned(17,8) ,
47198	 => std_logic_vector(to_unsigned(11,8) ,
47199	 => std_logic_vector(to_unsigned(10,8) ,
47200	 => std_logic_vector(to_unsigned(10,8) ,
47201	 => std_logic_vector(to_unsigned(9,8) ,
47202	 => std_logic_vector(to_unsigned(8,8) ,
47203	 => std_logic_vector(to_unsigned(8,8) ,
47204	 => std_logic_vector(to_unsigned(10,8) ,
47205	 => std_logic_vector(to_unsigned(11,8) ,
47206	 => std_logic_vector(to_unsigned(8,8) ,
47207	 => std_logic_vector(to_unsigned(17,8) ,
47208	 => std_logic_vector(to_unsigned(17,8) ,
47209	 => std_logic_vector(to_unsigned(18,8) ,
47210	 => std_logic_vector(to_unsigned(17,8) ,
47211	 => std_logic_vector(to_unsigned(23,8) ,
47212	 => std_logic_vector(to_unsigned(32,8) ,
47213	 => std_logic_vector(to_unsigned(17,8) ,
47214	 => std_logic_vector(to_unsigned(21,8) ,
47215	 => std_logic_vector(to_unsigned(54,8) ,
47216	 => std_logic_vector(to_unsigned(71,8) ,
47217	 => std_logic_vector(to_unsigned(92,8) ,
47218	 => std_logic_vector(to_unsigned(84,8) ,
47219	 => std_logic_vector(to_unsigned(74,8) ,
47220	 => std_logic_vector(to_unsigned(61,8) ,
47221	 => std_logic_vector(to_unsigned(57,8) ,
47222	 => std_logic_vector(to_unsigned(43,8) ,
47223	 => std_logic_vector(to_unsigned(37,8) ,
47224	 => std_logic_vector(to_unsigned(37,8) ,
47225	 => std_logic_vector(to_unsigned(21,8) ,
47226	 => std_logic_vector(to_unsigned(12,8) ,
47227	 => std_logic_vector(to_unsigned(15,8) ,
47228	 => std_logic_vector(to_unsigned(20,8) ,
47229	 => std_logic_vector(to_unsigned(16,8) ,
47230	 => std_logic_vector(to_unsigned(30,8) ,
47231	 => std_logic_vector(to_unsigned(61,8) ,
47232	 => std_logic_vector(to_unsigned(56,8) ,
47233	 => std_logic_vector(to_unsigned(45,8) ,
47234	 => std_logic_vector(to_unsigned(52,8) ,
47235	 => std_logic_vector(to_unsigned(52,8) ,
47236	 => std_logic_vector(to_unsigned(48,8) ,
47237	 => std_logic_vector(to_unsigned(56,8) ,
47238	 => std_logic_vector(to_unsigned(62,8) ,
47239	 => std_logic_vector(to_unsigned(52,8) ,
47240	 => std_logic_vector(to_unsigned(20,8) ,
47241	 => std_logic_vector(to_unsigned(17,8) ,
47242	 => std_logic_vector(to_unsigned(32,8) ,
47243	 => std_logic_vector(to_unsigned(44,8) ,
47244	 => std_logic_vector(to_unsigned(40,8) ,
47245	 => std_logic_vector(to_unsigned(39,8) ,
47246	 => std_logic_vector(to_unsigned(19,8) ,
47247	 => std_logic_vector(to_unsigned(6,8) ,
47248	 => std_logic_vector(to_unsigned(5,8) ,
47249	 => std_logic_vector(to_unsigned(18,8) ,
47250	 => std_logic_vector(to_unsigned(38,8) ,
47251	 => std_logic_vector(to_unsigned(44,8) ,
47252	 => std_logic_vector(to_unsigned(41,8) ,
47253	 => std_logic_vector(to_unsigned(24,8) ,
47254	 => std_logic_vector(to_unsigned(8,8) ,
47255	 => std_logic_vector(to_unsigned(6,8) ,
47256	 => std_logic_vector(to_unsigned(19,8) ,
47257	 => std_logic_vector(to_unsigned(61,8) ,
47258	 => std_logic_vector(to_unsigned(56,8) ,
47259	 => std_logic_vector(to_unsigned(69,8) ,
47260	 => std_logic_vector(to_unsigned(80,8) ,
47261	 => std_logic_vector(to_unsigned(63,8) ,
47262	 => std_logic_vector(to_unsigned(63,8) ,
47263	 => std_logic_vector(to_unsigned(66,8) ,
47264	 => std_logic_vector(to_unsigned(66,8) ,
47265	 => std_logic_vector(to_unsigned(82,8) ,
47266	 => std_logic_vector(to_unsigned(69,8) ,
47267	 => std_logic_vector(to_unsigned(59,8) ,
47268	 => std_logic_vector(to_unsigned(64,8) ,
47269	 => std_logic_vector(to_unsigned(64,8) ,
47270	 => std_logic_vector(to_unsigned(8,8) ,
47271	 => std_logic_vector(to_unsigned(1,8) ,
47272	 => std_logic_vector(to_unsigned(2,8) ,
47273	 => std_logic_vector(to_unsigned(2,8) ,
47274	 => std_logic_vector(to_unsigned(5,8) ,
47275	 => std_logic_vector(to_unsigned(40,8) ,
47276	 => std_logic_vector(to_unsigned(44,8) ,
47277	 => std_logic_vector(to_unsigned(2,8) ,
47278	 => std_logic_vector(to_unsigned(1,8) ,
47279	 => std_logic_vector(to_unsigned(1,8) ,
47280	 => std_logic_vector(to_unsigned(1,8) ,
47281	 => std_logic_vector(to_unsigned(4,8) ,
47282	 => std_logic_vector(to_unsigned(47,8) ,
47283	 => std_logic_vector(to_unsigned(112,8) ,
47284	 => std_logic_vector(to_unsigned(92,8) ,
47285	 => std_logic_vector(to_unsigned(100,8) ,
47286	 => std_logic_vector(to_unsigned(99,8) ,
47287	 => std_logic_vector(to_unsigned(107,8) ,
47288	 => std_logic_vector(to_unsigned(36,8) ,
47289	 => std_logic_vector(to_unsigned(1,8) ,
47290	 => std_logic_vector(to_unsigned(3,8) ,
47291	 => std_logic_vector(to_unsigned(88,8) ,
47292	 => std_logic_vector(to_unsigned(173,8) ,
47293	 => std_logic_vector(to_unsigned(141,8) ,
47294	 => std_logic_vector(to_unsigned(161,8) ,
47295	 => std_logic_vector(to_unsigned(130,8) ,
47296	 => std_logic_vector(to_unsigned(8,8) ,
47297	 => std_logic_vector(to_unsigned(1,8) ,
47298	 => std_logic_vector(to_unsigned(5,8) ,
47299	 => std_logic_vector(to_unsigned(6,8) ,
47300	 => std_logic_vector(to_unsigned(5,8) ,
47301	 => std_logic_vector(to_unsigned(2,8) ,
47302	 => std_logic_vector(to_unsigned(0,8) ,
47303	 => std_logic_vector(to_unsigned(21,8) ,
47304	 => std_logic_vector(to_unsigned(157,8) ,
47305	 => std_logic_vector(to_unsigned(133,8) ,
47306	 => std_logic_vector(to_unsigned(152,8) ,
47307	 => std_logic_vector(to_unsigned(179,8) ,
47308	 => std_logic_vector(to_unsigned(42,8) ,
47309	 => std_logic_vector(to_unsigned(2,8) ,
47310	 => std_logic_vector(to_unsigned(8,8) ,
47311	 => std_logic_vector(to_unsigned(3,8) ,
47312	 => std_logic_vector(to_unsigned(8,8) ,
47313	 => std_logic_vector(to_unsigned(6,8) ,
47314	 => std_logic_vector(to_unsigned(2,8) ,
47315	 => std_logic_vector(to_unsigned(1,8) ,
47316	 => std_logic_vector(to_unsigned(1,8) ,
47317	 => std_logic_vector(to_unsigned(1,8) ,
47318	 => std_logic_vector(to_unsigned(6,8) ,
47319	 => std_logic_vector(to_unsigned(52,8) ,
47320	 => std_logic_vector(to_unsigned(74,8) ,
47321	 => std_logic_vector(to_unsigned(92,8) ,
47322	 => std_logic_vector(to_unsigned(27,8) ,
47323	 => std_logic_vector(to_unsigned(0,8) ,
47324	 => std_logic_vector(to_unsigned(0,8) ,
47325	 => std_logic_vector(to_unsigned(2,8) ,
47326	 => std_logic_vector(to_unsigned(4,8) ,
47327	 => std_logic_vector(to_unsigned(2,8) ,
47328	 => std_logic_vector(to_unsigned(2,8) ,
47329	 => std_logic_vector(to_unsigned(34,8) ,
47330	 => std_logic_vector(to_unsigned(62,8) ,
47331	 => std_logic_vector(to_unsigned(88,8) ,
47332	 => std_logic_vector(to_unsigned(95,8) ,
47333	 => std_logic_vector(to_unsigned(91,8) ,
47334	 => std_logic_vector(to_unsigned(109,8) ,
47335	 => std_logic_vector(to_unsigned(56,8) ,
47336	 => std_logic_vector(to_unsigned(35,8) ,
47337	 => std_logic_vector(to_unsigned(45,8) ,
47338	 => std_logic_vector(to_unsigned(31,8) ,
47339	 => std_logic_vector(to_unsigned(15,8) ,
47340	 => std_logic_vector(to_unsigned(16,8) ,
47341	 => std_logic_vector(to_unsigned(16,8) ,
47342	 => std_logic_vector(to_unsigned(10,8) ,
47343	 => std_logic_vector(to_unsigned(11,8) ,
47344	 => std_logic_vector(to_unsigned(11,8) ,
47345	 => std_logic_vector(to_unsigned(6,8) ,
47346	 => std_logic_vector(to_unsigned(4,8) ,
47347	 => std_logic_vector(to_unsigned(4,8) ,
47348	 => std_logic_vector(to_unsigned(2,8) ,
47349	 => std_logic_vector(to_unsigned(2,8) ,
47350	 => std_logic_vector(to_unsigned(2,8) ,
47351	 => std_logic_vector(to_unsigned(1,8) ,
47352	 => std_logic_vector(to_unsigned(2,8) ,
47353	 => std_logic_vector(to_unsigned(2,8) ,
47354	 => std_logic_vector(to_unsigned(3,8) ,
47355	 => std_logic_vector(to_unsigned(2,8) ,
47356	 => std_logic_vector(to_unsigned(4,8) ,
47357	 => std_logic_vector(to_unsigned(7,8) ,
47358	 => std_logic_vector(to_unsigned(5,8) ,
47359	 => std_logic_vector(to_unsigned(4,8) ,
47360	 => std_logic_vector(to_unsigned(5,8) ,
47361	 => std_logic_vector(to_unsigned(80,8) ,
47362	 => std_logic_vector(to_unsigned(74,8) ,
47363	 => std_logic_vector(to_unsigned(56,8) ,
47364	 => std_logic_vector(to_unsigned(50,8) ,
47365	 => std_logic_vector(to_unsigned(55,8) ,
47366	 => std_logic_vector(to_unsigned(60,8) ,
47367	 => std_logic_vector(to_unsigned(51,8) ,
47368	 => std_logic_vector(to_unsigned(52,8) ,
47369	 => std_logic_vector(to_unsigned(36,8) ,
47370	 => std_logic_vector(to_unsigned(24,8) ,
47371	 => std_logic_vector(to_unsigned(28,8) ,
47372	 => std_logic_vector(to_unsigned(25,8) ,
47373	 => std_logic_vector(to_unsigned(25,8) ,
47374	 => std_logic_vector(to_unsigned(33,8) ,
47375	 => std_logic_vector(to_unsigned(69,8) ,
47376	 => std_logic_vector(to_unsigned(97,8) ,
47377	 => std_logic_vector(to_unsigned(92,8) ,
47378	 => std_logic_vector(to_unsigned(100,8) ,
47379	 => std_logic_vector(to_unsigned(97,8) ,
47380	 => std_logic_vector(to_unsigned(105,8) ,
47381	 => std_logic_vector(to_unsigned(109,8) ,
47382	 => std_logic_vector(to_unsigned(101,8) ,
47383	 => std_logic_vector(to_unsigned(100,8) ,
47384	 => std_logic_vector(to_unsigned(109,8) ,
47385	 => std_logic_vector(to_unsigned(104,8) ,
47386	 => std_logic_vector(to_unsigned(108,8) ,
47387	 => std_logic_vector(to_unsigned(112,8) ,
47388	 => std_logic_vector(to_unsigned(109,8) ,
47389	 => std_logic_vector(to_unsigned(114,8) ,
47390	 => std_logic_vector(to_unsigned(101,8) ,
47391	 => std_logic_vector(to_unsigned(108,8) ,
47392	 => std_logic_vector(to_unsigned(144,8) ,
47393	 => std_logic_vector(to_unsigned(157,8) ,
47394	 => std_logic_vector(to_unsigned(154,8) ,
47395	 => std_logic_vector(to_unsigned(151,8) ,
47396	 => std_logic_vector(to_unsigned(151,8) ,
47397	 => std_logic_vector(to_unsigned(151,8) ,
47398	 => std_logic_vector(to_unsigned(156,8) ,
47399	 => std_logic_vector(to_unsigned(154,8) ,
47400	 => std_logic_vector(to_unsigned(159,8) ,
47401	 => std_logic_vector(to_unsigned(144,8) ,
47402	 => std_logic_vector(to_unsigned(90,8) ,
47403	 => std_logic_vector(to_unsigned(81,8) ,
47404	 => std_logic_vector(to_unsigned(82,8) ,
47405	 => std_logic_vector(to_unsigned(71,8) ,
47406	 => std_logic_vector(to_unsigned(65,8) ,
47407	 => std_logic_vector(to_unsigned(90,8) ,
47408	 => std_logic_vector(to_unsigned(80,8) ,
47409	 => std_logic_vector(to_unsigned(71,8) ,
47410	 => std_logic_vector(to_unsigned(80,8) ,
47411	 => std_logic_vector(to_unsigned(80,8) ,
47412	 => std_logic_vector(to_unsigned(63,8) ,
47413	 => std_logic_vector(to_unsigned(59,8) ,
47414	 => std_logic_vector(to_unsigned(70,8) ,
47415	 => std_logic_vector(to_unsigned(77,8) ,
47416	 => std_logic_vector(to_unsigned(85,8) ,
47417	 => std_logic_vector(to_unsigned(92,8) ,
47418	 => std_logic_vector(to_unsigned(84,8) ,
47419	 => std_logic_vector(to_unsigned(74,8) ,
47420	 => std_logic_vector(to_unsigned(63,8) ,
47421	 => std_logic_vector(to_unsigned(77,8) ,
47422	 => std_logic_vector(to_unsigned(65,8) ,
47423	 => std_logic_vector(to_unsigned(51,8) ,
47424	 => std_logic_vector(to_unsigned(51,8) ,
47425	 => std_logic_vector(to_unsigned(46,8) ,
47426	 => std_logic_vector(to_unsigned(58,8) ,
47427	 => std_logic_vector(to_unsigned(77,8) ,
47428	 => std_logic_vector(to_unsigned(64,8) ,
47429	 => std_logic_vector(to_unsigned(55,8) ,
47430	 => std_logic_vector(to_unsigned(52,8) ,
47431	 => std_logic_vector(to_unsigned(49,8) ,
47432	 => std_logic_vector(to_unsigned(48,8) ,
47433	 => std_logic_vector(to_unsigned(59,8) ,
47434	 => std_logic_vector(to_unsigned(54,8) ,
47435	 => std_logic_vector(to_unsigned(44,8) ,
47436	 => std_logic_vector(to_unsigned(74,8) ,
47437	 => std_logic_vector(to_unsigned(97,8) ,
47438	 => std_logic_vector(to_unsigned(78,8) ,
47439	 => std_logic_vector(to_unsigned(79,8) ,
47440	 => std_logic_vector(to_unsigned(88,8) ,
47441	 => std_logic_vector(to_unsigned(74,8) ,
47442	 => std_logic_vector(to_unsigned(76,8) ,
47443	 => std_logic_vector(to_unsigned(80,8) ,
47444	 => std_logic_vector(to_unsigned(66,8) ,
47445	 => std_logic_vector(to_unsigned(71,8) ,
47446	 => std_logic_vector(to_unsigned(68,8) ,
47447	 => std_logic_vector(to_unsigned(61,8) ,
47448	 => std_logic_vector(to_unsigned(57,8) ,
47449	 => std_logic_vector(to_unsigned(51,8) ,
47450	 => std_logic_vector(to_unsigned(42,8) ,
47451	 => std_logic_vector(to_unsigned(42,8) ,
47452	 => std_logic_vector(to_unsigned(51,8) ,
47453	 => std_logic_vector(to_unsigned(55,8) ,
47454	 => std_logic_vector(to_unsigned(57,8) ,
47455	 => std_logic_vector(to_unsigned(73,8) ,
47456	 => std_logic_vector(to_unsigned(67,8) ,
47457	 => std_logic_vector(to_unsigned(74,8) ,
47458	 => std_logic_vector(to_unsigned(68,8) ,
47459	 => std_logic_vector(to_unsigned(60,8) ,
47460	 => std_logic_vector(to_unsigned(50,8) ,
47461	 => std_logic_vector(to_unsigned(61,8) ,
47462	 => std_logic_vector(to_unsigned(58,8) ,
47463	 => std_logic_vector(to_unsigned(67,8) ,
47464	 => std_logic_vector(to_unsigned(100,8) ,
47465	 => std_logic_vector(to_unsigned(85,8) ,
47466	 => std_logic_vector(to_unsigned(77,8) ,
47467	 => std_logic_vector(to_unsigned(76,8) ,
47468	 => std_logic_vector(to_unsigned(84,8) ,
47469	 => std_logic_vector(to_unsigned(74,8) ,
47470	 => std_logic_vector(to_unsigned(96,8) ,
47471	 => std_logic_vector(to_unsigned(118,8) ,
47472	 => std_logic_vector(to_unsigned(79,8) ,
47473	 => std_logic_vector(to_unsigned(71,8) ,
47474	 => std_logic_vector(to_unsigned(88,8) ,
47475	 => std_logic_vector(to_unsigned(88,8) ,
47476	 => std_logic_vector(to_unsigned(58,8) ,
47477	 => std_logic_vector(to_unsigned(60,8) ,
47478	 => std_logic_vector(to_unsigned(55,8) ,
47479	 => std_logic_vector(to_unsigned(51,8) ,
47480	 => std_logic_vector(to_unsigned(52,8) ,
47481	 => std_logic_vector(to_unsigned(44,8) ,
47482	 => std_logic_vector(to_unsigned(51,8) ,
47483	 => std_logic_vector(to_unsigned(48,8) ,
47484	 => std_logic_vector(to_unsigned(46,8) ,
47485	 => std_logic_vector(to_unsigned(73,8) ,
47486	 => std_logic_vector(to_unsigned(81,8) ,
47487	 => std_logic_vector(to_unsigned(82,8) ,
47488	 => std_logic_vector(to_unsigned(91,8) ,
47489	 => std_logic_vector(to_unsigned(74,8) ,
47490	 => std_logic_vector(to_unsigned(66,8) ,
47491	 => std_logic_vector(to_unsigned(77,8) ,
47492	 => std_logic_vector(to_unsigned(88,8) ,
47493	 => std_logic_vector(to_unsigned(74,8) ,
47494	 => std_logic_vector(to_unsigned(80,8) ,
47495	 => std_logic_vector(to_unsigned(64,8) ,
47496	 => std_logic_vector(to_unsigned(40,8) ,
47497	 => std_logic_vector(to_unsigned(29,8) ,
47498	 => std_logic_vector(to_unsigned(35,8) ,
47499	 => std_logic_vector(to_unsigned(46,8) ,
47500	 => std_logic_vector(to_unsigned(52,8) ,
47501	 => std_logic_vector(to_unsigned(82,8) ,
47502	 => std_logic_vector(to_unsigned(107,8) ,
47503	 => std_logic_vector(to_unsigned(73,8) ,
47504	 => std_logic_vector(to_unsigned(71,8) ,
47505	 => std_logic_vector(to_unsigned(86,8) ,
47506	 => std_logic_vector(to_unsigned(88,8) ,
47507	 => std_logic_vector(to_unsigned(30,8) ,
47508	 => std_logic_vector(to_unsigned(14,8) ,
47509	 => std_logic_vector(to_unsigned(46,8) ,
47510	 => std_logic_vector(to_unsigned(25,8) ,
47511	 => std_logic_vector(to_unsigned(22,8) ,
47512	 => std_logic_vector(to_unsigned(37,8) ,
47513	 => std_logic_vector(to_unsigned(32,8) ,
47514	 => std_logic_vector(to_unsigned(33,8) ,
47515	 => std_logic_vector(to_unsigned(29,8) ,
47516	 => std_logic_vector(to_unsigned(34,8) ,
47517	 => std_logic_vector(to_unsigned(33,8) ,
47518	 => std_logic_vector(to_unsigned(29,8) ,
47519	 => std_logic_vector(to_unsigned(32,8) ,
47520	 => std_logic_vector(to_unsigned(24,8) ,
47521	 => std_logic_vector(to_unsigned(22,8) ,
47522	 => std_logic_vector(to_unsigned(32,8) ,
47523	 => std_logic_vector(to_unsigned(35,8) ,
47524	 => std_logic_vector(to_unsigned(32,8) ,
47525	 => std_logic_vector(to_unsigned(25,8) ,
47526	 => std_logic_vector(to_unsigned(12,8) ,
47527	 => std_logic_vector(to_unsigned(27,8) ,
47528	 => std_logic_vector(to_unsigned(21,8) ,
47529	 => std_logic_vector(to_unsigned(14,8) ,
47530	 => std_logic_vector(to_unsigned(12,8) ,
47531	 => std_logic_vector(to_unsigned(15,8) ,
47532	 => std_logic_vector(to_unsigned(12,8) ,
47533	 => std_logic_vector(to_unsigned(9,8) ,
47534	 => std_logic_vector(to_unsigned(26,8) ,
47535	 => std_logic_vector(to_unsigned(52,8) ,
47536	 => std_logic_vector(to_unsigned(73,8) ,
47537	 => std_logic_vector(to_unsigned(82,8) ,
47538	 => std_logic_vector(to_unsigned(97,8) ,
47539	 => std_logic_vector(to_unsigned(97,8) ,
47540	 => std_logic_vector(to_unsigned(54,8) ,
47541	 => std_logic_vector(to_unsigned(81,8) ,
47542	 => std_logic_vector(to_unsigned(96,8) ,
47543	 => std_logic_vector(to_unsigned(63,8) ,
47544	 => std_logic_vector(to_unsigned(53,8) ,
47545	 => std_logic_vector(to_unsigned(43,8) ,
47546	 => std_logic_vector(to_unsigned(35,8) ,
47547	 => std_logic_vector(to_unsigned(30,8) ,
47548	 => std_logic_vector(to_unsigned(24,8) ,
47549	 => std_logic_vector(to_unsigned(12,8) ,
47550	 => std_logic_vector(to_unsigned(25,8) ,
47551	 => std_logic_vector(to_unsigned(50,8) ,
47552	 => std_logic_vector(to_unsigned(35,8) ,
47553	 => std_logic_vector(to_unsigned(35,8) ,
47554	 => std_logic_vector(to_unsigned(47,8) ,
47555	 => std_logic_vector(to_unsigned(52,8) ,
47556	 => std_logic_vector(to_unsigned(67,8) ,
47557	 => std_logic_vector(to_unsigned(71,8) ,
47558	 => std_logic_vector(to_unsigned(60,8) ,
47559	 => std_logic_vector(to_unsigned(61,8) ,
47560	 => std_logic_vector(to_unsigned(32,8) ,
47561	 => std_logic_vector(to_unsigned(27,8) ,
47562	 => std_logic_vector(to_unsigned(35,8) ,
47563	 => std_logic_vector(to_unsigned(37,8) ,
47564	 => std_logic_vector(to_unsigned(34,8) ,
47565	 => std_logic_vector(to_unsigned(37,8) ,
47566	 => std_logic_vector(to_unsigned(40,8) ,
47567	 => std_logic_vector(to_unsigned(41,8) ,
47568	 => std_logic_vector(to_unsigned(48,8) ,
47569	 => std_logic_vector(to_unsigned(41,8) ,
47570	 => std_logic_vector(to_unsigned(37,8) ,
47571	 => std_logic_vector(to_unsigned(39,8) ,
47572	 => std_logic_vector(to_unsigned(35,8) ,
47573	 => std_logic_vector(to_unsigned(36,8) ,
47574	 => std_logic_vector(to_unsigned(36,8) ,
47575	 => std_logic_vector(to_unsigned(41,8) ,
47576	 => std_logic_vector(to_unsigned(60,8) ,
47577	 => std_logic_vector(to_unsigned(51,8) ,
47578	 => std_logic_vector(to_unsigned(46,8) ,
47579	 => std_logic_vector(to_unsigned(69,8) ,
47580	 => std_logic_vector(to_unsigned(76,8) ,
47581	 => std_logic_vector(to_unsigned(81,8) ,
47582	 => std_logic_vector(to_unsigned(74,8) ,
47583	 => std_logic_vector(to_unsigned(58,8) ,
47584	 => std_logic_vector(to_unsigned(51,8) ,
47585	 => std_logic_vector(to_unsigned(61,8) ,
47586	 => std_logic_vector(to_unsigned(53,8) ,
47587	 => std_logic_vector(to_unsigned(55,8) ,
47588	 => std_logic_vector(to_unsigned(59,8) ,
47589	 => std_logic_vector(to_unsigned(57,8) ,
47590	 => std_logic_vector(to_unsigned(43,8) ,
47591	 => std_logic_vector(to_unsigned(19,8) ,
47592	 => std_logic_vector(to_unsigned(12,8) ,
47593	 => std_logic_vector(to_unsigned(24,8) ,
47594	 => std_logic_vector(to_unsigned(67,8) ,
47595	 => std_logic_vector(to_unsigned(73,8) ,
47596	 => std_logic_vector(to_unsigned(65,8) ,
47597	 => std_logic_vector(to_unsigned(33,8) ,
47598	 => std_logic_vector(to_unsigned(13,8) ,
47599	 => std_logic_vector(to_unsigned(6,8) ,
47600	 => std_logic_vector(to_unsigned(11,8) ,
47601	 => std_logic_vector(to_unsigned(47,8) ,
47602	 => std_logic_vector(to_unsigned(79,8) ,
47603	 => std_logic_vector(to_unsigned(87,8) ,
47604	 => std_logic_vector(to_unsigned(97,8) ,
47605	 => std_logic_vector(to_unsigned(95,8) ,
47606	 => std_logic_vector(to_unsigned(74,8) ,
47607	 => std_logic_vector(to_unsigned(82,8) ,
47608	 => std_logic_vector(to_unsigned(61,8) ,
47609	 => std_logic_vector(to_unsigned(4,8) ,
47610	 => std_logic_vector(to_unsigned(2,8) ,
47611	 => std_logic_vector(to_unsigned(29,8) ,
47612	 => std_logic_vector(to_unsigned(125,8) ,
47613	 => std_logic_vector(to_unsigned(111,8) ,
47614	 => std_logic_vector(to_unsigned(138,8) ,
47615	 => std_logic_vector(to_unsigned(81,8) ,
47616	 => std_logic_vector(to_unsigned(2,8) ,
47617	 => std_logic_vector(to_unsigned(2,8) ,
47618	 => std_logic_vector(to_unsigned(5,8) ,
47619	 => std_logic_vector(to_unsigned(6,8) ,
47620	 => std_logic_vector(to_unsigned(6,8) ,
47621	 => std_logic_vector(to_unsigned(2,8) ,
47622	 => std_logic_vector(to_unsigned(1,8) ,
47623	 => std_logic_vector(to_unsigned(61,8) ,
47624	 => std_logic_vector(to_unsigned(188,8) ,
47625	 => std_logic_vector(to_unsigned(151,8) ,
47626	 => std_logic_vector(to_unsigned(170,8) ,
47627	 => std_logic_vector(to_unsigned(151,8) ,
47628	 => std_logic_vector(to_unsigned(14,8) ,
47629	 => std_logic_vector(to_unsigned(2,8) ,
47630	 => std_logic_vector(to_unsigned(10,8) ,
47631	 => std_logic_vector(to_unsigned(8,8) ,
47632	 => std_logic_vector(to_unsigned(9,8) ,
47633	 => std_logic_vector(to_unsigned(5,8) ,
47634	 => std_logic_vector(to_unsigned(2,8) ,
47635	 => std_logic_vector(to_unsigned(1,8) ,
47636	 => std_logic_vector(to_unsigned(0,8) ,
47637	 => std_logic_vector(to_unsigned(1,8) ,
47638	 => std_logic_vector(to_unsigned(2,8) ,
47639	 => std_logic_vector(to_unsigned(35,8) ,
47640	 => std_logic_vector(to_unsigned(81,8) ,
47641	 => std_logic_vector(to_unsigned(77,8) ,
47642	 => std_logic_vector(to_unsigned(9,8) ,
47643	 => std_logic_vector(to_unsigned(1,8) ,
47644	 => std_logic_vector(to_unsigned(1,8) ,
47645	 => std_logic_vector(to_unsigned(3,8) ,
47646	 => std_logic_vector(to_unsigned(7,8) ,
47647	 => std_logic_vector(to_unsigned(3,8) ,
47648	 => std_logic_vector(to_unsigned(3,8) ,
47649	 => std_logic_vector(to_unsigned(37,8) ,
47650	 => std_logic_vector(to_unsigned(64,8) ,
47651	 => std_logic_vector(to_unsigned(64,8) ,
47652	 => std_logic_vector(to_unsigned(70,8) ,
47653	 => std_logic_vector(to_unsigned(86,8) ,
47654	 => std_logic_vector(to_unsigned(95,8) ,
47655	 => std_logic_vector(to_unsigned(49,8) ,
47656	 => std_logic_vector(to_unsigned(41,8) ,
47657	 => std_logic_vector(to_unsigned(73,8) ,
47658	 => std_logic_vector(to_unsigned(65,8) ,
47659	 => std_logic_vector(to_unsigned(51,8) ,
47660	 => std_logic_vector(to_unsigned(55,8) ,
47661	 => std_logic_vector(to_unsigned(51,8) ,
47662	 => std_logic_vector(to_unsigned(34,8) ,
47663	 => std_logic_vector(to_unsigned(46,8) ,
47664	 => std_logic_vector(to_unsigned(56,8) ,
47665	 => std_logic_vector(to_unsigned(41,8) ,
47666	 => std_logic_vector(to_unsigned(27,8) ,
47667	 => std_logic_vector(to_unsigned(27,8) ,
47668	 => std_logic_vector(to_unsigned(40,8) ,
47669	 => std_logic_vector(to_unsigned(26,8) ,
47670	 => std_logic_vector(to_unsigned(25,8) ,
47671	 => std_logic_vector(to_unsigned(18,8) ,
47672	 => std_logic_vector(to_unsigned(9,8) ,
47673	 => std_logic_vector(to_unsigned(10,8) ,
47674	 => std_logic_vector(to_unsigned(6,8) ,
47675	 => std_logic_vector(to_unsigned(4,8) ,
47676	 => std_logic_vector(to_unsigned(4,8) ,
47677	 => std_logic_vector(to_unsigned(3,8) ,
47678	 => std_logic_vector(to_unsigned(2,8) ,
47679	 => std_logic_vector(to_unsigned(2,8) ,
47680	 => std_logic_vector(to_unsigned(2,8) ,
47681	 => std_logic_vector(to_unsigned(82,8) ,
47682	 => std_logic_vector(to_unsigned(78,8) ,
47683	 => std_logic_vector(to_unsigned(78,8) ,
47684	 => std_logic_vector(to_unsigned(77,8) ,
47685	 => std_logic_vector(to_unsigned(68,8) ,
47686	 => std_logic_vector(to_unsigned(65,8) ,
47687	 => std_logic_vector(to_unsigned(55,8) ,
47688	 => std_logic_vector(to_unsigned(57,8) ,
47689	 => std_logic_vector(to_unsigned(41,8) ,
47690	 => std_logic_vector(to_unsigned(29,8) ,
47691	 => std_logic_vector(to_unsigned(25,8) ,
47692	 => std_logic_vector(to_unsigned(21,8) ,
47693	 => std_logic_vector(to_unsigned(24,8) ,
47694	 => std_logic_vector(to_unsigned(29,8) ,
47695	 => std_logic_vector(to_unsigned(61,8) ,
47696	 => std_logic_vector(to_unsigned(112,8) ,
47697	 => std_logic_vector(to_unsigned(100,8) ,
47698	 => std_logic_vector(to_unsigned(101,8) ,
47699	 => std_logic_vector(to_unsigned(101,8) ,
47700	 => std_logic_vector(to_unsigned(100,8) ,
47701	 => std_logic_vector(to_unsigned(100,8) ,
47702	 => std_logic_vector(to_unsigned(103,8) ,
47703	 => std_logic_vector(to_unsigned(105,8) ,
47704	 => std_logic_vector(to_unsigned(107,8) ,
47705	 => std_logic_vector(to_unsigned(90,8) ,
47706	 => std_logic_vector(to_unsigned(105,8) ,
47707	 => std_logic_vector(to_unsigned(105,8) ,
47708	 => std_logic_vector(to_unsigned(101,8) ,
47709	 => std_logic_vector(to_unsigned(114,8) ,
47710	 => std_logic_vector(to_unsigned(105,8) ,
47711	 => std_logic_vector(to_unsigned(105,8) ,
47712	 => std_logic_vector(to_unsigned(134,8) ,
47713	 => std_logic_vector(to_unsigned(146,8) ,
47714	 => std_logic_vector(to_unsigned(152,8) ,
47715	 => std_logic_vector(to_unsigned(151,8) ,
47716	 => std_logic_vector(to_unsigned(154,8) ,
47717	 => std_logic_vector(to_unsigned(156,8) ,
47718	 => std_logic_vector(to_unsigned(154,8) ,
47719	 => std_logic_vector(to_unsigned(151,8) ,
47720	 => std_logic_vector(to_unsigned(154,8) ,
47721	 => std_logic_vector(to_unsigned(138,8) ,
47722	 => std_logic_vector(to_unsigned(91,8) ,
47723	 => std_logic_vector(to_unsigned(122,8) ,
47724	 => std_logic_vector(to_unsigned(112,8) ,
47725	 => std_logic_vector(to_unsigned(82,8) ,
47726	 => std_logic_vector(to_unsigned(78,8) ,
47727	 => std_logic_vector(to_unsigned(84,8) ,
47728	 => std_logic_vector(to_unsigned(73,8) ,
47729	 => std_logic_vector(to_unsigned(45,8) ,
47730	 => std_logic_vector(to_unsigned(48,8) ,
47731	 => std_logic_vector(to_unsigned(82,8) ,
47732	 => std_logic_vector(to_unsigned(72,8) ,
47733	 => std_logic_vector(to_unsigned(56,8) ,
47734	 => std_logic_vector(to_unsigned(64,8) ,
47735	 => std_logic_vector(to_unsigned(74,8) ,
47736	 => std_logic_vector(to_unsigned(69,8) ,
47737	 => std_logic_vector(to_unsigned(63,8) ,
47738	 => std_logic_vector(to_unsigned(80,8) ,
47739	 => std_logic_vector(to_unsigned(86,8) ,
47740	 => std_logic_vector(to_unsigned(77,8) ,
47741	 => std_logic_vector(to_unsigned(88,8) ,
47742	 => std_logic_vector(to_unsigned(87,8) ,
47743	 => std_logic_vector(to_unsigned(78,8) ,
47744	 => std_logic_vector(to_unsigned(74,8) ,
47745	 => std_logic_vector(to_unsigned(69,8) ,
47746	 => std_logic_vector(to_unsigned(65,8) ,
47747	 => std_logic_vector(to_unsigned(70,8) ,
47748	 => std_logic_vector(to_unsigned(63,8) ,
47749	 => std_logic_vector(to_unsigned(45,8) ,
47750	 => std_logic_vector(to_unsigned(43,8) ,
47751	 => std_logic_vector(to_unsigned(45,8) ,
47752	 => std_logic_vector(to_unsigned(47,8) ,
47753	 => std_logic_vector(to_unsigned(51,8) ,
47754	 => std_logic_vector(to_unsigned(52,8) ,
47755	 => std_logic_vector(to_unsigned(44,8) ,
47756	 => std_logic_vector(to_unsigned(70,8) ,
47757	 => std_logic_vector(to_unsigned(91,8) ,
47758	 => std_logic_vector(to_unsigned(70,8) ,
47759	 => std_logic_vector(to_unsigned(73,8) ,
47760	 => std_logic_vector(to_unsigned(84,8) ,
47761	 => std_logic_vector(to_unsigned(72,8) ,
47762	 => std_logic_vector(to_unsigned(60,8) ,
47763	 => std_logic_vector(to_unsigned(69,8) ,
47764	 => std_logic_vector(to_unsigned(73,8) ,
47765	 => std_logic_vector(to_unsigned(64,8) ,
47766	 => std_logic_vector(to_unsigned(53,8) ,
47767	 => std_logic_vector(to_unsigned(58,8) ,
47768	 => std_logic_vector(to_unsigned(56,8) ,
47769	 => std_logic_vector(to_unsigned(42,8) ,
47770	 => std_logic_vector(to_unsigned(39,8) ,
47771	 => std_logic_vector(to_unsigned(46,8) ,
47772	 => std_logic_vector(to_unsigned(50,8) ,
47773	 => std_logic_vector(to_unsigned(49,8) ,
47774	 => std_logic_vector(to_unsigned(54,8) ,
47775	 => std_logic_vector(to_unsigned(72,8) ,
47776	 => std_logic_vector(to_unsigned(72,8) ,
47777	 => std_logic_vector(to_unsigned(90,8) ,
47778	 => std_logic_vector(to_unsigned(90,8) ,
47779	 => std_logic_vector(to_unsigned(92,8) ,
47780	 => std_logic_vector(to_unsigned(59,8) ,
47781	 => std_logic_vector(to_unsigned(59,8) ,
47782	 => std_logic_vector(to_unsigned(61,8) ,
47783	 => std_logic_vector(to_unsigned(64,8) ,
47784	 => std_logic_vector(to_unsigned(95,8) ,
47785	 => std_logic_vector(to_unsigned(84,8) ,
47786	 => std_logic_vector(to_unsigned(81,8) ,
47787	 => std_logic_vector(to_unsigned(78,8) ,
47788	 => std_logic_vector(to_unsigned(73,8) ,
47789	 => std_logic_vector(to_unsigned(68,8) ,
47790	 => std_logic_vector(to_unsigned(82,8) ,
47791	 => std_logic_vector(to_unsigned(107,8) ,
47792	 => std_logic_vector(to_unsigned(84,8) ,
47793	 => std_logic_vector(to_unsigned(72,8) ,
47794	 => std_logic_vector(to_unsigned(79,8) ,
47795	 => std_logic_vector(to_unsigned(96,8) ,
47796	 => std_logic_vector(to_unsigned(73,8) ,
47797	 => std_logic_vector(to_unsigned(68,8) ,
47798	 => std_logic_vector(to_unsigned(66,8) ,
47799	 => std_logic_vector(to_unsigned(53,8) ,
47800	 => std_logic_vector(to_unsigned(47,8) ,
47801	 => std_logic_vector(to_unsigned(46,8) ,
47802	 => std_logic_vector(to_unsigned(42,8) ,
47803	 => std_logic_vector(to_unsigned(41,8) ,
47804	 => std_logic_vector(to_unsigned(47,8) ,
47805	 => std_logic_vector(to_unsigned(74,8) ,
47806	 => std_logic_vector(to_unsigned(73,8) ,
47807	 => std_logic_vector(to_unsigned(79,8) ,
47808	 => std_logic_vector(to_unsigned(76,8) ,
47809	 => std_logic_vector(to_unsigned(67,8) ,
47810	 => std_logic_vector(to_unsigned(71,8) ,
47811	 => std_logic_vector(to_unsigned(90,8) ,
47812	 => std_logic_vector(to_unsigned(81,8) ,
47813	 => std_logic_vector(to_unsigned(57,8) ,
47814	 => std_logic_vector(to_unsigned(67,8) ,
47815	 => std_logic_vector(to_unsigned(61,8) ,
47816	 => std_logic_vector(to_unsigned(37,8) ,
47817	 => std_logic_vector(to_unsigned(27,8) ,
47818	 => std_logic_vector(to_unsigned(27,8) ,
47819	 => std_logic_vector(to_unsigned(33,8) ,
47820	 => std_logic_vector(to_unsigned(61,8) ,
47821	 => std_logic_vector(to_unsigned(82,8) ,
47822	 => std_logic_vector(to_unsigned(101,8) ,
47823	 => std_logic_vector(to_unsigned(104,8) ,
47824	 => std_logic_vector(to_unsigned(101,8) ,
47825	 => std_logic_vector(to_unsigned(108,8) ,
47826	 => std_logic_vector(to_unsigned(136,8) ,
47827	 => std_logic_vector(to_unsigned(84,8) ,
47828	 => std_logic_vector(to_unsigned(88,8) ,
47829	 => std_logic_vector(to_unsigned(130,8) ,
47830	 => std_logic_vector(to_unsigned(87,8) ,
47831	 => std_logic_vector(to_unsigned(73,8) ,
47832	 => std_logic_vector(to_unsigned(74,8) ,
47833	 => std_logic_vector(to_unsigned(25,8) ,
47834	 => std_logic_vector(to_unsigned(24,8) ,
47835	 => std_logic_vector(to_unsigned(48,8) ,
47836	 => std_logic_vector(to_unsigned(48,8) ,
47837	 => std_logic_vector(to_unsigned(55,8) ,
47838	 => std_logic_vector(to_unsigned(53,8) ,
47839	 => std_logic_vector(to_unsigned(45,8) ,
47840	 => std_logic_vector(to_unsigned(52,8) ,
47841	 => std_logic_vector(to_unsigned(72,8) ,
47842	 => std_logic_vector(to_unsigned(96,8) ,
47843	 => std_logic_vector(to_unsigned(92,8) ,
47844	 => std_logic_vector(to_unsigned(95,8) ,
47845	 => std_logic_vector(to_unsigned(80,8) ,
47846	 => std_logic_vector(to_unsigned(34,8) ,
47847	 => std_logic_vector(to_unsigned(30,8) ,
47848	 => std_logic_vector(to_unsigned(32,8) ,
47849	 => std_logic_vector(to_unsigned(28,8) ,
47850	 => std_logic_vector(to_unsigned(20,8) ,
47851	 => std_logic_vector(to_unsigned(24,8) ,
47852	 => std_logic_vector(to_unsigned(16,8) ,
47853	 => std_logic_vector(to_unsigned(10,8) ,
47854	 => std_logic_vector(to_unsigned(33,8) ,
47855	 => std_logic_vector(to_unsigned(58,8) ,
47856	 => std_logic_vector(to_unsigned(62,8) ,
47857	 => std_logic_vector(to_unsigned(43,8) ,
47858	 => std_logic_vector(to_unsigned(48,8) ,
47859	 => std_logic_vector(to_unsigned(43,8) ,
47860	 => std_logic_vector(to_unsigned(35,8) ,
47861	 => std_logic_vector(to_unsigned(46,8) ,
47862	 => std_logic_vector(to_unsigned(55,8) ,
47863	 => std_logic_vector(to_unsigned(45,8) ,
47864	 => std_logic_vector(to_unsigned(50,8) ,
47865	 => std_logic_vector(to_unsigned(99,8) ,
47866	 => std_logic_vector(to_unsigned(90,8) ,
47867	 => std_logic_vector(to_unsigned(27,8) ,
47868	 => std_logic_vector(to_unsigned(18,8) ,
47869	 => std_logic_vector(to_unsigned(9,8) ,
47870	 => std_logic_vector(to_unsigned(25,8) ,
47871	 => std_logic_vector(to_unsigned(45,8) ,
47872	 => std_logic_vector(to_unsigned(24,8) ,
47873	 => std_logic_vector(to_unsigned(25,8) ,
47874	 => std_logic_vector(to_unsigned(38,8) ,
47875	 => std_logic_vector(to_unsigned(35,8) ,
47876	 => std_logic_vector(to_unsigned(35,8) ,
47877	 => std_logic_vector(to_unsigned(51,8) ,
47878	 => std_logic_vector(to_unsigned(68,8) ,
47879	 => std_logic_vector(to_unsigned(56,8) ,
47880	 => std_logic_vector(to_unsigned(37,8) ,
47881	 => std_logic_vector(to_unsigned(33,8) ,
47882	 => std_logic_vector(to_unsigned(32,8) ,
47883	 => std_logic_vector(to_unsigned(30,8) ,
47884	 => std_logic_vector(to_unsigned(32,8) ,
47885	 => std_logic_vector(to_unsigned(33,8) ,
47886	 => std_logic_vector(to_unsigned(37,8) ,
47887	 => std_logic_vector(to_unsigned(52,8) ,
47888	 => std_logic_vector(to_unsigned(62,8) ,
47889	 => std_logic_vector(to_unsigned(35,8) ,
47890	 => std_logic_vector(to_unsigned(31,8) ,
47891	 => std_logic_vector(to_unsigned(34,8) ,
47892	 => std_logic_vector(to_unsigned(34,8) ,
47893	 => std_logic_vector(to_unsigned(33,8) ,
47894	 => std_logic_vector(to_unsigned(29,8) ,
47895	 => std_logic_vector(to_unsigned(37,8) ,
47896	 => std_logic_vector(to_unsigned(52,8) ,
47897	 => std_logic_vector(to_unsigned(45,8) ,
47898	 => std_logic_vector(to_unsigned(54,8) ,
47899	 => std_logic_vector(to_unsigned(97,8) ,
47900	 => std_logic_vector(to_unsigned(81,8) ,
47901	 => std_logic_vector(to_unsigned(81,8) ,
47902	 => std_logic_vector(to_unsigned(73,8) ,
47903	 => std_logic_vector(to_unsigned(51,8) ,
47904	 => std_logic_vector(to_unsigned(52,8) ,
47905	 => std_logic_vector(to_unsigned(55,8) ,
47906	 => std_logic_vector(to_unsigned(52,8) ,
47907	 => std_logic_vector(to_unsigned(52,8) ,
47908	 => std_logic_vector(to_unsigned(56,8) ,
47909	 => std_logic_vector(to_unsigned(54,8) ,
47910	 => std_logic_vector(to_unsigned(69,8) ,
47911	 => std_logic_vector(to_unsigned(79,8) ,
47912	 => std_logic_vector(to_unsigned(76,8) ,
47913	 => std_logic_vector(to_unsigned(79,8) ,
47914	 => std_logic_vector(to_unsigned(74,8) ,
47915	 => std_logic_vector(to_unsigned(54,8) ,
47916	 => std_logic_vector(to_unsigned(49,8) ,
47917	 => std_logic_vector(to_unsigned(64,8) ,
47918	 => std_logic_vector(to_unsigned(63,8) ,
47919	 => std_logic_vector(to_unsigned(57,8) ,
47920	 => std_logic_vector(to_unsigned(71,8) ,
47921	 => std_logic_vector(to_unsigned(81,8) ,
47922	 => std_logic_vector(to_unsigned(74,8) ,
47923	 => std_logic_vector(to_unsigned(96,8) ,
47924	 => std_logic_vector(to_unsigned(103,8) ,
47925	 => std_logic_vector(to_unsigned(69,8) ,
47926	 => std_logic_vector(to_unsigned(63,8) ,
47927	 => std_logic_vector(to_unsigned(57,8) ,
47928	 => std_logic_vector(to_unsigned(52,8) ,
47929	 => std_logic_vector(to_unsigned(7,8) ,
47930	 => std_logic_vector(to_unsigned(1,8) ,
47931	 => std_logic_vector(to_unsigned(8,8) ,
47932	 => std_logic_vector(to_unsigned(103,8) ,
47933	 => std_logic_vector(to_unsigned(99,8) ,
47934	 => std_logic_vector(to_unsigned(121,8) ,
47935	 => std_logic_vector(to_unsigned(66,8) ,
47936	 => std_logic_vector(to_unsigned(1,8) ,
47937	 => std_logic_vector(to_unsigned(2,8) ,
47938	 => std_logic_vector(to_unsigned(4,8) ,
47939	 => std_logic_vector(to_unsigned(5,8) ,
47940	 => std_logic_vector(to_unsigned(2,8) ,
47941	 => std_logic_vector(to_unsigned(1,8) ,
47942	 => std_logic_vector(to_unsigned(12,8) ,
47943	 => std_logic_vector(to_unsigned(107,8) ,
47944	 => std_logic_vector(to_unsigned(146,8) ,
47945	 => std_logic_vector(to_unsigned(119,8) ,
47946	 => std_logic_vector(to_unsigned(161,8) ,
47947	 => std_logic_vector(to_unsigned(134,8) ,
47948	 => std_logic_vector(to_unsigned(9,8) ,
47949	 => std_logic_vector(to_unsigned(3,8) ,
47950	 => std_logic_vector(to_unsigned(8,8) ,
47951	 => std_logic_vector(to_unsigned(7,8) ,
47952	 => std_logic_vector(to_unsigned(5,8) ,
47953	 => std_logic_vector(to_unsigned(2,8) ,
47954	 => std_logic_vector(to_unsigned(1,8) ,
47955	 => std_logic_vector(to_unsigned(1,8) ,
47956	 => std_logic_vector(to_unsigned(1,8) ,
47957	 => std_logic_vector(to_unsigned(1,8) ,
47958	 => std_logic_vector(to_unsigned(1,8) ,
47959	 => std_logic_vector(to_unsigned(11,8) ,
47960	 => std_logic_vector(to_unsigned(80,8) ,
47961	 => std_logic_vector(to_unsigned(71,8) ,
47962	 => std_logic_vector(to_unsigned(3,8) ,
47963	 => std_logic_vector(to_unsigned(0,8) ,
47964	 => std_logic_vector(to_unsigned(1,8) ,
47965	 => std_logic_vector(to_unsigned(2,8) ,
47966	 => std_logic_vector(to_unsigned(6,8) ,
47967	 => std_logic_vector(to_unsigned(4,8) ,
47968	 => std_logic_vector(to_unsigned(3,8) ,
47969	 => std_logic_vector(to_unsigned(42,8) ,
47970	 => std_logic_vector(to_unsigned(82,8) ,
47971	 => std_logic_vector(to_unsigned(53,8) ,
47972	 => std_logic_vector(to_unsigned(58,8) ,
47973	 => std_logic_vector(to_unsigned(74,8) ,
47974	 => std_logic_vector(to_unsigned(80,8) ,
47975	 => std_logic_vector(to_unsigned(70,8) ,
47976	 => std_logic_vector(to_unsigned(54,8) ,
47977	 => std_logic_vector(to_unsigned(74,8) ,
47978	 => std_logic_vector(to_unsigned(87,8) ,
47979	 => std_logic_vector(to_unsigned(79,8) ,
47980	 => std_logic_vector(to_unsigned(73,8) ,
47981	 => std_logic_vector(to_unsigned(61,8) ,
47982	 => std_logic_vector(to_unsigned(57,8) ,
47983	 => std_logic_vector(to_unsigned(59,8) ,
47984	 => std_logic_vector(to_unsigned(52,8) ,
47985	 => std_logic_vector(to_unsigned(47,8) ,
47986	 => std_logic_vector(to_unsigned(46,8) ,
47987	 => std_logic_vector(to_unsigned(50,8) ,
47988	 => std_logic_vector(to_unsigned(86,8) ,
47989	 => std_logic_vector(to_unsigned(56,8) ,
47990	 => std_logic_vector(to_unsigned(73,8) ,
47991	 => std_logic_vector(to_unsigned(103,8) ,
47992	 => std_logic_vector(to_unsigned(82,8) ,
47993	 => std_logic_vector(to_unsigned(105,8) ,
47994	 => std_logic_vector(to_unsigned(60,8) ,
47995	 => std_logic_vector(to_unsigned(38,8) ,
47996	 => std_logic_vector(to_unsigned(51,8) ,
47997	 => std_logic_vector(to_unsigned(46,8) ,
47998	 => std_logic_vector(to_unsigned(25,8) ,
47999	 => std_logic_vector(to_unsigned(31,8) ,
48000	 => std_logic_vector(to_unsigned(22,8) ,
48001	 => std_logic_vector(to_unsigned(101,8) ,
48002	 => std_logic_vector(to_unsigned(95,8) ,
48003	 => std_logic_vector(to_unsigned(87,8) ,
48004	 => std_logic_vector(to_unsigned(90,8) ,
48005	 => std_logic_vector(to_unsigned(86,8) ,
48006	 => std_logic_vector(to_unsigned(77,8) ,
48007	 => std_logic_vector(to_unsigned(69,8) ,
48008	 => std_logic_vector(to_unsigned(69,8) ,
48009	 => std_logic_vector(to_unsigned(46,8) ,
48010	 => std_logic_vector(to_unsigned(29,8) ,
48011	 => std_logic_vector(to_unsigned(34,8) ,
48012	 => std_logic_vector(to_unsigned(30,8) ,
48013	 => std_logic_vector(to_unsigned(25,8) ,
48014	 => std_logic_vector(to_unsigned(29,8) ,
48015	 => std_logic_vector(to_unsigned(47,8) ,
48016	 => std_logic_vector(to_unsigned(99,8) ,
48017	 => std_logic_vector(to_unsigned(96,8) ,
48018	 => std_logic_vector(to_unsigned(97,8) ,
48019	 => std_logic_vector(to_unsigned(101,8) ,
48020	 => std_logic_vector(to_unsigned(99,8) ,
48021	 => std_logic_vector(to_unsigned(104,8) ,
48022	 => std_logic_vector(to_unsigned(105,8) ,
48023	 => std_logic_vector(to_unsigned(105,8) ,
48024	 => std_logic_vector(to_unsigned(105,8) ,
48025	 => std_logic_vector(to_unsigned(90,8) ,
48026	 => std_logic_vector(to_unsigned(103,8) ,
48027	 => std_logic_vector(to_unsigned(101,8) ,
48028	 => std_logic_vector(to_unsigned(93,8) ,
48029	 => std_logic_vector(to_unsigned(93,8) ,
48030	 => std_logic_vector(to_unsigned(92,8) ,
48031	 => std_logic_vector(to_unsigned(90,8) ,
48032	 => std_logic_vector(to_unsigned(100,8) ,
48033	 => std_logic_vector(to_unsigned(115,8) ,
48034	 => std_logic_vector(to_unsigned(146,8) ,
48035	 => std_logic_vector(to_unsigned(144,8) ,
48036	 => std_logic_vector(to_unsigned(142,8) ,
48037	 => std_logic_vector(to_unsigned(151,8) ,
48038	 => std_logic_vector(to_unsigned(144,8) ,
48039	 => std_logic_vector(to_unsigned(149,8) ,
48040	 => std_logic_vector(to_unsigned(156,8) ,
48041	 => std_logic_vector(to_unsigned(141,8) ,
48042	 => std_logic_vector(to_unsigned(128,8) ,
48043	 => std_logic_vector(to_unsigned(149,8) ,
48044	 => std_logic_vector(to_unsigned(114,8) ,
48045	 => std_logic_vector(to_unsigned(104,8) ,
48046	 => std_logic_vector(to_unsigned(97,8) ,
48047	 => std_logic_vector(to_unsigned(81,8) ,
48048	 => std_logic_vector(to_unsigned(69,8) ,
48049	 => std_logic_vector(to_unsigned(58,8) ,
48050	 => std_logic_vector(to_unsigned(67,8) ,
48051	 => std_logic_vector(to_unsigned(76,8) ,
48052	 => std_logic_vector(to_unsigned(71,8) ,
48053	 => std_logic_vector(to_unsigned(54,8) ,
48054	 => std_logic_vector(to_unsigned(60,8) ,
48055	 => std_logic_vector(to_unsigned(65,8) ,
48056	 => std_logic_vector(to_unsigned(69,8) ,
48057	 => std_logic_vector(to_unsigned(66,8) ,
48058	 => std_logic_vector(to_unsigned(72,8) ,
48059	 => std_logic_vector(to_unsigned(82,8) ,
48060	 => std_logic_vector(to_unsigned(81,8) ,
48061	 => std_logic_vector(to_unsigned(93,8) ,
48062	 => std_logic_vector(to_unsigned(97,8) ,
48063	 => std_logic_vector(to_unsigned(88,8) ,
48064	 => std_logic_vector(to_unsigned(92,8) ,
48065	 => std_logic_vector(to_unsigned(85,8) ,
48066	 => std_logic_vector(to_unsigned(90,8) ,
48067	 => std_logic_vector(to_unsigned(93,8) ,
48068	 => std_logic_vector(to_unsigned(74,8) ,
48069	 => std_logic_vector(to_unsigned(49,8) ,
48070	 => std_logic_vector(to_unsigned(51,8) ,
48071	 => std_logic_vector(to_unsigned(47,8) ,
48072	 => std_logic_vector(to_unsigned(49,8) ,
48073	 => std_logic_vector(to_unsigned(58,8) ,
48074	 => std_logic_vector(to_unsigned(57,8) ,
48075	 => std_logic_vector(to_unsigned(45,8) ,
48076	 => std_logic_vector(to_unsigned(61,8) ,
48077	 => std_logic_vector(to_unsigned(86,8) ,
48078	 => std_logic_vector(to_unsigned(73,8) ,
48079	 => std_logic_vector(to_unsigned(68,8) ,
48080	 => std_logic_vector(to_unsigned(77,8) ,
48081	 => std_logic_vector(to_unsigned(64,8) ,
48082	 => std_logic_vector(to_unsigned(58,8) ,
48083	 => std_logic_vector(to_unsigned(66,8) ,
48084	 => std_logic_vector(to_unsigned(72,8) ,
48085	 => std_logic_vector(to_unsigned(69,8) ,
48086	 => std_logic_vector(to_unsigned(60,8) ,
48087	 => std_logic_vector(to_unsigned(58,8) ,
48088	 => std_logic_vector(to_unsigned(52,8) ,
48089	 => std_logic_vector(to_unsigned(40,8) ,
48090	 => std_logic_vector(to_unsigned(42,8) ,
48091	 => std_logic_vector(to_unsigned(42,8) ,
48092	 => std_logic_vector(to_unsigned(45,8) ,
48093	 => std_logic_vector(to_unsigned(43,8) ,
48094	 => std_logic_vector(to_unsigned(38,8) ,
48095	 => std_logic_vector(to_unsigned(53,8) ,
48096	 => std_logic_vector(to_unsigned(47,8) ,
48097	 => std_logic_vector(to_unsigned(54,8) ,
48098	 => std_logic_vector(to_unsigned(61,8) ,
48099	 => std_logic_vector(to_unsigned(61,8) ,
48100	 => std_logic_vector(to_unsigned(55,8) ,
48101	 => std_logic_vector(to_unsigned(50,8) ,
48102	 => std_logic_vector(to_unsigned(51,8) ,
48103	 => std_logic_vector(to_unsigned(72,8) ,
48104	 => std_logic_vector(to_unsigned(100,8) ,
48105	 => std_logic_vector(to_unsigned(78,8) ,
48106	 => std_logic_vector(to_unsigned(76,8) ,
48107	 => std_logic_vector(to_unsigned(74,8) ,
48108	 => std_logic_vector(to_unsigned(72,8) ,
48109	 => std_logic_vector(to_unsigned(67,8) ,
48110	 => std_logic_vector(to_unsigned(79,8) ,
48111	 => std_logic_vector(to_unsigned(111,8) ,
48112	 => std_logic_vector(to_unsigned(86,8) ,
48113	 => std_logic_vector(to_unsigned(76,8) ,
48114	 => std_logic_vector(to_unsigned(81,8) ,
48115	 => std_logic_vector(to_unsigned(101,8) ,
48116	 => std_logic_vector(to_unsigned(76,8) ,
48117	 => std_logic_vector(to_unsigned(61,8) ,
48118	 => std_logic_vector(to_unsigned(57,8) ,
48119	 => std_logic_vector(to_unsigned(53,8) ,
48120	 => std_logic_vector(to_unsigned(51,8) ,
48121	 => std_logic_vector(to_unsigned(49,8) ,
48122	 => std_logic_vector(to_unsigned(41,8) ,
48123	 => std_logic_vector(to_unsigned(40,8) ,
48124	 => std_logic_vector(to_unsigned(38,8) ,
48125	 => std_logic_vector(to_unsigned(65,8) ,
48126	 => std_logic_vector(to_unsigned(63,8) ,
48127	 => std_logic_vector(to_unsigned(69,8) ,
48128	 => std_logic_vector(to_unsigned(77,8) ,
48129	 => std_logic_vector(to_unsigned(71,8) ,
48130	 => std_logic_vector(to_unsigned(72,8) ,
48131	 => std_logic_vector(to_unsigned(92,8) ,
48132	 => std_logic_vector(to_unsigned(93,8) ,
48133	 => std_logic_vector(to_unsigned(78,8) ,
48134	 => std_logic_vector(to_unsigned(76,8) ,
48135	 => std_logic_vector(to_unsigned(56,8) ,
48136	 => std_logic_vector(to_unsigned(35,8) ,
48137	 => std_logic_vector(to_unsigned(25,8) ,
48138	 => std_logic_vector(to_unsigned(28,8) ,
48139	 => std_logic_vector(to_unsigned(29,8) ,
48140	 => std_logic_vector(to_unsigned(46,8) ,
48141	 => std_logic_vector(to_unsigned(45,8) ,
48142	 => std_logic_vector(to_unsigned(49,8) ,
48143	 => std_logic_vector(to_unsigned(50,8) ,
48144	 => std_logic_vector(to_unsigned(51,8) ,
48145	 => std_logic_vector(to_unsigned(59,8) ,
48146	 => std_logic_vector(to_unsigned(70,8) ,
48147	 => std_logic_vector(to_unsigned(87,8) ,
48148	 => std_logic_vector(to_unsigned(92,8) ,
48149	 => std_logic_vector(to_unsigned(62,8) ,
48150	 => std_logic_vector(to_unsigned(78,8) ,
48151	 => std_logic_vector(to_unsigned(88,8) ,
48152	 => std_logic_vector(to_unsigned(68,8) ,
48153	 => std_logic_vector(to_unsigned(51,8) ,
48154	 => std_logic_vector(to_unsigned(72,8) ,
48155	 => std_logic_vector(to_unsigned(67,8) ,
48156	 => std_logic_vector(to_unsigned(68,8) ,
48157	 => std_logic_vector(to_unsigned(87,8) ,
48158	 => std_logic_vector(to_unsigned(69,8) ,
48159	 => std_logic_vector(to_unsigned(61,8) ,
48160	 => std_logic_vector(to_unsigned(97,8) ,
48161	 => std_logic_vector(to_unsigned(99,8) ,
48162	 => std_logic_vector(to_unsigned(36,8) ,
48163	 => std_logic_vector(to_unsigned(34,8) ,
48164	 => std_logic_vector(to_unsigned(51,8) ,
48165	 => std_logic_vector(to_unsigned(22,8) ,
48166	 => std_logic_vector(to_unsigned(21,8) ,
48167	 => std_logic_vector(to_unsigned(34,8) ,
48168	 => std_logic_vector(to_unsigned(39,8) ,
48169	 => std_logic_vector(to_unsigned(37,8) ,
48170	 => std_logic_vector(to_unsigned(45,8) ,
48171	 => std_logic_vector(to_unsigned(36,8) ,
48172	 => std_logic_vector(to_unsigned(45,8) ,
48173	 => std_logic_vector(to_unsigned(59,8) ,
48174	 => std_logic_vector(to_unsigned(50,8) ,
48175	 => std_logic_vector(to_unsigned(54,8) ,
48176	 => std_logic_vector(to_unsigned(62,8) ,
48177	 => std_logic_vector(to_unsigned(45,8) ,
48178	 => std_logic_vector(to_unsigned(27,8) ,
48179	 => std_logic_vector(to_unsigned(30,8) ,
48180	 => std_logic_vector(to_unsigned(43,8) ,
48181	 => std_logic_vector(to_unsigned(51,8) ,
48182	 => std_logic_vector(to_unsigned(34,8) ,
48183	 => std_logic_vector(to_unsigned(47,8) ,
48184	 => std_logic_vector(to_unsigned(57,8) ,
48185	 => std_logic_vector(to_unsigned(69,8) ,
48186	 => std_logic_vector(to_unsigned(60,8) ,
48187	 => std_logic_vector(to_unsigned(24,8) ,
48188	 => std_logic_vector(to_unsigned(21,8) ,
48189	 => std_logic_vector(to_unsigned(10,8) ,
48190	 => std_logic_vector(to_unsigned(22,8) ,
48191	 => std_logic_vector(to_unsigned(41,8) ,
48192	 => std_logic_vector(to_unsigned(40,8) ,
48193	 => std_logic_vector(to_unsigned(39,8) ,
48194	 => std_logic_vector(to_unsigned(41,8) ,
48195	 => std_logic_vector(to_unsigned(37,8) ,
48196	 => std_logic_vector(to_unsigned(40,8) ,
48197	 => std_logic_vector(to_unsigned(71,8) ,
48198	 => std_logic_vector(to_unsigned(87,8) ,
48199	 => std_logic_vector(to_unsigned(29,8) ,
48200	 => std_logic_vector(to_unsigned(25,8) ,
48201	 => std_logic_vector(to_unsigned(31,8) ,
48202	 => std_logic_vector(to_unsigned(29,8) ,
48203	 => std_logic_vector(to_unsigned(32,8) ,
48204	 => std_logic_vector(to_unsigned(29,8) ,
48205	 => std_logic_vector(to_unsigned(24,8) ,
48206	 => std_logic_vector(to_unsigned(42,8) ,
48207	 => std_logic_vector(to_unsigned(47,8) ,
48208	 => std_logic_vector(to_unsigned(51,8) ,
48209	 => std_logic_vector(to_unsigned(51,8) ,
48210	 => std_logic_vector(to_unsigned(30,8) ,
48211	 => std_logic_vector(to_unsigned(26,8) ,
48212	 => std_logic_vector(to_unsigned(30,8) ,
48213	 => std_logic_vector(to_unsigned(34,8) ,
48214	 => std_logic_vector(to_unsigned(27,8) ,
48215	 => std_logic_vector(to_unsigned(29,8) ,
48216	 => std_logic_vector(to_unsigned(49,8) ,
48217	 => std_logic_vector(to_unsigned(30,8) ,
48218	 => std_logic_vector(to_unsigned(24,8) ,
48219	 => std_logic_vector(to_unsigned(52,8) ,
48220	 => std_logic_vector(to_unsigned(51,8) ,
48221	 => std_logic_vector(to_unsigned(55,8) ,
48222	 => std_logic_vector(to_unsigned(53,8) ,
48223	 => std_logic_vector(to_unsigned(43,8) ,
48224	 => std_logic_vector(to_unsigned(51,8) ,
48225	 => std_logic_vector(to_unsigned(54,8) ,
48226	 => std_logic_vector(to_unsigned(54,8) ,
48227	 => std_logic_vector(to_unsigned(49,8) ,
48228	 => std_logic_vector(to_unsigned(62,8) ,
48229	 => std_logic_vector(to_unsigned(55,8) ,
48230	 => std_logic_vector(to_unsigned(53,8) ,
48231	 => std_logic_vector(to_unsigned(64,8) ,
48232	 => std_logic_vector(to_unsigned(70,8) ,
48233	 => std_logic_vector(to_unsigned(62,8) ,
48234	 => std_logic_vector(to_unsigned(59,8) ,
48235	 => std_logic_vector(to_unsigned(55,8) ,
48236	 => std_logic_vector(to_unsigned(54,8) ,
48237	 => std_logic_vector(to_unsigned(54,8) ,
48238	 => std_logic_vector(to_unsigned(52,8) ,
48239	 => std_logic_vector(to_unsigned(54,8) ,
48240	 => std_logic_vector(to_unsigned(60,8) ,
48241	 => std_logic_vector(to_unsigned(48,8) ,
48242	 => std_logic_vector(to_unsigned(63,8) ,
48243	 => std_logic_vector(to_unsigned(91,8) ,
48244	 => std_logic_vector(to_unsigned(78,8) ,
48245	 => std_logic_vector(to_unsigned(64,8) ,
48246	 => std_logic_vector(to_unsigned(48,8) ,
48247	 => std_logic_vector(to_unsigned(48,8) ,
48248	 => std_logic_vector(to_unsigned(49,8) ,
48249	 => std_logic_vector(to_unsigned(12,8) ,
48250	 => std_logic_vector(to_unsigned(1,8) ,
48251	 => std_logic_vector(to_unsigned(3,8) ,
48252	 => std_logic_vector(to_unsigned(65,8) ,
48253	 => std_logic_vector(to_unsigned(92,8) ,
48254	 => std_logic_vector(to_unsigned(107,8) ,
48255	 => std_logic_vector(to_unsigned(74,8) ,
48256	 => std_logic_vector(to_unsigned(1,8) ,
48257	 => std_logic_vector(to_unsigned(1,8) ,
48258	 => std_logic_vector(to_unsigned(3,8) ,
48259	 => std_logic_vector(to_unsigned(4,8) ,
48260	 => std_logic_vector(to_unsigned(1,8) ,
48261	 => std_logic_vector(to_unsigned(5,8) ,
48262	 => std_logic_vector(to_unsigned(80,8) ,
48263	 => std_logic_vector(to_unsigned(114,8) ,
48264	 => std_logic_vector(to_unsigned(119,8) ,
48265	 => std_logic_vector(to_unsigned(86,8) ,
48266	 => std_logic_vector(to_unsigned(151,8) ,
48267	 => std_logic_vector(to_unsigned(141,8) ,
48268	 => std_logic_vector(to_unsigned(8,8) ,
48269	 => std_logic_vector(to_unsigned(3,8) ,
48270	 => std_logic_vector(to_unsigned(11,8) ,
48271	 => std_logic_vector(to_unsigned(8,8) ,
48272	 => std_logic_vector(to_unsigned(5,8) ,
48273	 => std_logic_vector(to_unsigned(1,8) ,
48274	 => std_logic_vector(to_unsigned(7,8) ,
48275	 => std_logic_vector(to_unsigned(8,8) ,
48276	 => std_logic_vector(to_unsigned(0,8) ,
48277	 => std_logic_vector(to_unsigned(1,8) ,
48278	 => std_logic_vector(to_unsigned(1,8) ,
48279	 => std_logic_vector(to_unsigned(5,8) ,
48280	 => std_logic_vector(to_unsigned(54,8) ,
48281	 => std_logic_vector(to_unsigned(54,8) ,
48282	 => std_logic_vector(to_unsigned(6,8) ,
48283	 => std_logic_vector(to_unsigned(2,8) ,
48284	 => std_logic_vector(to_unsigned(4,8) ,
48285	 => std_logic_vector(to_unsigned(5,8) ,
48286	 => std_logic_vector(to_unsigned(6,8) ,
48287	 => std_logic_vector(to_unsigned(9,8) ,
48288	 => std_logic_vector(to_unsigned(9,8) ,
48289	 => std_logic_vector(to_unsigned(31,8) ,
48290	 => std_logic_vector(to_unsigned(47,8) ,
48291	 => std_logic_vector(to_unsigned(48,8) ,
48292	 => std_logic_vector(to_unsigned(51,8) ,
48293	 => std_logic_vector(to_unsigned(66,8) ,
48294	 => std_logic_vector(to_unsigned(79,8) ,
48295	 => std_logic_vector(to_unsigned(70,8) ,
48296	 => std_logic_vector(to_unsigned(48,8) ,
48297	 => std_logic_vector(to_unsigned(53,8) ,
48298	 => std_logic_vector(to_unsigned(69,8) ,
48299	 => std_logic_vector(to_unsigned(46,8) ,
48300	 => std_logic_vector(to_unsigned(24,8) ,
48301	 => std_logic_vector(to_unsigned(36,8) ,
48302	 => std_logic_vector(to_unsigned(52,8) ,
48303	 => std_logic_vector(to_unsigned(49,8) ,
48304	 => std_logic_vector(to_unsigned(51,8) ,
48305	 => std_logic_vector(to_unsigned(53,8) ,
48306	 => std_logic_vector(to_unsigned(41,8) ,
48307	 => std_logic_vector(to_unsigned(31,8) ,
48308	 => std_logic_vector(to_unsigned(61,8) ,
48309	 => std_logic_vector(to_unsigned(90,8) ,
48310	 => std_logic_vector(to_unsigned(78,8) ,
48311	 => std_logic_vector(to_unsigned(88,8) ,
48312	 => std_logic_vector(to_unsigned(96,8) ,
48313	 => std_logic_vector(to_unsigned(93,8) ,
48314	 => std_logic_vector(to_unsigned(86,8) ,
48315	 => std_logic_vector(to_unsigned(67,8) ,
48316	 => std_logic_vector(to_unsigned(84,8) ,
48317	 => std_logic_vector(to_unsigned(105,8) ,
48318	 => std_logic_vector(to_unsigned(88,8) ,
48319	 => std_logic_vector(to_unsigned(109,8) ,
48320	 => std_logic_vector(to_unsigned(92,8) ,
48321	 => std_logic_vector(to_unsigned(97,8) ,
48322	 => std_logic_vector(to_unsigned(97,8) ,
48323	 => std_logic_vector(to_unsigned(97,8) ,
48324	 => std_logic_vector(to_unsigned(91,8) ,
48325	 => std_logic_vector(to_unsigned(85,8) ,
48326	 => std_logic_vector(to_unsigned(84,8) ,
48327	 => std_logic_vector(to_unsigned(86,8) ,
48328	 => std_logic_vector(to_unsigned(82,8) ,
48329	 => std_logic_vector(to_unsigned(61,8) ,
48330	 => std_logic_vector(to_unsigned(34,8) ,
48331	 => std_logic_vector(to_unsigned(39,8) ,
48332	 => std_logic_vector(to_unsigned(38,8) ,
48333	 => std_logic_vector(to_unsigned(28,8) ,
48334	 => std_logic_vector(to_unsigned(29,8) ,
48335	 => std_logic_vector(to_unsigned(61,8) ,
48336	 => std_logic_vector(to_unsigned(103,8) ,
48337	 => std_logic_vector(to_unsigned(97,8) ,
48338	 => std_logic_vector(to_unsigned(101,8) ,
48339	 => std_logic_vector(to_unsigned(100,8) ,
48340	 => std_logic_vector(to_unsigned(97,8) ,
48341	 => std_logic_vector(to_unsigned(99,8) ,
48342	 => std_logic_vector(to_unsigned(99,8) ,
48343	 => std_logic_vector(to_unsigned(104,8) ,
48344	 => std_logic_vector(to_unsigned(108,8) ,
48345	 => std_logic_vector(to_unsigned(96,8) ,
48346	 => std_logic_vector(to_unsigned(104,8) ,
48347	 => std_logic_vector(to_unsigned(101,8) ,
48348	 => std_logic_vector(to_unsigned(100,8) ,
48349	 => std_logic_vector(to_unsigned(108,8) ,
48350	 => std_logic_vector(to_unsigned(100,8) ,
48351	 => std_logic_vector(to_unsigned(99,8) ,
48352	 => std_logic_vector(to_unsigned(103,8) ,
48353	 => std_logic_vector(to_unsigned(115,8) ,
48354	 => std_logic_vector(to_unsigned(139,8) ,
48355	 => std_logic_vector(to_unsigned(130,8) ,
48356	 => std_logic_vector(to_unsigned(125,8) ,
48357	 => std_logic_vector(to_unsigned(136,8) ,
48358	 => std_logic_vector(to_unsigned(133,8) ,
48359	 => std_logic_vector(to_unsigned(139,8) ,
48360	 => std_logic_vector(to_unsigned(142,8) ,
48361	 => std_logic_vector(to_unsigned(104,8) ,
48362	 => std_logic_vector(to_unsigned(101,8) ,
48363	 => std_logic_vector(to_unsigned(119,8) ,
48364	 => std_logic_vector(to_unsigned(90,8) ,
48365	 => std_logic_vector(to_unsigned(100,8) ,
48366	 => std_logic_vector(to_unsigned(107,8) ,
48367	 => std_logic_vector(to_unsigned(84,8) ,
48368	 => std_logic_vector(to_unsigned(76,8) ,
48369	 => std_logic_vector(to_unsigned(100,8) ,
48370	 => std_logic_vector(to_unsigned(76,8) ,
48371	 => std_logic_vector(to_unsigned(64,8) ,
48372	 => std_logic_vector(to_unsigned(69,8) ,
48373	 => std_logic_vector(to_unsigned(68,8) ,
48374	 => std_logic_vector(to_unsigned(72,8) ,
48375	 => std_logic_vector(to_unsigned(73,8) ,
48376	 => std_logic_vector(to_unsigned(86,8) ,
48377	 => std_logic_vector(to_unsigned(90,8) ,
48378	 => std_logic_vector(to_unsigned(85,8) ,
48379	 => std_logic_vector(to_unsigned(91,8) ,
48380	 => std_logic_vector(to_unsigned(96,8) ,
48381	 => std_logic_vector(to_unsigned(116,8) ,
48382	 => std_logic_vector(to_unsigned(111,8) ,
48383	 => std_logic_vector(to_unsigned(101,8) ,
48384	 => std_logic_vector(to_unsigned(109,8) ,
48385	 => std_logic_vector(to_unsigned(95,8) ,
48386	 => std_logic_vector(to_unsigned(74,8) ,
48387	 => std_logic_vector(to_unsigned(82,8) ,
48388	 => std_logic_vector(to_unsigned(79,8) ,
48389	 => std_logic_vector(to_unsigned(50,8) ,
48390	 => std_logic_vector(to_unsigned(43,8) ,
48391	 => std_logic_vector(to_unsigned(49,8) ,
48392	 => std_logic_vector(to_unsigned(48,8) ,
48393	 => std_logic_vector(to_unsigned(47,8) ,
48394	 => std_logic_vector(to_unsigned(46,8) ,
48395	 => std_logic_vector(to_unsigned(41,8) ,
48396	 => std_logic_vector(to_unsigned(57,8) ,
48397	 => std_logic_vector(to_unsigned(86,8) ,
48398	 => std_logic_vector(to_unsigned(71,8) ,
48399	 => std_logic_vector(to_unsigned(59,8) ,
48400	 => std_logic_vector(to_unsigned(71,8) ,
48401	 => std_logic_vector(to_unsigned(61,8) ,
48402	 => std_logic_vector(to_unsigned(62,8) ,
48403	 => std_logic_vector(to_unsigned(69,8) ,
48404	 => std_logic_vector(to_unsigned(61,8) ,
48405	 => std_logic_vector(to_unsigned(65,8) ,
48406	 => std_logic_vector(to_unsigned(72,8) ,
48407	 => std_logic_vector(to_unsigned(58,8) ,
48408	 => std_logic_vector(to_unsigned(50,8) ,
48409	 => std_logic_vector(to_unsigned(42,8) ,
48410	 => std_logic_vector(to_unsigned(44,8) ,
48411	 => std_logic_vector(to_unsigned(41,8) ,
48412	 => std_logic_vector(to_unsigned(45,8) ,
48413	 => std_logic_vector(to_unsigned(42,8) ,
48414	 => std_logic_vector(to_unsigned(40,8) ,
48415	 => std_logic_vector(to_unsigned(54,8) ,
48416	 => std_logic_vector(to_unsigned(48,8) ,
48417	 => std_logic_vector(to_unsigned(48,8) ,
48418	 => std_logic_vector(to_unsigned(45,8) ,
48419	 => std_logic_vector(to_unsigned(50,8) ,
48420	 => std_logic_vector(to_unsigned(62,8) ,
48421	 => std_logic_vector(to_unsigned(68,8) ,
48422	 => std_logic_vector(to_unsigned(54,8) ,
48423	 => std_logic_vector(to_unsigned(56,8) ,
48424	 => std_logic_vector(to_unsigned(95,8) ,
48425	 => std_logic_vector(to_unsigned(81,8) ,
48426	 => std_logic_vector(to_unsigned(71,8) ,
48427	 => std_logic_vector(to_unsigned(76,8) ,
48428	 => std_logic_vector(to_unsigned(77,8) ,
48429	 => std_logic_vector(to_unsigned(73,8) ,
48430	 => std_logic_vector(to_unsigned(76,8) ,
48431	 => std_logic_vector(to_unsigned(109,8) ,
48432	 => std_logic_vector(to_unsigned(97,8) ,
48433	 => std_logic_vector(to_unsigned(68,8) ,
48434	 => std_logic_vector(to_unsigned(73,8) ,
48435	 => std_logic_vector(to_unsigned(82,8) ,
48436	 => std_logic_vector(to_unsigned(58,8) ,
48437	 => std_logic_vector(to_unsigned(66,8) ,
48438	 => std_logic_vector(to_unsigned(62,8) ,
48439	 => std_logic_vector(to_unsigned(81,8) ,
48440	 => std_logic_vector(to_unsigned(93,8) ,
48441	 => std_logic_vector(to_unsigned(68,8) ,
48442	 => std_logic_vector(to_unsigned(55,8) ,
48443	 => std_logic_vector(to_unsigned(48,8) ,
48444	 => std_logic_vector(to_unsigned(47,8) ,
48445	 => std_logic_vector(to_unsigned(72,8) ,
48446	 => std_logic_vector(to_unsigned(67,8) ,
48447	 => std_logic_vector(to_unsigned(70,8) ,
48448	 => std_logic_vector(to_unsigned(68,8) ,
48449	 => std_logic_vector(to_unsigned(55,8) ,
48450	 => std_logic_vector(to_unsigned(58,8) ,
48451	 => std_logic_vector(to_unsigned(73,8) ,
48452	 => std_logic_vector(to_unsigned(91,8) ,
48453	 => std_logic_vector(to_unsigned(95,8) ,
48454	 => std_logic_vector(to_unsigned(74,8) ,
48455	 => std_logic_vector(to_unsigned(42,8) ,
48456	 => std_logic_vector(to_unsigned(30,8) ,
48457	 => std_logic_vector(to_unsigned(21,8) ,
48458	 => std_logic_vector(to_unsigned(25,8) ,
48459	 => std_logic_vector(to_unsigned(31,8) ,
48460	 => std_logic_vector(to_unsigned(51,8) ,
48461	 => std_logic_vector(to_unsigned(37,8) ,
48462	 => std_logic_vector(to_unsigned(30,8) ,
48463	 => std_logic_vector(to_unsigned(36,8) ,
48464	 => std_logic_vector(to_unsigned(31,8) ,
48465	 => std_logic_vector(to_unsigned(23,8) ,
48466	 => std_logic_vector(to_unsigned(36,8) ,
48467	 => std_logic_vector(to_unsigned(43,8) ,
48468	 => std_logic_vector(to_unsigned(37,8) ,
48469	 => std_logic_vector(to_unsigned(30,8) ,
48470	 => std_logic_vector(to_unsigned(35,8) ,
48471	 => std_logic_vector(to_unsigned(41,8) ,
48472	 => std_logic_vector(to_unsigned(43,8) ,
48473	 => std_logic_vector(to_unsigned(56,8) ,
48474	 => std_logic_vector(to_unsigned(51,8) ,
48475	 => std_logic_vector(to_unsigned(44,8) ,
48476	 => std_logic_vector(to_unsigned(58,8) ,
48477	 => std_logic_vector(to_unsigned(84,8) ,
48478	 => std_logic_vector(to_unsigned(92,8) ,
48479	 => std_logic_vector(to_unsigned(88,8) ,
48480	 => std_logic_vector(to_unsigned(70,8) ,
48481	 => std_logic_vector(to_unsigned(78,8) ,
48482	 => std_logic_vector(to_unsigned(51,8) ,
48483	 => std_logic_vector(to_unsigned(51,8) ,
48484	 => std_logic_vector(to_unsigned(41,8) ,
48485	 => std_logic_vector(to_unsigned(40,8) ,
48486	 => std_logic_vector(to_unsigned(63,8) ,
48487	 => std_logic_vector(to_unsigned(59,8) ,
48488	 => std_logic_vector(to_unsigned(63,8) ,
48489	 => std_logic_vector(to_unsigned(58,8) ,
48490	 => std_logic_vector(to_unsigned(43,8) ,
48491	 => std_logic_vector(to_unsigned(58,8) ,
48492	 => std_logic_vector(to_unsigned(85,8) ,
48493	 => std_logic_vector(to_unsigned(70,8) ,
48494	 => std_logic_vector(to_unsigned(39,8) ,
48495	 => std_logic_vector(to_unsigned(33,8) ,
48496	 => std_logic_vector(to_unsigned(54,8) ,
48497	 => std_logic_vector(to_unsigned(37,8) ,
48498	 => std_logic_vector(to_unsigned(16,8) ,
48499	 => std_logic_vector(to_unsigned(18,8) ,
48500	 => std_logic_vector(to_unsigned(23,8) ,
48501	 => std_logic_vector(to_unsigned(59,8) ,
48502	 => std_logic_vector(to_unsigned(51,8) ,
48503	 => std_logic_vector(to_unsigned(61,8) ,
48504	 => std_logic_vector(to_unsigned(59,8) ,
48505	 => std_logic_vector(to_unsigned(41,8) ,
48506	 => std_logic_vector(to_unsigned(52,8) ,
48507	 => std_logic_vector(to_unsigned(52,8) ,
48508	 => std_logic_vector(to_unsigned(46,8) ,
48509	 => std_logic_vector(to_unsigned(70,8) ,
48510	 => std_logic_vector(to_unsigned(48,8) ,
48511	 => std_logic_vector(to_unsigned(32,8) ,
48512	 => std_logic_vector(to_unsigned(22,8) ,
48513	 => std_logic_vector(to_unsigned(19,8) ,
48514	 => std_logic_vector(to_unsigned(32,8) ,
48515	 => std_logic_vector(to_unsigned(34,8) ,
48516	 => std_logic_vector(to_unsigned(27,8) ,
48517	 => std_logic_vector(to_unsigned(54,8) ,
48518	 => std_logic_vector(to_unsigned(62,8) ,
48519	 => std_logic_vector(to_unsigned(21,8) ,
48520	 => std_logic_vector(to_unsigned(27,8) ,
48521	 => std_logic_vector(to_unsigned(33,8) ,
48522	 => std_logic_vector(to_unsigned(32,8) ,
48523	 => std_logic_vector(to_unsigned(27,8) ,
48524	 => std_logic_vector(to_unsigned(24,8) ,
48525	 => std_logic_vector(to_unsigned(27,8) ,
48526	 => std_logic_vector(to_unsigned(41,8) ,
48527	 => std_logic_vector(to_unsigned(29,8) ,
48528	 => std_logic_vector(to_unsigned(34,8) ,
48529	 => std_logic_vector(to_unsigned(52,8) ,
48530	 => std_logic_vector(to_unsigned(25,8) ,
48531	 => std_logic_vector(to_unsigned(26,8) ,
48532	 => std_logic_vector(to_unsigned(27,8) ,
48533	 => std_logic_vector(to_unsigned(27,8) ,
48534	 => std_logic_vector(to_unsigned(29,8) ,
48535	 => std_logic_vector(to_unsigned(24,8) ,
48536	 => std_logic_vector(to_unsigned(37,8) ,
48537	 => std_logic_vector(to_unsigned(36,8) ,
48538	 => std_logic_vector(to_unsigned(20,8) ,
48539	 => std_logic_vector(to_unsigned(30,8) ,
48540	 => std_logic_vector(to_unsigned(41,8) ,
48541	 => std_logic_vector(to_unsigned(52,8) ,
48542	 => std_logic_vector(to_unsigned(48,8) ,
48543	 => std_logic_vector(to_unsigned(37,8) ,
48544	 => std_logic_vector(to_unsigned(51,8) ,
48545	 => std_logic_vector(to_unsigned(67,8) ,
48546	 => std_logic_vector(to_unsigned(56,8) ,
48547	 => std_logic_vector(to_unsigned(51,8) ,
48548	 => std_logic_vector(to_unsigned(65,8) ,
48549	 => std_logic_vector(to_unsigned(50,8) ,
48550	 => std_logic_vector(to_unsigned(54,8) ,
48551	 => std_logic_vector(to_unsigned(60,8) ,
48552	 => std_logic_vector(to_unsigned(55,8) ,
48553	 => std_logic_vector(to_unsigned(54,8) ,
48554	 => std_logic_vector(to_unsigned(54,8) ,
48555	 => std_logic_vector(to_unsigned(49,8) ,
48556	 => std_logic_vector(to_unsigned(51,8) ,
48557	 => std_logic_vector(to_unsigned(53,8) ,
48558	 => std_logic_vector(to_unsigned(51,8) ,
48559	 => std_logic_vector(to_unsigned(50,8) ,
48560	 => std_logic_vector(to_unsigned(50,8) ,
48561	 => std_logic_vector(to_unsigned(38,8) ,
48562	 => std_logic_vector(to_unsigned(36,8) ,
48563	 => std_logic_vector(to_unsigned(61,8) ,
48564	 => std_logic_vector(to_unsigned(65,8) ,
48565	 => std_logic_vector(to_unsigned(53,8) ,
48566	 => std_logic_vector(to_unsigned(54,8) ,
48567	 => std_logic_vector(to_unsigned(59,8) ,
48568	 => std_logic_vector(to_unsigned(50,8) ,
48569	 => std_logic_vector(to_unsigned(45,8) ,
48570	 => std_logic_vector(to_unsigned(4,8) ,
48571	 => std_logic_vector(to_unsigned(0,8) ,
48572	 => std_logic_vector(to_unsigned(17,8) ,
48573	 => std_logic_vector(to_unsigned(82,8) ,
48574	 => std_logic_vector(to_unsigned(112,8) ,
48575	 => std_logic_vector(to_unsigned(96,8) ,
48576	 => std_logic_vector(to_unsigned(42,8) ,
48577	 => std_logic_vector(to_unsigned(7,8) ,
48578	 => std_logic_vector(to_unsigned(9,8) ,
48579	 => std_logic_vector(to_unsigned(10,8) ,
48580	 => std_logic_vector(to_unsigned(22,8) ,
48581	 => std_logic_vector(to_unsigned(50,8) ,
48582	 => std_logic_vector(to_unsigned(125,8) ,
48583	 => std_logic_vector(to_unsigned(90,8) ,
48584	 => std_logic_vector(to_unsigned(103,8) ,
48585	 => std_logic_vector(to_unsigned(81,8) ,
48586	 => std_logic_vector(to_unsigned(139,8) ,
48587	 => std_logic_vector(to_unsigned(159,8) ,
48588	 => std_logic_vector(to_unsigned(42,8) ,
48589	 => std_logic_vector(to_unsigned(2,8) ,
48590	 => std_logic_vector(to_unsigned(3,8) ,
48591	 => std_logic_vector(to_unsigned(4,8) ,
48592	 => std_logic_vector(to_unsigned(3,8) ,
48593	 => std_logic_vector(to_unsigned(2,8) ,
48594	 => std_logic_vector(to_unsigned(51,8) ,
48595	 => std_logic_vector(to_unsigned(37,8) ,
48596	 => std_logic_vector(to_unsigned(1,8) ,
48597	 => std_logic_vector(to_unsigned(0,8) ,
48598	 => std_logic_vector(to_unsigned(3,8) ,
48599	 => std_logic_vector(to_unsigned(35,8) ,
48600	 => std_logic_vector(to_unsigned(32,8) ,
48601	 => std_logic_vector(to_unsigned(13,8) ,
48602	 => std_logic_vector(to_unsigned(15,8) ,
48603	 => std_logic_vector(to_unsigned(17,8) ,
48604	 => std_logic_vector(to_unsigned(13,8) ,
48605	 => std_logic_vector(to_unsigned(11,8) ,
48606	 => std_logic_vector(to_unsigned(8,8) ,
48607	 => std_logic_vector(to_unsigned(17,8) ,
48608	 => std_logic_vector(to_unsigned(20,8) ,
48609	 => std_logic_vector(to_unsigned(22,8) ,
48610	 => std_logic_vector(to_unsigned(25,8) ,
48611	 => std_logic_vector(to_unsigned(35,8) ,
48612	 => std_logic_vector(to_unsigned(47,8) ,
48613	 => std_logic_vector(to_unsigned(65,8) ,
48614	 => std_logic_vector(to_unsigned(71,8) ,
48615	 => std_logic_vector(to_unsigned(51,8) ,
48616	 => std_logic_vector(to_unsigned(22,8) ,
48617	 => std_logic_vector(to_unsigned(28,8) ,
48618	 => std_logic_vector(to_unsigned(37,8) ,
48619	 => std_logic_vector(to_unsigned(30,8) ,
48620	 => std_logic_vector(to_unsigned(15,8) ,
48621	 => std_logic_vector(to_unsigned(19,8) ,
48622	 => std_logic_vector(to_unsigned(25,8) ,
48623	 => std_logic_vector(to_unsigned(18,8) ,
48624	 => std_logic_vector(to_unsigned(17,8) ,
48625	 => std_logic_vector(to_unsigned(32,8) ,
48626	 => std_logic_vector(to_unsigned(24,8) ,
48627	 => std_logic_vector(to_unsigned(13,8) ,
48628	 => std_logic_vector(to_unsigned(45,8) ,
48629	 => std_logic_vector(to_unsigned(73,8) ,
48630	 => std_logic_vector(to_unsigned(77,8) ,
48631	 => std_logic_vector(to_unsigned(71,8) ,
48632	 => std_logic_vector(to_unsigned(73,8) ,
48633	 => std_logic_vector(to_unsigned(86,8) ,
48634	 => std_logic_vector(to_unsigned(100,8) ,
48635	 => std_logic_vector(to_unsigned(96,8) ,
48636	 => std_logic_vector(to_unsigned(87,8) ,
48637	 => std_logic_vector(to_unsigned(81,8) ,
48638	 => std_logic_vector(to_unsigned(93,8) ,
48639	 => std_logic_vector(to_unsigned(88,8) ,
48640	 => std_logic_vector(to_unsigned(87,8) ,
48641	 => std_logic_vector(to_unsigned(104,8) ,
48642	 => std_logic_vector(to_unsigned(100,8) ,
48643	 => std_logic_vector(to_unsigned(93,8) ,
48644	 => std_logic_vector(to_unsigned(85,8) ,
48645	 => std_logic_vector(to_unsigned(80,8) ,
48646	 => std_logic_vector(to_unsigned(82,8) ,
48647	 => std_logic_vector(to_unsigned(86,8) ,
48648	 => std_logic_vector(to_unsigned(84,8) ,
48649	 => std_logic_vector(to_unsigned(69,8) ,
48650	 => std_logic_vector(to_unsigned(42,8) ,
48651	 => std_logic_vector(to_unsigned(41,8) ,
48652	 => std_logic_vector(to_unsigned(35,8) ,
48653	 => std_logic_vector(to_unsigned(32,8) ,
48654	 => std_logic_vector(to_unsigned(29,8) ,
48655	 => std_logic_vector(to_unsigned(56,8) ,
48656	 => std_logic_vector(to_unsigned(100,8) ,
48657	 => std_logic_vector(to_unsigned(93,8) ,
48658	 => std_logic_vector(to_unsigned(109,8) ,
48659	 => std_logic_vector(to_unsigned(103,8) ,
48660	 => std_logic_vector(to_unsigned(100,8) ,
48661	 => std_logic_vector(to_unsigned(105,8) ,
48662	 => std_logic_vector(to_unsigned(99,8) ,
48663	 => std_logic_vector(to_unsigned(103,8) ,
48664	 => std_logic_vector(to_unsigned(104,8) ,
48665	 => std_logic_vector(to_unsigned(91,8) ,
48666	 => std_logic_vector(to_unsigned(101,8) ,
48667	 => std_logic_vector(to_unsigned(107,8) ,
48668	 => std_logic_vector(to_unsigned(103,8) ,
48669	 => std_logic_vector(to_unsigned(107,8) ,
48670	 => std_logic_vector(to_unsigned(103,8) ,
48671	 => std_logic_vector(to_unsigned(107,8) ,
48672	 => std_logic_vector(to_unsigned(111,8) ,
48673	 => std_logic_vector(to_unsigned(114,8) ,
48674	 => std_logic_vector(to_unsigned(127,8) ,
48675	 => std_logic_vector(to_unsigned(125,8) ,
48676	 => std_logic_vector(to_unsigned(125,8) ,
48677	 => std_logic_vector(to_unsigned(130,8) ,
48678	 => std_logic_vector(to_unsigned(136,8) ,
48679	 => std_logic_vector(to_unsigned(121,8) ,
48680	 => std_logic_vector(to_unsigned(87,8) ,
48681	 => std_logic_vector(to_unsigned(51,8) ,
48682	 => std_logic_vector(to_unsigned(87,8) ,
48683	 => std_logic_vector(to_unsigned(133,8) ,
48684	 => std_logic_vector(to_unsigned(91,8) ,
48685	 => std_logic_vector(to_unsigned(97,8) ,
48686	 => std_logic_vector(to_unsigned(90,8) ,
48687	 => std_logic_vector(to_unsigned(82,8) ,
48688	 => std_logic_vector(to_unsigned(100,8) ,
48689	 => std_logic_vector(to_unsigned(112,8) ,
48690	 => std_logic_vector(to_unsigned(74,8) ,
48691	 => std_logic_vector(to_unsigned(68,8) ,
48692	 => std_logic_vector(to_unsigned(79,8) ,
48693	 => std_logic_vector(to_unsigned(84,8) ,
48694	 => std_logic_vector(to_unsigned(91,8) ,
48695	 => std_logic_vector(to_unsigned(90,8) ,
48696	 => std_logic_vector(to_unsigned(86,8) ,
48697	 => std_logic_vector(to_unsigned(86,8) ,
48698	 => std_logic_vector(to_unsigned(100,8) ,
48699	 => std_logic_vector(to_unsigned(114,8) ,
48700	 => std_logic_vector(to_unsigned(130,8) ,
48701	 => std_logic_vector(to_unsigned(131,8) ,
48702	 => std_logic_vector(to_unsigned(112,8) ,
48703	 => std_logic_vector(to_unsigned(118,8) ,
48704	 => std_logic_vector(to_unsigned(136,8) ,
48705	 => std_logic_vector(to_unsigned(127,8) ,
48706	 => std_logic_vector(to_unsigned(52,8) ,
48707	 => std_logic_vector(to_unsigned(73,8) ,
48708	 => std_logic_vector(to_unsigned(80,8) ,
48709	 => std_logic_vector(to_unsigned(55,8) ,
48710	 => std_logic_vector(to_unsigned(47,8) ,
48711	 => std_logic_vector(to_unsigned(57,8) ,
48712	 => std_logic_vector(to_unsigned(55,8) ,
48713	 => std_logic_vector(to_unsigned(33,8) ,
48714	 => std_logic_vector(to_unsigned(30,8) ,
48715	 => std_logic_vector(to_unsigned(35,8) ,
48716	 => std_logic_vector(to_unsigned(55,8) ,
48717	 => std_logic_vector(to_unsigned(78,8) ,
48718	 => std_logic_vector(to_unsigned(70,8) ,
48719	 => std_logic_vector(to_unsigned(67,8) ,
48720	 => std_logic_vector(to_unsigned(71,8) ,
48721	 => std_logic_vector(to_unsigned(55,8) ,
48722	 => std_logic_vector(to_unsigned(57,8) ,
48723	 => std_logic_vector(to_unsigned(67,8) ,
48724	 => std_logic_vector(to_unsigned(65,8) ,
48725	 => std_logic_vector(to_unsigned(70,8) ,
48726	 => std_logic_vector(to_unsigned(66,8) ,
48727	 => std_logic_vector(to_unsigned(53,8) ,
48728	 => std_logic_vector(to_unsigned(51,8) ,
48729	 => std_logic_vector(to_unsigned(42,8) ,
48730	 => std_logic_vector(to_unsigned(41,8) ,
48731	 => std_logic_vector(to_unsigned(41,8) ,
48732	 => std_logic_vector(to_unsigned(43,8) ,
48733	 => std_logic_vector(to_unsigned(42,8) ,
48734	 => std_logic_vector(to_unsigned(36,8) ,
48735	 => std_logic_vector(to_unsigned(32,8) ,
48736	 => std_logic_vector(to_unsigned(41,8) ,
48737	 => std_logic_vector(to_unsigned(46,8) ,
48738	 => std_logic_vector(to_unsigned(41,8) ,
48739	 => std_logic_vector(to_unsigned(56,8) ,
48740	 => std_logic_vector(to_unsigned(68,8) ,
48741	 => std_logic_vector(to_unsigned(69,8) ,
48742	 => std_logic_vector(to_unsigned(51,8) ,
48743	 => std_logic_vector(to_unsigned(54,8) ,
48744	 => std_logic_vector(to_unsigned(95,8) ,
48745	 => std_logic_vector(to_unsigned(73,8) ,
48746	 => std_logic_vector(to_unsigned(69,8) ,
48747	 => std_logic_vector(to_unsigned(76,8) ,
48748	 => std_logic_vector(to_unsigned(73,8) ,
48749	 => std_logic_vector(to_unsigned(70,8) ,
48750	 => std_logic_vector(to_unsigned(71,8) ,
48751	 => std_logic_vector(to_unsigned(108,8) ,
48752	 => std_logic_vector(to_unsigned(93,8) ,
48753	 => std_logic_vector(to_unsigned(64,8) ,
48754	 => std_logic_vector(to_unsigned(71,8) ,
48755	 => std_logic_vector(to_unsigned(69,8) ,
48756	 => std_logic_vector(to_unsigned(40,8) ,
48757	 => std_logic_vector(to_unsigned(48,8) ,
48758	 => std_logic_vector(to_unsigned(51,8) ,
48759	 => std_logic_vector(to_unsigned(52,8) ,
48760	 => std_logic_vector(to_unsigned(64,8) ,
48761	 => std_logic_vector(to_unsigned(65,8) ,
48762	 => std_logic_vector(to_unsigned(60,8) ,
48763	 => std_logic_vector(to_unsigned(66,8) ,
48764	 => std_logic_vector(to_unsigned(70,8) ,
48765	 => std_logic_vector(to_unsigned(77,8) ,
48766	 => std_logic_vector(to_unsigned(85,8) ,
48767	 => std_logic_vector(to_unsigned(88,8) ,
48768	 => std_logic_vector(to_unsigned(91,8) ,
48769	 => std_logic_vector(to_unsigned(72,8) ,
48770	 => std_logic_vector(to_unsigned(50,8) ,
48771	 => std_logic_vector(to_unsigned(60,8) ,
48772	 => std_logic_vector(to_unsigned(68,8) ,
48773	 => std_logic_vector(to_unsigned(56,8) ,
48774	 => std_logic_vector(to_unsigned(62,8) ,
48775	 => std_logic_vector(to_unsigned(44,8) ,
48776	 => std_logic_vector(to_unsigned(28,8) ,
48777	 => std_logic_vector(to_unsigned(17,8) ,
48778	 => std_logic_vector(to_unsigned(22,8) ,
48779	 => std_logic_vector(to_unsigned(30,8) ,
48780	 => std_logic_vector(to_unsigned(37,8) ,
48781	 => std_logic_vector(to_unsigned(33,8) ,
48782	 => std_logic_vector(to_unsigned(33,8) ,
48783	 => std_logic_vector(to_unsigned(32,8) ,
48784	 => std_logic_vector(to_unsigned(32,8) ,
48785	 => std_logic_vector(to_unsigned(32,8) ,
48786	 => std_logic_vector(to_unsigned(66,8) ,
48787	 => std_logic_vector(to_unsigned(65,8) ,
48788	 => std_logic_vector(to_unsigned(42,8) ,
48789	 => std_logic_vector(to_unsigned(25,8) ,
48790	 => std_logic_vector(to_unsigned(25,8) ,
48791	 => std_logic_vector(to_unsigned(31,8) ,
48792	 => std_logic_vector(to_unsigned(27,8) ,
48793	 => std_logic_vector(to_unsigned(26,8) ,
48794	 => std_logic_vector(to_unsigned(23,8) ,
48795	 => std_logic_vector(to_unsigned(23,8) ,
48796	 => std_logic_vector(to_unsigned(19,8) ,
48797	 => std_logic_vector(to_unsigned(28,8) ,
48798	 => std_logic_vector(to_unsigned(41,8) ,
48799	 => std_logic_vector(to_unsigned(39,8) ,
48800	 => std_logic_vector(to_unsigned(31,8) ,
48801	 => std_logic_vector(to_unsigned(33,8) ,
48802	 => std_logic_vector(to_unsigned(45,8) ,
48803	 => std_logic_vector(to_unsigned(49,8) ,
48804	 => std_logic_vector(to_unsigned(48,8) ,
48805	 => std_logic_vector(to_unsigned(63,8) ,
48806	 => std_logic_vector(to_unsigned(65,8) ,
48807	 => std_logic_vector(to_unsigned(71,8) ,
48808	 => std_logic_vector(to_unsigned(86,8) ,
48809	 => std_logic_vector(to_unsigned(80,8) ,
48810	 => std_logic_vector(to_unsigned(72,8) ,
48811	 => std_logic_vector(to_unsigned(84,8) ,
48812	 => std_logic_vector(to_unsigned(62,8) ,
48813	 => std_logic_vector(to_unsigned(63,8) ,
48814	 => std_logic_vector(to_unsigned(54,8) ,
48815	 => std_logic_vector(to_unsigned(45,8) ,
48816	 => std_logic_vector(to_unsigned(56,8) ,
48817	 => std_logic_vector(to_unsigned(67,8) ,
48818	 => std_logic_vector(to_unsigned(47,8) ,
48819	 => std_logic_vector(to_unsigned(26,8) ,
48820	 => std_logic_vector(to_unsigned(36,8) ,
48821	 => std_logic_vector(to_unsigned(60,8) ,
48822	 => std_logic_vector(to_unsigned(61,8) ,
48823	 => std_logic_vector(to_unsigned(52,8) ,
48824	 => std_logic_vector(to_unsigned(51,8) ,
48825	 => std_logic_vector(to_unsigned(56,8) ,
48826	 => std_logic_vector(to_unsigned(59,8) ,
48827	 => std_logic_vector(to_unsigned(22,8) ,
48828	 => std_logic_vector(to_unsigned(32,8) ,
48829	 => std_logic_vector(to_unsigned(146,8) ,
48830	 => std_logic_vector(to_unsigned(95,8) ,
48831	 => std_logic_vector(to_unsigned(42,8) ,
48832	 => std_logic_vector(to_unsigned(39,8) ,
48833	 => std_logic_vector(to_unsigned(31,8) ,
48834	 => std_logic_vector(to_unsigned(35,8) ,
48835	 => std_logic_vector(to_unsigned(30,8) ,
48836	 => std_logic_vector(to_unsigned(25,8) ,
48837	 => std_logic_vector(to_unsigned(30,8) ,
48838	 => std_logic_vector(to_unsigned(31,8) ,
48839	 => std_logic_vector(to_unsigned(26,8) ,
48840	 => std_logic_vector(to_unsigned(24,8) ,
48841	 => std_logic_vector(to_unsigned(27,8) ,
48842	 => std_logic_vector(to_unsigned(33,8) ,
48843	 => std_logic_vector(to_unsigned(29,8) ,
48844	 => std_logic_vector(to_unsigned(27,8) ,
48845	 => std_logic_vector(to_unsigned(30,8) ,
48846	 => std_logic_vector(to_unsigned(45,8) ,
48847	 => std_logic_vector(to_unsigned(45,8) ,
48848	 => std_logic_vector(to_unsigned(48,8) ,
48849	 => std_logic_vector(to_unsigned(51,8) ,
48850	 => std_logic_vector(to_unsigned(29,8) ,
48851	 => std_logic_vector(to_unsigned(22,8) ,
48852	 => std_logic_vector(to_unsigned(25,8) ,
48853	 => std_logic_vector(to_unsigned(24,8) ,
48854	 => std_logic_vector(to_unsigned(25,8) ,
48855	 => std_logic_vector(to_unsigned(25,8) ,
48856	 => std_logic_vector(to_unsigned(25,8) ,
48857	 => std_logic_vector(to_unsigned(64,8) ,
48858	 => std_logic_vector(to_unsigned(46,8) ,
48859	 => std_logic_vector(to_unsigned(35,8) ,
48860	 => std_logic_vector(to_unsigned(51,8) ,
48861	 => std_logic_vector(to_unsigned(65,8) ,
48862	 => std_logic_vector(to_unsigned(50,8) ,
48863	 => std_logic_vector(to_unsigned(30,8) ,
48864	 => std_logic_vector(to_unsigned(46,8) ,
48865	 => std_logic_vector(to_unsigned(68,8) ,
48866	 => std_logic_vector(to_unsigned(53,8) ,
48867	 => std_logic_vector(to_unsigned(45,8) ,
48868	 => std_logic_vector(to_unsigned(65,8) ,
48869	 => std_logic_vector(to_unsigned(46,8) ,
48870	 => std_logic_vector(to_unsigned(55,8) ,
48871	 => std_logic_vector(to_unsigned(59,8) ,
48872	 => std_logic_vector(to_unsigned(48,8) ,
48873	 => std_logic_vector(to_unsigned(50,8) ,
48874	 => std_logic_vector(to_unsigned(50,8) ,
48875	 => std_logic_vector(to_unsigned(42,8) ,
48876	 => std_logic_vector(to_unsigned(45,8) ,
48877	 => std_logic_vector(to_unsigned(50,8) ,
48878	 => std_logic_vector(to_unsigned(46,8) ,
48879	 => std_logic_vector(to_unsigned(46,8) ,
48880	 => std_logic_vector(to_unsigned(43,8) ,
48881	 => std_logic_vector(to_unsigned(40,8) ,
48882	 => std_logic_vector(to_unsigned(44,8) ,
48883	 => std_logic_vector(to_unsigned(56,8) ,
48884	 => std_logic_vector(to_unsigned(52,8) ,
48885	 => std_logic_vector(to_unsigned(41,8) ,
48886	 => std_logic_vector(to_unsigned(49,8) ,
48887	 => std_logic_vector(to_unsigned(54,8) ,
48888	 => std_logic_vector(to_unsigned(51,8) ,
48889	 => std_logic_vector(to_unsigned(87,8) ,
48890	 => std_logic_vector(to_unsigned(30,8) ,
48891	 => std_logic_vector(to_unsigned(1,8) ,
48892	 => std_logic_vector(to_unsigned(3,8) ,
48893	 => std_logic_vector(to_unsigned(28,8) ,
48894	 => std_logic_vector(to_unsigned(125,8) ,
48895	 => std_logic_vector(to_unsigned(85,8) ,
48896	 => std_logic_vector(to_unsigned(109,8) ,
48897	 => std_logic_vector(to_unsigned(97,8) ,
48898	 => std_logic_vector(to_unsigned(92,8) ,
48899	 => std_logic_vector(to_unsigned(87,8) ,
48900	 => std_logic_vector(to_unsigned(119,8) ,
48901	 => std_logic_vector(to_unsigned(84,8) ,
48902	 => std_logic_vector(to_unsigned(97,8) ,
48903	 => std_logic_vector(to_unsigned(85,8) ,
48904	 => std_logic_vector(to_unsigned(93,8) ,
48905	 => std_logic_vector(to_unsigned(71,8) ,
48906	 => std_logic_vector(to_unsigned(141,8) ,
48907	 => std_logic_vector(to_unsigned(152,8) ,
48908	 => std_logic_vector(to_unsigned(133,8) ,
48909	 => std_logic_vector(to_unsigned(27,8) ,
48910	 => std_logic_vector(to_unsigned(3,8) ,
48911	 => std_logic_vector(to_unsigned(4,8) ,
48912	 => std_logic_vector(to_unsigned(4,8) ,
48913	 => std_logic_vector(to_unsigned(27,8) ,
48914	 => std_logic_vector(to_unsigned(72,8) ,
48915	 => std_logic_vector(to_unsigned(26,8) ,
48916	 => std_logic_vector(to_unsigned(1,8) ,
48917	 => std_logic_vector(to_unsigned(1,8) ,
48918	 => std_logic_vector(to_unsigned(17,8) ,
48919	 => std_logic_vector(to_unsigned(35,8) ,
48920	 => std_logic_vector(to_unsigned(7,8) ,
48921	 => std_logic_vector(to_unsigned(1,8) ,
48922	 => std_logic_vector(to_unsigned(5,8) ,
48923	 => std_logic_vector(to_unsigned(6,8) ,
48924	 => std_logic_vector(to_unsigned(6,8) ,
48925	 => std_logic_vector(to_unsigned(12,8) ,
48926	 => std_logic_vector(to_unsigned(13,8) ,
48927	 => std_logic_vector(to_unsigned(10,8) ,
48928	 => std_logic_vector(to_unsigned(21,8) ,
48929	 => std_logic_vector(to_unsigned(56,8) ,
48930	 => std_logic_vector(to_unsigned(49,8) ,
48931	 => std_logic_vector(to_unsigned(49,8) ,
48932	 => std_logic_vector(to_unsigned(60,8) ,
48933	 => std_logic_vector(to_unsigned(66,8) ,
48934	 => std_logic_vector(to_unsigned(64,8) ,
48935	 => std_logic_vector(to_unsigned(45,8) ,
48936	 => std_logic_vector(to_unsigned(25,8) ,
48937	 => std_logic_vector(to_unsigned(27,8) ,
48938	 => std_logic_vector(to_unsigned(52,8) ,
48939	 => std_logic_vector(to_unsigned(46,8) ,
48940	 => std_logic_vector(to_unsigned(29,8) ,
48941	 => std_logic_vector(to_unsigned(25,8) ,
48942	 => std_logic_vector(to_unsigned(28,8) ,
48943	 => std_logic_vector(to_unsigned(16,8) ,
48944	 => std_logic_vector(to_unsigned(18,8) ,
48945	 => std_logic_vector(to_unsigned(30,8) ,
48946	 => std_logic_vector(to_unsigned(32,8) ,
48947	 => std_logic_vector(to_unsigned(26,8) ,
48948	 => std_logic_vector(to_unsigned(47,8) ,
48949	 => std_logic_vector(to_unsigned(43,8) ,
48950	 => std_logic_vector(to_unsigned(38,8) ,
48951	 => std_logic_vector(to_unsigned(12,8) ,
48952	 => std_logic_vector(to_unsigned(12,8) ,
48953	 => std_logic_vector(to_unsigned(43,8) ,
48954	 => std_logic_vector(to_unsigned(58,8) ,
48955	 => std_logic_vector(to_unsigned(50,8) ,
48956	 => std_logic_vector(to_unsigned(62,8) ,
48957	 => std_logic_vector(to_unsigned(41,8) ,
48958	 => std_logic_vector(to_unsigned(30,8) ,
48959	 => std_logic_vector(to_unsigned(62,8) ,
48960	 => std_logic_vector(to_unsigned(91,8) ,
48961	 => std_logic_vector(to_unsigned(95,8) ,
48962	 => std_logic_vector(to_unsigned(92,8) ,
48963	 => std_logic_vector(to_unsigned(88,8) ,
48964	 => std_logic_vector(to_unsigned(86,8) ,
48965	 => std_logic_vector(to_unsigned(86,8) ,
48966	 => std_logic_vector(to_unsigned(81,8) ,
48967	 => std_logic_vector(to_unsigned(80,8) ,
48968	 => std_logic_vector(to_unsigned(81,8) ,
48969	 => std_logic_vector(to_unsigned(72,8) ,
48970	 => std_logic_vector(to_unsigned(51,8) ,
48971	 => std_logic_vector(to_unsigned(51,8) ,
48972	 => std_logic_vector(to_unsigned(42,8) ,
48973	 => std_logic_vector(to_unsigned(37,8) ,
48974	 => std_logic_vector(to_unsigned(35,8) ,
48975	 => std_logic_vector(to_unsigned(40,8) ,
48976	 => std_logic_vector(to_unsigned(91,8) ,
48977	 => std_logic_vector(to_unsigned(104,8) ,
48978	 => std_logic_vector(to_unsigned(97,8) ,
48979	 => std_logic_vector(to_unsigned(99,8) ,
48980	 => std_logic_vector(to_unsigned(91,8) ,
48981	 => std_logic_vector(to_unsigned(104,8) ,
48982	 => std_logic_vector(to_unsigned(99,8) ,
48983	 => std_logic_vector(to_unsigned(91,8) ,
48984	 => std_logic_vector(to_unsigned(99,8) ,
48985	 => std_logic_vector(to_unsigned(92,8) ,
48986	 => std_logic_vector(to_unsigned(95,8) ,
48987	 => std_logic_vector(to_unsigned(100,8) ,
48988	 => std_logic_vector(to_unsigned(92,8) ,
48989	 => std_logic_vector(to_unsigned(91,8) ,
48990	 => std_logic_vector(to_unsigned(100,8) ,
48991	 => std_logic_vector(to_unsigned(100,8) ,
48992	 => std_logic_vector(to_unsigned(107,8) ,
48993	 => std_logic_vector(to_unsigned(103,8) ,
48994	 => std_logic_vector(to_unsigned(119,8) ,
48995	 => std_logic_vector(to_unsigned(114,8) ,
48996	 => std_logic_vector(to_unsigned(112,8) ,
48997	 => std_logic_vector(to_unsigned(108,8) ,
48998	 => std_logic_vector(to_unsigned(93,8) ,
48999	 => std_logic_vector(to_unsigned(64,8) ,
49000	 => std_logic_vector(to_unsigned(43,8) ,
49001	 => std_logic_vector(to_unsigned(60,8) ,
49002	 => std_logic_vector(to_unsigned(139,8) ,
49003	 => std_logic_vector(to_unsigned(146,8) ,
49004	 => std_logic_vector(to_unsigned(118,8) ,
49005	 => std_logic_vector(to_unsigned(103,8) ,
49006	 => std_logic_vector(to_unsigned(57,8) ,
49007	 => std_logic_vector(to_unsigned(58,8) ,
49008	 => std_logic_vector(to_unsigned(97,8) ,
49009	 => std_logic_vector(to_unsigned(105,8) ,
49010	 => std_logic_vector(to_unsigned(81,8) ,
49011	 => std_logic_vector(to_unsigned(81,8) ,
49012	 => std_logic_vector(to_unsigned(97,8) ,
49013	 => std_logic_vector(to_unsigned(91,8) ,
49014	 => std_logic_vector(to_unsigned(90,8) ,
49015	 => std_logic_vector(to_unsigned(104,8) ,
49016	 => std_logic_vector(to_unsigned(85,8) ,
49017	 => std_logic_vector(to_unsigned(65,8) ,
49018	 => std_logic_vector(to_unsigned(55,8) ,
49019	 => std_logic_vector(to_unsigned(71,8) ,
49020	 => std_logic_vector(to_unsigned(103,8) ,
49021	 => std_logic_vector(to_unsigned(115,8) ,
49022	 => std_logic_vector(to_unsigned(119,8) ,
49023	 => std_logic_vector(to_unsigned(107,8) ,
49024	 => std_logic_vector(to_unsigned(115,8) ,
49025	 => std_logic_vector(to_unsigned(147,8) ,
49026	 => std_logic_vector(to_unsigned(88,8) ,
49027	 => std_logic_vector(to_unsigned(91,8) ,
49028	 => std_logic_vector(to_unsigned(68,8) ,
49029	 => std_logic_vector(to_unsigned(50,8) ,
49030	 => std_logic_vector(to_unsigned(64,8) ,
49031	 => std_logic_vector(to_unsigned(86,8) ,
49032	 => std_logic_vector(to_unsigned(86,8) ,
49033	 => std_logic_vector(to_unsigned(59,8) ,
49034	 => std_logic_vector(to_unsigned(47,8) ,
49035	 => std_logic_vector(to_unsigned(43,8) ,
49036	 => std_logic_vector(to_unsigned(57,8) ,
49037	 => std_logic_vector(to_unsigned(79,8) ,
49038	 => std_logic_vector(to_unsigned(68,8) ,
49039	 => std_logic_vector(to_unsigned(53,8) ,
49040	 => std_logic_vector(to_unsigned(69,8) ,
49041	 => std_logic_vector(to_unsigned(66,8) ,
49042	 => std_logic_vector(to_unsigned(68,8) ,
49043	 => std_logic_vector(to_unsigned(76,8) ,
49044	 => std_logic_vector(to_unsigned(61,8) ,
49045	 => std_logic_vector(to_unsigned(67,8) ,
49046	 => std_logic_vector(to_unsigned(73,8) ,
49047	 => std_logic_vector(to_unsigned(54,8) ,
49048	 => std_logic_vector(to_unsigned(45,8) ,
49049	 => std_logic_vector(to_unsigned(39,8) ,
49050	 => std_logic_vector(to_unsigned(40,8) ,
49051	 => std_logic_vector(to_unsigned(41,8) ,
49052	 => std_logic_vector(to_unsigned(39,8) ,
49053	 => std_logic_vector(to_unsigned(41,8) ,
49054	 => std_logic_vector(to_unsigned(38,8) ,
49055	 => std_logic_vector(to_unsigned(38,8) ,
49056	 => std_logic_vector(to_unsigned(52,8) ,
49057	 => std_logic_vector(to_unsigned(45,8) ,
49058	 => std_logic_vector(to_unsigned(43,8) ,
49059	 => std_logic_vector(to_unsigned(45,8) ,
49060	 => std_logic_vector(to_unsigned(43,8) ,
49061	 => std_logic_vector(to_unsigned(63,8) ,
49062	 => std_logic_vector(to_unsigned(51,8) ,
49063	 => std_logic_vector(to_unsigned(50,8) ,
49064	 => std_logic_vector(to_unsigned(93,8) ,
49065	 => std_logic_vector(to_unsigned(95,8) ,
49066	 => std_logic_vector(to_unsigned(84,8) ,
49067	 => std_logic_vector(to_unsigned(72,8) ,
49068	 => std_logic_vector(to_unsigned(69,8) ,
49069	 => std_logic_vector(to_unsigned(65,8) ,
49070	 => std_logic_vector(to_unsigned(70,8) ,
49071	 => std_logic_vector(to_unsigned(97,8) ,
49072	 => std_logic_vector(to_unsigned(74,8) ,
49073	 => std_logic_vector(to_unsigned(48,8) ,
49074	 => std_logic_vector(to_unsigned(56,8) ,
49075	 => std_logic_vector(to_unsigned(68,8) ,
49076	 => std_logic_vector(to_unsigned(77,8) ,
49077	 => std_logic_vector(to_unsigned(76,8) ,
49078	 => std_logic_vector(to_unsigned(74,8) ,
49079	 => std_logic_vector(to_unsigned(64,8) ,
49080	 => std_logic_vector(to_unsigned(51,8) ,
49081	 => std_logic_vector(to_unsigned(57,8) ,
49082	 => std_logic_vector(to_unsigned(56,8) ,
49083	 => std_logic_vector(to_unsigned(54,8) ,
49084	 => std_logic_vector(to_unsigned(52,8) ,
49085	 => std_logic_vector(to_unsigned(54,8) ,
49086	 => std_logic_vector(to_unsigned(51,8) ,
49087	 => std_logic_vector(to_unsigned(64,8) ,
49088	 => std_logic_vector(to_unsigned(101,8) ,
49089	 => std_logic_vector(to_unsigned(72,8) ,
49090	 => std_logic_vector(to_unsigned(37,8) ,
49091	 => std_logic_vector(to_unsigned(52,8) ,
49092	 => std_logic_vector(to_unsigned(62,8) ,
49093	 => std_logic_vector(to_unsigned(44,8) ,
49094	 => std_logic_vector(to_unsigned(55,8) ,
49095	 => std_logic_vector(to_unsigned(41,8) ,
49096	 => std_logic_vector(to_unsigned(24,8) ,
49097	 => std_logic_vector(to_unsigned(16,8) ,
49098	 => std_logic_vector(to_unsigned(19,8) ,
49099	 => std_logic_vector(to_unsigned(23,8) ,
49100	 => std_logic_vector(to_unsigned(41,8) ,
49101	 => std_logic_vector(to_unsigned(49,8) ,
49102	 => std_logic_vector(to_unsigned(58,8) ,
49103	 => std_logic_vector(to_unsigned(51,8) ,
49104	 => std_logic_vector(to_unsigned(43,8) ,
49105	 => std_logic_vector(to_unsigned(44,8) ,
49106	 => std_logic_vector(to_unsigned(68,8) ,
49107	 => std_logic_vector(to_unsigned(58,8) ,
49108	 => std_logic_vector(to_unsigned(40,8) ,
49109	 => std_logic_vector(to_unsigned(30,8) ,
49110	 => std_logic_vector(to_unsigned(34,8) ,
49111	 => std_logic_vector(to_unsigned(43,8) ,
49112	 => std_logic_vector(to_unsigned(46,8) ,
49113	 => std_logic_vector(to_unsigned(44,8) ,
49114	 => std_logic_vector(to_unsigned(37,8) ,
49115	 => std_logic_vector(to_unsigned(32,8) ,
49116	 => std_logic_vector(to_unsigned(19,8) ,
49117	 => std_logic_vector(to_unsigned(24,8) ,
49118	 => std_logic_vector(to_unsigned(35,8) ,
49119	 => std_logic_vector(to_unsigned(31,8) ,
49120	 => std_logic_vector(to_unsigned(24,8) ,
49121	 => std_logic_vector(to_unsigned(13,8) ,
49122	 => std_logic_vector(to_unsigned(17,8) ,
49123	 => std_logic_vector(to_unsigned(18,8) ,
49124	 => std_logic_vector(to_unsigned(14,8) ,
49125	 => std_logic_vector(to_unsigned(17,8) ,
49126	 => std_logic_vector(to_unsigned(16,8) ,
49127	 => std_logic_vector(to_unsigned(23,8) ,
49128	 => std_logic_vector(to_unsigned(35,8) ,
49129	 => std_logic_vector(to_unsigned(53,8) ,
49130	 => std_logic_vector(to_unsigned(79,8) ,
49131	 => std_logic_vector(to_unsigned(52,8) ,
49132	 => std_logic_vector(to_unsigned(35,8) ,
49133	 => std_logic_vector(to_unsigned(60,8) ,
49134	 => std_logic_vector(to_unsigned(67,8) ,
49135	 => std_logic_vector(to_unsigned(79,8) ,
49136	 => std_logic_vector(to_unsigned(80,8) ,
49137	 => std_logic_vector(to_unsigned(93,8) ,
49138	 => std_logic_vector(to_unsigned(73,8) ,
49139	 => std_logic_vector(to_unsigned(45,8) ,
49140	 => std_logic_vector(to_unsigned(54,8) ,
49141	 => std_logic_vector(to_unsigned(60,8) ,
49142	 => std_logic_vector(to_unsigned(51,8) ,
49143	 => std_logic_vector(to_unsigned(55,8) ,
49144	 => std_logic_vector(to_unsigned(53,8) ,
49145	 => std_logic_vector(to_unsigned(66,8) ,
49146	 => std_logic_vector(to_unsigned(32,8) ,
49147	 => std_logic_vector(to_unsigned(20,8) ,
49148	 => std_logic_vector(to_unsigned(33,8) ,
49149	 => std_logic_vector(to_unsigned(63,8) ,
49150	 => std_logic_vector(to_unsigned(70,8) ,
49151	 => std_logic_vector(to_unsigned(44,8) ,
49152	 => std_logic_vector(to_unsigned(30,8) ,
49153	 => std_logic_vector(to_unsigned(30,8) ,
49154	 => std_logic_vector(to_unsigned(34,8) ,
49155	 => std_logic_vector(to_unsigned(35,8) ,
49156	 => std_logic_vector(to_unsigned(37,8) ,
49157	 => std_logic_vector(to_unsigned(44,8) ,
49158	 => std_logic_vector(to_unsigned(45,8) ,
49159	 => std_logic_vector(to_unsigned(42,8) ,
49160	 => std_logic_vector(to_unsigned(33,8) ,
49161	 => std_logic_vector(to_unsigned(37,8) ,
49162	 => std_logic_vector(to_unsigned(35,8) ,
49163	 => std_logic_vector(to_unsigned(34,8) ,
49164	 => std_logic_vector(to_unsigned(29,8) ,
49165	 => std_logic_vector(to_unsigned(26,8) ,
49166	 => std_logic_vector(to_unsigned(44,8) ,
49167	 => std_logic_vector(to_unsigned(68,8) ,
49168	 => std_logic_vector(to_unsigned(65,8) ,
49169	 => std_logic_vector(to_unsigned(41,8) ,
49170	 => std_logic_vector(to_unsigned(28,8) ,
49171	 => std_logic_vector(to_unsigned(17,8) ,
49172	 => std_logic_vector(to_unsigned(22,8) ,
49173	 => std_logic_vector(to_unsigned(23,8) ,
49174	 => std_logic_vector(to_unsigned(24,8) ,
49175	 => std_logic_vector(to_unsigned(22,8) ,
49176	 => std_logic_vector(to_unsigned(17,8) ,
49177	 => std_logic_vector(to_unsigned(67,8) ,
49178	 => std_logic_vector(to_unsigned(58,8) ,
49179	 => std_logic_vector(to_unsigned(25,8) ,
49180	 => std_logic_vector(to_unsigned(49,8) ,
49181	 => std_logic_vector(to_unsigned(63,8) ,
49182	 => std_logic_vector(to_unsigned(59,8) ,
49183	 => std_logic_vector(to_unsigned(33,8) ,
49184	 => std_logic_vector(to_unsigned(35,8) ,
49185	 => std_logic_vector(to_unsigned(41,8) ,
49186	 => std_logic_vector(to_unsigned(35,8) ,
49187	 => std_logic_vector(to_unsigned(39,8) ,
49188	 => std_logic_vector(to_unsigned(45,8) ,
49189	 => std_logic_vector(to_unsigned(43,8) ,
49190	 => std_logic_vector(to_unsigned(48,8) ,
49191	 => std_logic_vector(to_unsigned(52,8) ,
49192	 => std_logic_vector(to_unsigned(52,8) ,
49193	 => std_logic_vector(to_unsigned(47,8) ,
49194	 => std_logic_vector(to_unsigned(44,8) ,
49195	 => std_logic_vector(to_unsigned(38,8) ,
49196	 => std_logic_vector(to_unsigned(39,8) ,
49197	 => std_logic_vector(to_unsigned(40,8) ,
49198	 => std_logic_vector(to_unsigned(35,8) ,
49199	 => std_logic_vector(to_unsigned(38,8) ,
49200	 => std_logic_vector(to_unsigned(37,8) ,
49201	 => std_logic_vector(to_unsigned(20,8) ,
49202	 => std_logic_vector(to_unsigned(22,8) ,
49203	 => std_logic_vector(to_unsigned(38,8) ,
49204	 => std_logic_vector(to_unsigned(37,8) ,
49205	 => std_logic_vector(to_unsigned(33,8) ,
49206	 => std_logic_vector(to_unsigned(34,8) ,
49207	 => std_logic_vector(to_unsigned(42,8) ,
49208	 => std_logic_vector(to_unsigned(58,8) ,
49209	 => std_logic_vector(to_unsigned(76,8) ,
49210	 => std_logic_vector(to_unsigned(69,8) ,
49211	 => std_logic_vector(to_unsigned(8,8) ,
49212	 => std_logic_vector(to_unsigned(1,8) ,
49213	 => std_logic_vector(to_unsigned(5,8) ,
49214	 => std_logic_vector(to_unsigned(96,8) ,
49215	 => std_logic_vector(to_unsigned(82,8) ,
49216	 => std_logic_vector(to_unsigned(104,8) ,
49217	 => std_logic_vector(to_unsigned(146,8) ,
49218	 => std_logic_vector(to_unsigned(142,8) ,
49219	 => std_logic_vector(to_unsigned(121,8) ,
49220	 => std_logic_vector(to_unsigned(111,8) ,
49221	 => std_logic_vector(to_unsigned(70,8) ,
49222	 => std_logic_vector(to_unsigned(93,8) ,
49223	 => std_logic_vector(to_unsigned(63,8) ,
49224	 => std_logic_vector(to_unsigned(87,8) ,
49225	 => std_logic_vector(to_unsigned(64,8) ,
49226	 => std_logic_vector(to_unsigned(131,8) ,
49227	 => std_logic_vector(to_unsigned(130,8) ,
49228	 => std_logic_vector(to_unsigned(101,8) ,
49229	 => std_logic_vector(to_unsigned(61,8) ,
49230	 => std_logic_vector(to_unsigned(32,8) ,
49231	 => std_logic_vector(to_unsigned(34,8) ,
49232	 => std_logic_vector(to_unsigned(34,8) ,
49233	 => std_logic_vector(to_unsigned(37,8) ,
49234	 => std_logic_vector(to_unsigned(36,8) ,
49235	 => std_logic_vector(to_unsigned(7,8) ,
49236	 => std_logic_vector(to_unsigned(1,8) ,
49237	 => std_logic_vector(to_unsigned(1,8) ,
49238	 => std_logic_vector(to_unsigned(2,8) ,
49239	 => std_logic_vector(to_unsigned(6,8) ,
49240	 => std_logic_vector(to_unsigned(9,8) ,
49241	 => std_logic_vector(to_unsigned(4,8) ,
49242	 => std_logic_vector(to_unsigned(1,8) ,
49243	 => std_logic_vector(to_unsigned(1,8) ,
49244	 => std_logic_vector(to_unsigned(0,8) ,
49245	 => std_logic_vector(to_unsigned(1,8) ,
49246	 => std_logic_vector(to_unsigned(5,8) ,
49247	 => std_logic_vector(to_unsigned(9,8) ,
49248	 => std_logic_vector(to_unsigned(32,8) ,
49249	 => std_logic_vector(to_unsigned(37,8) ,
49250	 => std_logic_vector(to_unsigned(35,8) ,
49251	 => std_logic_vector(to_unsigned(43,8) ,
49252	 => std_logic_vector(to_unsigned(43,8) ,
49253	 => std_logic_vector(to_unsigned(56,8) ,
49254	 => std_logic_vector(to_unsigned(63,8) ,
49255	 => std_logic_vector(to_unsigned(47,8) ,
49256	 => std_logic_vector(to_unsigned(35,8) ,
49257	 => std_logic_vector(to_unsigned(37,8) ,
49258	 => std_logic_vector(to_unsigned(38,8) ,
49259	 => std_logic_vector(to_unsigned(38,8) ,
49260	 => std_logic_vector(to_unsigned(32,8) ,
49261	 => std_logic_vector(to_unsigned(41,8) ,
49262	 => std_logic_vector(to_unsigned(67,8) ,
49263	 => std_logic_vector(to_unsigned(26,8) ,
49264	 => std_logic_vector(to_unsigned(27,8) ,
49265	 => std_logic_vector(to_unsigned(35,8) ,
49266	 => std_logic_vector(to_unsigned(29,8) ,
49267	 => std_logic_vector(to_unsigned(19,8) ,
49268	 => std_logic_vector(to_unsigned(48,8) ,
49269	 => std_logic_vector(to_unsigned(80,8) ,
49270	 => std_logic_vector(to_unsigned(66,8) ,
49271	 => std_logic_vector(to_unsigned(35,8) ,
49272	 => std_logic_vector(to_unsigned(35,8) ,
49273	 => std_logic_vector(to_unsigned(47,8) ,
49274	 => std_logic_vector(to_unsigned(54,8) ,
49275	 => std_logic_vector(to_unsigned(47,8) ,
49276	 => std_logic_vector(to_unsigned(51,8) ,
49277	 => std_logic_vector(to_unsigned(37,8) ,
49278	 => std_logic_vector(to_unsigned(13,8) ,
49279	 => std_logic_vector(to_unsigned(31,8) ,
49280	 => std_logic_vector(to_unsigned(58,8) ,
49281	 => std_logic_vector(to_unsigned(95,8) ,
49282	 => std_logic_vector(to_unsigned(95,8) ,
49283	 => std_logic_vector(to_unsigned(96,8) ,
49284	 => std_logic_vector(to_unsigned(90,8) ,
49285	 => std_logic_vector(to_unsigned(79,8) ,
49286	 => std_logic_vector(to_unsigned(77,8) ,
49287	 => std_logic_vector(to_unsigned(81,8) ,
49288	 => std_logic_vector(to_unsigned(81,8) ,
49289	 => std_logic_vector(to_unsigned(72,8) ,
49290	 => std_logic_vector(to_unsigned(55,8) ,
49291	 => std_logic_vector(to_unsigned(51,8) ,
49292	 => std_logic_vector(to_unsigned(46,8) ,
49293	 => std_logic_vector(to_unsigned(48,8) ,
49294	 => std_logic_vector(to_unsigned(44,8) ,
49295	 => std_logic_vector(to_unsigned(48,8) ,
49296	 => std_logic_vector(to_unsigned(90,8) ,
49297	 => std_logic_vector(to_unsigned(111,8) ,
49298	 => std_logic_vector(to_unsigned(101,8) ,
49299	 => std_logic_vector(to_unsigned(101,8) ,
49300	 => std_logic_vector(to_unsigned(99,8) ,
49301	 => std_logic_vector(to_unsigned(107,8) ,
49302	 => std_logic_vector(to_unsigned(107,8) ,
49303	 => std_logic_vector(to_unsigned(96,8) ,
49304	 => std_logic_vector(to_unsigned(101,8) ,
49305	 => std_logic_vector(to_unsigned(91,8) ,
49306	 => std_logic_vector(to_unsigned(88,8) ,
49307	 => std_logic_vector(to_unsigned(84,8) ,
49308	 => std_logic_vector(to_unsigned(85,8) ,
49309	 => std_logic_vector(to_unsigned(96,8) ,
49310	 => std_logic_vector(to_unsigned(97,8) ,
49311	 => std_logic_vector(to_unsigned(92,8) ,
49312	 => std_logic_vector(to_unsigned(99,8) ,
49313	 => std_logic_vector(to_unsigned(99,8) ,
49314	 => std_logic_vector(to_unsigned(121,8) ,
49315	 => std_logic_vector(to_unsigned(97,8) ,
49316	 => std_logic_vector(to_unsigned(73,8) ,
49317	 => std_logic_vector(to_unsigned(52,8) ,
49318	 => std_logic_vector(to_unsigned(48,8) ,
49319	 => std_logic_vector(to_unsigned(54,8) ,
49320	 => std_logic_vector(to_unsigned(57,8) ,
49321	 => std_logic_vector(to_unsigned(56,8) ,
49322	 => std_logic_vector(to_unsigned(109,8) ,
49323	 => std_logic_vector(to_unsigned(131,8) ,
49324	 => std_logic_vector(to_unsigned(95,8) ,
49325	 => std_logic_vector(to_unsigned(76,8) ,
49326	 => std_logic_vector(to_unsigned(66,8) ,
49327	 => std_logic_vector(to_unsigned(56,8) ,
49328	 => std_logic_vector(to_unsigned(82,8) ,
49329	 => std_logic_vector(to_unsigned(103,8) ,
49330	 => std_logic_vector(to_unsigned(103,8) ,
49331	 => std_logic_vector(to_unsigned(86,8) ,
49332	 => std_logic_vector(to_unsigned(65,8) ,
49333	 => std_logic_vector(to_unsigned(67,8) ,
49334	 => std_logic_vector(to_unsigned(76,8) ,
49335	 => std_logic_vector(to_unsigned(97,8) ,
49336	 => std_logic_vector(to_unsigned(100,8) ,
49337	 => std_logic_vector(to_unsigned(65,8) ,
49338	 => std_logic_vector(to_unsigned(45,8) ,
49339	 => std_logic_vector(to_unsigned(62,8) ,
49340	 => std_logic_vector(to_unsigned(109,8) ,
49341	 => std_logic_vector(to_unsigned(122,8) ,
49342	 => std_logic_vector(to_unsigned(115,8) ,
49343	 => std_logic_vector(to_unsigned(79,8) ,
49344	 => std_logic_vector(to_unsigned(93,8) ,
49345	 => std_logic_vector(to_unsigned(100,8) ,
49346	 => std_logic_vector(to_unsigned(78,8) ,
49347	 => std_logic_vector(to_unsigned(74,8) ,
49348	 => std_logic_vector(to_unsigned(71,8) ,
49349	 => std_logic_vector(to_unsigned(60,8) ,
49350	 => std_logic_vector(to_unsigned(88,8) ,
49351	 => std_logic_vector(to_unsigned(119,8) ,
49352	 => std_logic_vector(to_unsigned(116,8) ,
49353	 => std_logic_vector(to_unsigned(116,8) ,
49354	 => std_logic_vector(to_unsigned(116,8) ,
49355	 => std_logic_vector(to_unsigned(91,8) ,
49356	 => std_logic_vector(to_unsigned(54,8) ,
49357	 => std_logic_vector(to_unsigned(57,8) ,
49358	 => std_logic_vector(to_unsigned(69,8) ,
49359	 => std_logic_vector(to_unsigned(55,8) ,
49360	 => std_logic_vector(to_unsigned(66,8) ,
49361	 => std_logic_vector(to_unsigned(76,8) ,
49362	 => std_logic_vector(to_unsigned(72,8) ,
49363	 => std_logic_vector(to_unsigned(70,8) ,
49364	 => std_logic_vector(to_unsigned(57,8) ,
49365	 => std_logic_vector(to_unsigned(64,8) ,
49366	 => std_logic_vector(to_unsigned(67,8) ,
49367	 => std_logic_vector(to_unsigned(50,8) ,
49368	 => std_logic_vector(to_unsigned(45,8) ,
49369	 => std_logic_vector(to_unsigned(41,8) ,
49370	 => std_logic_vector(to_unsigned(42,8) ,
49371	 => std_logic_vector(to_unsigned(43,8) ,
49372	 => std_logic_vector(to_unsigned(40,8) ,
49373	 => std_logic_vector(to_unsigned(42,8) ,
49374	 => std_logic_vector(to_unsigned(39,8) ,
49375	 => std_logic_vector(to_unsigned(44,8) ,
49376	 => std_logic_vector(to_unsigned(42,8) ,
49377	 => std_logic_vector(to_unsigned(42,8) ,
49378	 => std_logic_vector(to_unsigned(47,8) ,
49379	 => std_logic_vector(to_unsigned(46,8) ,
49380	 => std_logic_vector(to_unsigned(52,8) ,
49381	 => std_logic_vector(to_unsigned(63,8) ,
49382	 => std_logic_vector(to_unsigned(53,8) ,
49383	 => std_logic_vector(to_unsigned(45,8) ,
49384	 => std_logic_vector(to_unsigned(96,8) ,
49385	 => std_logic_vector(to_unsigned(136,8) ,
49386	 => std_logic_vector(to_unsigned(121,8) ,
49387	 => std_logic_vector(to_unsigned(116,8) ,
49388	 => std_logic_vector(to_unsigned(115,8) ,
49389	 => std_logic_vector(to_unsigned(105,8) ,
49390	 => std_logic_vector(to_unsigned(99,8) ,
49391	 => std_logic_vector(to_unsigned(109,8) ,
49392	 => std_logic_vector(to_unsigned(81,8) ,
49393	 => std_logic_vector(to_unsigned(57,8) ,
49394	 => std_logic_vector(to_unsigned(66,8) ,
49395	 => std_logic_vector(to_unsigned(79,8) ,
49396	 => std_logic_vector(to_unsigned(91,8) ,
49397	 => std_logic_vector(to_unsigned(100,8) ,
49398	 => std_logic_vector(to_unsigned(90,8) ,
49399	 => std_logic_vector(to_unsigned(58,8) ,
49400	 => std_logic_vector(to_unsigned(52,8) ,
49401	 => std_logic_vector(to_unsigned(73,8) ,
49402	 => std_logic_vector(to_unsigned(88,8) ,
49403	 => std_logic_vector(to_unsigned(80,8) ,
49404	 => std_logic_vector(to_unsigned(72,8) ,
49405	 => std_logic_vector(to_unsigned(66,8) ,
49406	 => std_logic_vector(to_unsigned(64,8) ,
49407	 => std_logic_vector(to_unsigned(84,8) ,
49408	 => std_logic_vector(to_unsigned(100,8) ,
49409	 => std_logic_vector(to_unsigned(72,8) ,
49410	 => std_logic_vector(to_unsigned(51,8) ,
49411	 => std_logic_vector(to_unsigned(59,8) ,
49412	 => std_logic_vector(to_unsigned(65,8) ,
49413	 => std_logic_vector(to_unsigned(42,8) ,
49414	 => std_logic_vector(to_unsigned(52,8) ,
49415	 => std_logic_vector(to_unsigned(45,8) ,
49416	 => std_logic_vector(to_unsigned(21,8) ,
49417	 => std_logic_vector(to_unsigned(14,8) ,
49418	 => std_logic_vector(to_unsigned(17,8) ,
49419	 => std_logic_vector(to_unsigned(19,8) ,
49420	 => std_logic_vector(to_unsigned(32,8) ,
49421	 => std_logic_vector(to_unsigned(69,8) ,
49422	 => std_logic_vector(to_unsigned(84,8) ,
49423	 => std_logic_vector(to_unsigned(37,8) ,
49424	 => std_logic_vector(to_unsigned(63,8) ,
49425	 => std_logic_vector(to_unsigned(85,8) ,
49426	 => std_logic_vector(to_unsigned(61,8) ,
49427	 => std_logic_vector(to_unsigned(33,8) ,
49428	 => std_logic_vector(to_unsigned(19,8) ,
49429	 => std_logic_vector(to_unsigned(25,8) ,
49430	 => std_logic_vector(to_unsigned(51,8) ,
49431	 => std_logic_vector(to_unsigned(56,8) ,
49432	 => std_logic_vector(to_unsigned(45,8) ,
49433	 => std_logic_vector(to_unsigned(47,8) ,
49434	 => std_logic_vector(to_unsigned(32,8) ,
49435	 => std_logic_vector(to_unsigned(13,8) ,
49436	 => std_logic_vector(to_unsigned(23,8) ,
49437	 => std_logic_vector(to_unsigned(48,8) ,
49438	 => std_logic_vector(to_unsigned(74,8) ,
49439	 => std_logic_vector(to_unsigned(51,8) ,
49440	 => std_logic_vector(to_unsigned(32,8) ,
49441	 => std_logic_vector(to_unsigned(19,8) ,
49442	 => std_logic_vector(to_unsigned(29,8) ,
49443	 => std_logic_vector(to_unsigned(32,8) ,
49444	 => std_logic_vector(to_unsigned(25,8) ,
49445	 => std_logic_vector(to_unsigned(27,8) ,
49446	 => std_logic_vector(to_unsigned(24,8) ,
49447	 => std_logic_vector(to_unsigned(15,8) ,
49448	 => std_logic_vector(to_unsigned(12,8) ,
49449	 => std_logic_vector(to_unsigned(22,8) ,
49450	 => std_logic_vector(to_unsigned(25,8) ,
49451	 => std_logic_vector(to_unsigned(23,8) ,
49452	 => std_logic_vector(to_unsigned(22,8) ,
49453	 => std_logic_vector(to_unsigned(20,8) ,
49454	 => std_logic_vector(to_unsigned(22,8) ,
49455	 => std_logic_vector(to_unsigned(30,8) ,
49456	 => std_logic_vector(to_unsigned(38,8) ,
49457	 => std_logic_vector(to_unsigned(66,8) ,
49458	 => std_logic_vector(to_unsigned(73,8) ,
49459	 => std_logic_vector(to_unsigned(50,8) ,
49460	 => std_logic_vector(to_unsigned(49,8) ,
49461	 => std_logic_vector(to_unsigned(62,8) ,
49462	 => std_logic_vector(to_unsigned(57,8) ,
49463	 => std_logic_vector(to_unsigned(55,8) ,
49464	 => std_logic_vector(to_unsigned(61,8) ,
49465	 => std_logic_vector(to_unsigned(47,8) ,
49466	 => std_logic_vector(to_unsigned(25,8) ,
49467	 => std_logic_vector(to_unsigned(37,8) ,
49468	 => std_logic_vector(to_unsigned(17,8) ,
49469	 => std_logic_vector(to_unsigned(11,8) ,
49470	 => std_logic_vector(to_unsigned(35,8) ,
49471	 => std_logic_vector(to_unsigned(37,8) ,
49472	 => std_logic_vector(to_unsigned(24,8) ,
49473	 => std_logic_vector(to_unsigned(19,8) ,
49474	 => std_logic_vector(to_unsigned(25,8) ,
49475	 => std_logic_vector(to_unsigned(37,8) ,
49476	 => std_logic_vector(to_unsigned(27,8) ,
49477	 => std_logic_vector(to_unsigned(31,8) ,
49478	 => std_logic_vector(to_unsigned(45,8) ,
49479	 => std_logic_vector(to_unsigned(37,8) ,
49480	 => std_logic_vector(to_unsigned(32,8) ,
49481	 => std_logic_vector(to_unsigned(42,8) ,
49482	 => std_logic_vector(to_unsigned(48,8) ,
49483	 => std_logic_vector(to_unsigned(46,8) ,
49484	 => std_logic_vector(to_unsigned(40,8) ,
49485	 => std_logic_vector(to_unsigned(41,8) ,
49486	 => std_logic_vector(to_unsigned(30,8) ,
49487	 => std_logic_vector(to_unsigned(32,8) ,
49488	 => std_logic_vector(to_unsigned(46,8) ,
49489	 => std_logic_vector(to_unsigned(45,8) ,
49490	 => std_logic_vector(to_unsigned(30,8) ,
49491	 => std_logic_vector(to_unsigned(26,8) ,
49492	 => std_logic_vector(to_unsigned(21,8) ,
49493	 => std_logic_vector(to_unsigned(21,8) ,
49494	 => std_logic_vector(to_unsigned(25,8) ,
49495	 => std_logic_vector(to_unsigned(17,8) ,
49496	 => std_logic_vector(to_unsigned(17,8) ,
49497	 => std_logic_vector(to_unsigned(45,8) ,
49498	 => std_logic_vector(to_unsigned(45,8) ,
49499	 => std_logic_vector(to_unsigned(31,8) ,
49500	 => std_logic_vector(to_unsigned(45,8) ,
49501	 => std_logic_vector(to_unsigned(47,8) ,
49502	 => std_logic_vector(to_unsigned(47,8) ,
49503	 => std_logic_vector(to_unsigned(35,8) ,
49504	 => std_logic_vector(to_unsigned(35,8) ,
49505	 => std_logic_vector(to_unsigned(46,8) ,
49506	 => std_logic_vector(to_unsigned(41,8) ,
49507	 => std_logic_vector(to_unsigned(35,8) ,
49508	 => std_logic_vector(to_unsigned(48,8) ,
49509	 => std_logic_vector(to_unsigned(35,8) ,
49510	 => std_logic_vector(to_unsigned(42,8) ,
49511	 => std_logic_vector(to_unsigned(45,8) ,
49512	 => std_logic_vector(to_unsigned(46,8) ,
49513	 => std_logic_vector(to_unsigned(44,8) ,
49514	 => std_logic_vector(to_unsigned(32,8) ,
49515	 => std_logic_vector(to_unsigned(34,8) ,
49516	 => std_logic_vector(to_unsigned(43,8) ,
49517	 => std_logic_vector(to_unsigned(41,8) ,
49518	 => std_logic_vector(to_unsigned(37,8) ,
49519	 => std_logic_vector(to_unsigned(41,8) ,
49520	 => std_logic_vector(to_unsigned(39,8) ,
49521	 => std_logic_vector(to_unsigned(20,8) ,
49522	 => std_logic_vector(to_unsigned(20,8) ,
49523	 => std_logic_vector(to_unsigned(35,8) ,
49524	 => std_logic_vector(to_unsigned(35,8) ,
49525	 => std_logic_vector(to_unsigned(40,8) ,
49526	 => std_logic_vector(to_unsigned(47,8) ,
49527	 => std_logic_vector(to_unsigned(51,8) ,
49528	 => std_logic_vector(to_unsigned(58,8) ,
49529	 => std_logic_vector(to_unsigned(25,8) ,
49530	 => std_logic_vector(to_unsigned(74,8) ,
49531	 => std_logic_vector(to_unsigned(36,8) ,
49532	 => std_logic_vector(to_unsigned(0,8) ,
49533	 => std_logic_vector(to_unsigned(2,8) ,
49534	 => std_logic_vector(to_unsigned(36,8) ,
49535	 => std_logic_vector(to_unsigned(93,8) ,
49536	 => std_logic_vector(to_unsigned(108,8) ,
49537	 => std_logic_vector(to_unsigned(87,8) ,
49538	 => std_logic_vector(to_unsigned(104,8) ,
49539	 => std_logic_vector(to_unsigned(70,8) ,
49540	 => std_logic_vector(to_unsigned(93,8) ,
49541	 => std_logic_vector(to_unsigned(77,8) ,
49542	 => std_logic_vector(to_unsigned(96,8) ,
49543	 => std_logic_vector(to_unsigned(71,8) ,
49544	 => std_logic_vector(to_unsigned(84,8) ,
49545	 => std_logic_vector(to_unsigned(56,8) ,
49546	 => std_logic_vector(to_unsigned(125,8) ,
49547	 => std_logic_vector(to_unsigned(130,8) ,
49548	 => std_logic_vector(to_unsigned(114,8) ,
49549	 => std_logic_vector(to_unsigned(61,8) ,
49550	 => std_logic_vector(to_unsigned(37,8) ,
49551	 => std_logic_vector(to_unsigned(45,8) ,
49552	 => std_logic_vector(to_unsigned(33,8) ,
49553	 => std_logic_vector(to_unsigned(25,8) ,
49554	 => std_logic_vector(to_unsigned(22,8) ,
49555	 => std_logic_vector(to_unsigned(3,8) ,
49556	 => std_logic_vector(to_unsigned(2,8) ,
49557	 => std_logic_vector(to_unsigned(4,8) ,
49558	 => std_logic_vector(to_unsigned(2,8) ,
49559	 => std_logic_vector(to_unsigned(7,8) ,
49560	 => std_logic_vector(to_unsigned(22,8) ,
49561	 => std_logic_vector(to_unsigned(13,8) ,
49562	 => std_logic_vector(to_unsigned(2,8) ,
49563	 => std_logic_vector(to_unsigned(2,8) ,
49564	 => std_logic_vector(to_unsigned(3,8) ,
49565	 => std_logic_vector(to_unsigned(3,8) ,
49566	 => std_logic_vector(to_unsigned(8,8) ,
49567	 => std_logic_vector(to_unsigned(22,8) ,
49568	 => std_logic_vector(to_unsigned(15,8) ,
49569	 => std_logic_vector(to_unsigned(5,8) ,
49570	 => std_logic_vector(to_unsigned(12,8) ,
49571	 => std_logic_vector(to_unsigned(30,8) ,
49572	 => std_logic_vector(to_unsigned(42,8) ,
49573	 => std_logic_vector(to_unsigned(58,8) ,
49574	 => std_logic_vector(to_unsigned(50,8) ,
49575	 => std_logic_vector(to_unsigned(33,8) ,
49576	 => std_logic_vector(to_unsigned(24,8) ,
49577	 => std_logic_vector(to_unsigned(23,8) ,
49578	 => std_logic_vector(to_unsigned(17,8) ,
49579	 => std_logic_vector(to_unsigned(38,8) ,
49580	 => std_logic_vector(to_unsigned(65,8) ,
49581	 => std_logic_vector(to_unsigned(55,8) ,
49582	 => std_logic_vector(to_unsigned(46,8) ,
49583	 => std_logic_vector(to_unsigned(25,8) ,
49584	 => std_logic_vector(to_unsigned(20,8) ,
49585	 => std_logic_vector(to_unsigned(28,8) ,
49586	 => std_logic_vector(to_unsigned(24,8) ,
49587	 => std_logic_vector(to_unsigned(18,8) ,
49588	 => std_logic_vector(to_unsigned(45,8) ,
49589	 => std_logic_vector(to_unsigned(60,8) ,
49590	 => std_logic_vector(to_unsigned(77,8) ,
49591	 => std_logic_vector(to_unsigned(109,8) ,
49592	 => std_logic_vector(to_unsigned(112,8) ,
49593	 => std_logic_vector(to_unsigned(86,8) ,
49594	 => std_logic_vector(to_unsigned(82,8) ,
49595	 => std_logic_vector(to_unsigned(71,8) ,
49596	 => std_logic_vector(to_unsigned(80,8) ,
49597	 => std_logic_vector(to_unsigned(96,8) ,
49598	 => std_logic_vector(to_unsigned(72,8) ,
49599	 => std_logic_vector(to_unsigned(71,8) ,
49600	 => std_logic_vector(to_unsigned(71,8) ,
49601	 => std_logic_vector(to_unsigned(97,8) ,
49602	 => std_logic_vector(to_unsigned(90,8) ,
49603	 => std_logic_vector(to_unsigned(88,8) ,
49604	 => std_logic_vector(to_unsigned(100,8) ,
49605	 => std_logic_vector(to_unsigned(105,8) ,
49606	 => std_logic_vector(to_unsigned(107,8) ,
49607	 => std_logic_vector(to_unsigned(93,8) ,
49608	 => std_logic_vector(to_unsigned(85,8) ,
49609	 => std_logic_vector(to_unsigned(81,8) ,
49610	 => std_logic_vector(to_unsigned(63,8) ,
49611	 => std_logic_vector(to_unsigned(52,8) ,
49612	 => std_logic_vector(to_unsigned(52,8) ,
49613	 => std_logic_vector(to_unsigned(54,8) ,
49614	 => std_logic_vector(to_unsigned(49,8) ,
49615	 => std_logic_vector(to_unsigned(66,8) ,
49616	 => std_logic_vector(to_unsigned(112,8) ,
49617	 => std_logic_vector(to_unsigned(125,8) ,
49618	 => std_logic_vector(to_unsigned(111,8) ,
49619	 => std_logic_vector(to_unsigned(111,8) ,
49620	 => std_logic_vector(to_unsigned(105,8) ,
49621	 => std_logic_vector(to_unsigned(115,8) ,
49622	 => std_logic_vector(to_unsigned(107,8) ,
49623	 => std_logic_vector(to_unsigned(93,8) ,
49624	 => std_logic_vector(to_unsigned(97,8) ,
49625	 => std_logic_vector(to_unsigned(93,8) ,
49626	 => std_logic_vector(to_unsigned(92,8) ,
49627	 => std_logic_vector(to_unsigned(99,8) ,
49628	 => std_logic_vector(to_unsigned(97,8) ,
49629	 => std_logic_vector(to_unsigned(99,8) ,
49630	 => std_logic_vector(to_unsigned(93,8) ,
49631	 => std_logic_vector(to_unsigned(84,8) ,
49632	 => std_logic_vector(to_unsigned(88,8) ,
49633	 => std_logic_vector(to_unsigned(91,8) ,
49634	 => std_logic_vector(to_unsigned(97,8) ,
49635	 => std_logic_vector(to_unsigned(78,8) ,
49636	 => std_logic_vector(to_unsigned(63,8) ,
49637	 => std_logic_vector(to_unsigned(60,8) ,
49638	 => std_logic_vector(to_unsigned(71,8) ,
49639	 => std_logic_vector(to_unsigned(68,8) ,
49640	 => std_logic_vector(to_unsigned(70,8) ,
49641	 => std_logic_vector(to_unsigned(78,8) ,
49642	 => std_logic_vector(to_unsigned(86,8) ,
49643	 => std_logic_vector(to_unsigned(100,8) ,
49644	 => std_logic_vector(to_unsigned(79,8) ,
49645	 => std_logic_vector(to_unsigned(77,8) ,
49646	 => std_logic_vector(to_unsigned(70,8) ,
49647	 => std_logic_vector(to_unsigned(49,8) ,
49648	 => std_logic_vector(to_unsigned(62,8) ,
49649	 => std_logic_vector(to_unsigned(80,8) ,
49650	 => std_logic_vector(to_unsigned(101,8) ,
49651	 => std_logic_vector(to_unsigned(72,8) ,
49652	 => std_logic_vector(to_unsigned(39,8) ,
49653	 => std_logic_vector(to_unsigned(66,8) ,
49654	 => std_logic_vector(to_unsigned(81,8) ,
49655	 => std_logic_vector(to_unsigned(76,8) ,
49656	 => std_logic_vector(to_unsigned(82,8) ,
49657	 => std_logic_vector(to_unsigned(76,8) ,
49658	 => std_logic_vector(to_unsigned(81,8) ,
49659	 => std_logic_vector(to_unsigned(91,8) ,
49660	 => std_logic_vector(to_unsigned(92,8) ,
49661	 => std_logic_vector(to_unsigned(95,8) ,
49662	 => std_logic_vector(to_unsigned(85,8) ,
49663	 => std_logic_vector(to_unsigned(70,8) ,
49664	 => std_logic_vector(to_unsigned(82,8) ,
49665	 => std_logic_vector(to_unsigned(81,8) ,
49666	 => std_logic_vector(to_unsigned(67,8) ,
49667	 => std_logic_vector(to_unsigned(58,8) ,
49668	 => std_logic_vector(to_unsigned(60,8) ,
49669	 => std_logic_vector(to_unsigned(58,8) ,
49670	 => std_logic_vector(to_unsigned(63,8) ,
49671	 => std_logic_vector(to_unsigned(68,8) ,
49672	 => std_logic_vector(to_unsigned(84,8) ,
49673	 => std_logic_vector(to_unsigned(97,8) ,
49674	 => std_logic_vector(to_unsigned(103,8) ,
49675	 => std_logic_vector(to_unsigned(46,8) ,
49676	 => std_logic_vector(to_unsigned(35,8) ,
49677	 => std_logic_vector(to_unsigned(88,8) ,
49678	 => std_logic_vector(to_unsigned(88,8) ,
49679	 => std_logic_vector(to_unsigned(76,8) ,
49680	 => std_logic_vector(to_unsigned(70,8) ,
49681	 => std_logic_vector(to_unsigned(59,8) ,
49682	 => std_logic_vector(to_unsigned(50,8) ,
49683	 => std_logic_vector(to_unsigned(58,8) ,
49684	 => std_logic_vector(to_unsigned(65,8) ,
49685	 => std_logic_vector(to_unsigned(65,8) ,
49686	 => std_logic_vector(to_unsigned(61,8) ,
49687	 => std_logic_vector(to_unsigned(50,8) ,
49688	 => std_logic_vector(to_unsigned(45,8) ,
49689	 => std_logic_vector(to_unsigned(41,8) ,
49690	 => std_logic_vector(to_unsigned(37,8) ,
49691	 => std_logic_vector(to_unsigned(41,8) ,
49692	 => std_logic_vector(to_unsigned(42,8) ,
49693	 => std_logic_vector(to_unsigned(44,8) ,
49694	 => std_logic_vector(to_unsigned(40,8) ,
49695	 => std_logic_vector(to_unsigned(40,8) ,
49696	 => std_logic_vector(to_unsigned(34,8) ,
49697	 => std_logic_vector(to_unsigned(35,8) ,
49698	 => std_logic_vector(to_unsigned(37,8) ,
49699	 => std_logic_vector(to_unsigned(39,8) ,
49700	 => std_logic_vector(to_unsigned(36,8) ,
49701	 => std_logic_vector(to_unsigned(41,8) ,
49702	 => std_logic_vector(to_unsigned(42,8) ,
49703	 => std_logic_vector(to_unsigned(41,8) ,
49704	 => std_logic_vector(to_unsigned(86,8) ,
49705	 => std_logic_vector(to_unsigned(100,8) ,
49706	 => std_logic_vector(to_unsigned(92,8) ,
49707	 => std_logic_vector(to_unsigned(107,8) ,
49708	 => std_logic_vector(to_unsigned(112,8) ,
49709	 => std_logic_vector(to_unsigned(118,8) ,
49710	 => std_logic_vector(to_unsigned(119,8) ,
49711	 => std_logic_vector(to_unsigned(118,8) ,
49712	 => std_logic_vector(to_unsigned(111,8) ,
49713	 => std_logic_vector(to_unsigned(111,8) ,
49714	 => std_logic_vector(to_unsigned(115,8) ,
49715	 => std_logic_vector(to_unsigned(111,8) ,
49716	 => std_logic_vector(to_unsigned(103,8) ,
49717	 => std_logic_vector(to_unsigned(105,8) ,
49718	 => std_logic_vector(to_unsigned(73,8) ,
49719	 => std_logic_vector(to_unsigned(29,8) ,
49720	 => std_logic_vector(to_unsigned(60,8) ,
49721	 => std_logic_vector(to_unsigned(90,8) ,
49722	 => std_logic_vector(to_unsigned(91,8) ,
49723	 => std_logic_vector(to_unsigned(96,8) ,
49724	 => std_logic_vector(to_unsigned(93,8) ,
49725	 => std_logic_vector(to_unsigned(92,8) ,
49726	 => std_logic_vector(to_unsigned(107,8) ,
49727	 => std_logic_vector(to_unsigned(100,8) ,
49728	 => std_logic_vector(to_unsigned(76,8) ,
49729	 => std_logic_vector(to_unsigned(62,8) ,
49730	 => std_logic_vector(to_unsigned(45,8) ,
49731	 => std_logic_vector(to_unsigned(41,8) ,
49732	 => std_logic_vector(to_unsigned(58,8) ,
49733	 => std_logic_vector(to_unsigned(35,8) ,
49734	 => std_logic_vector(to_unsigned(45,8) ,
49735	 => std_logic_vector(to_unsigned(44,8) ,
49736	 => std_logic_vector(to_unsigned(19,8) ,
49737	 => std_logic_vector(to_unsigned(14,8) ,
49738	 => std_logic_vector(to_unsigned(20,8) ,
49739	 => std_logic_vector(to_unsigned(28,8) ,
49740	 => std_logic_vector(to_unsigned(29,8) ,
49741	 => std_logic_vector(to_unsigned(72,8) ,
49742	 => std_logic_vector(to_unsigned(84,8) ,
49743	 => std_logic_vector(to_unsigned(17,8) ,
49744	 => std_logic_vector(to_unsigned(43,8) ,
49745	 => std_logic_vector(to_unsigned(112,8) ,
49746	 => std_logic_vector(to_unsigned(62,8) ,
49747	 => std_logic_vector(to_unsigned(32,8) ,
49748	 => std_logic_vector(to_unsigned(14,8) ,
49749	 => std_logic_vector(to_unsigned(32,8) ,
49750	 => std_logic_vector(to_unsigned(70,8) ,
49751	 => std_logic_vector(to_unsigned(45,8) ,
49752	 => std_logic_vector(to_unsigned(51,8) ,
49753	 => std_logic_vector(to_unsigned(45,8) ,
49754	 => std_logic_vector(to_unsigned(43,8) ,
49755	 => std_logic_vector(to_unsigned(32,8) ,
49756	 => std_logic_vector(to_unsigned(47,8) ,
49757	 => std_logic_vector(to_unsigned(62,8) ,
49758	 => std_logic_vector(to_unsigned(43,8) ,
49759	 => std_logic_vector(to_unsigned(24,8) ,
49760	 => std_logic_vector(to_unsigned(23,8) ,
49761	 => std_logic_vector(to_unsigned(26,8) ,
49762	 => std_logic_vector(to_unsigned(41,8) ,
49763	 => std_logic_vector(to_unsigned(41,8) ,
49764	 => std_logic_vector(to_unsigned(35,8) ,
49765	 => std_logic_vector(to_unsigned(40,8) ,
49766	 => std_logic_vector(to_unsigned(36,8) ,
49767	 => std_logic_vector(to_unsigned(26,8) ,
49768	 => std_logic_vector(to_unsigned(19,8) ,
49769	 => std_logic_vector(to_unsigned(46,8) ,
49770	 => std_logic_vector(to_unsigned(51,8) ,
49771	 => std_logic_vector(to_unsigned(30,8) ,
49772	 => std_logic_vector(to_unsigned(17,8) ,
49773	 => std_logic_vector(to_unsigned(17,8) ,
49774	 => std_logic_vector(to_unsigned(20,8) ,
49775	 => std_logic_vector(to_unsigned(19,8) ,
49776	 => std_logic_vector(to_unsigned(16,8) ,
49777	 => std_logic_vector(to_unsigned(44,8) ,
49778	 => std_logic_vector(to_unsigned(59,8) ,
49779	 => std_logic_vector(to_unsigned(57,8) ,
49780	 => std_logic_vector(to_unsigned(55,8) ,
49781	 => std_logic_vector(to_unsigned(62,8) ,
49782	 => std_logic_vector(to_unsigned(56,8) ,
49783	 => std_logic_vector(to_unsigned(51,8) ,
49784	 => std_logic_vector(to_unsigned(60,8) ,
49785	 => std_logic_vector(to_unsigned(45,8) ,
49786	 => std_logic_vector(to_unsigned(41,8) ,
49787	 => std_logic_vector(to_unsigned(32,8) ,
49788	 => std_logic_vector(to_unsigned(17,8) ,
49789	 => std_logic_vector(to_unsigned(19,8) ,
49790	 => std_logic_vector(to_unsigned(35,8) ,
49791	 => std_logic_vector(to_unsigned(32,8) ,
49792	 => std_logic_vector(to_unsigned(28,8) ,
49793	 => std_logic_vector(to_unsigned(29,8) ,
49794	 => std_logic_vector(to_unsigned(32,8) ,
49795	 => std_logic_vector(to_unsigned(43,8) ,
49796	 => std_logic_vector(to_unsigned(36,8) ,
49797	 => std_logic_vector(to_unsigned(37,8) ,
49798	 => std_logic_vector(to_unsigned(42,8) ,
49799	 => std_logic_vector(to_unsigned(46,8) ,
49800	 => std_logic_vector(to_unsigned(56,8) ,
49801	 => std_logic_vector(to_unsigned(48,8) ,
49802	 => std_logic_vector(to_unsigned(40,8) ,
49803	 => std_logic_vector(to_unsigned(41,8) ,
49804	 => std_logic_vector(to_unsigned(44,8) ,
49805	 => std_logic_vector(to_unsigned(41,8) ,
49806	 => std_logic_vector(to_unsigned(12,8) ,
49807	 => std_logic_vector(to_unsigned(11,8) ,
49808	 => std_logic_vector(to_unsigned(17,8) ,
49809	 => std_logic_vector(to_unsigned(23,8) ,
49810	 => std_logic_vector(to_unsigned(38,8) ,
49811	 => std_logic_vector(to_unsigned(42,8) ,
49812	 => std_logic_vector(to_unsigned(40,8) ,
49813	 => std_logic_vector(to_unsigned(34,8) ,
49814	 => std_logic_vector(to_unsigned(30,8) ,
49815	 => std_logic_vector(to_unsigned(24,8) ,
49816	 => std_logic_vector(to_unsigned(30,8) ,
49817	 => std_logic_vector(to_unsigned(39,8) ,
49818	 => std_logic_vector(to_unsigned(45,8) ,
49819	 => std_logic_vector(to_unsigned(34,8) ,
49820	 => std_logic_vector(to_unsigned(38,8) ,
49821	 => std_logic_vector(to_unsigned(48,8) ,
49822	 => std_logic_vector(to_unsigned(42,8) ,
49823	 => std_logic_vector(to_unsigned(28,8) ,
49824	 => std_logic_vector(to_unsigned(28,8) ,
49825	 => std_logic_vector(to_unsigned(38,8) ,
49826	 => std_logic_vector(to_unsigned(37,8) ,
49827	 => std_logic_vector(to_unsigned(30,8) ,
49828	 => std_logic_vector(to_unsigned(38,8) ,
49829	 => std_logic_vector(to_unsigned(34,8) ,
49830	 => std_logic_vector(to_unsigned(37,8) ,
49831	 => std_logic_vector(to_unsigned(42,8) ,
49832	 => std_logic_vector(to_unsigned(42,8) ,
49833	 => std_logic_vector(to_unsigned(38,8) ,
49834	 => std_logic_vector(to_unsigned(27,8) ,
49835	 => std_logic_vector(to_unsigned(33,8) ,
49836	 => std_logic_vector(to_unsigned(41,8) ,
49837	 => std_logic_vector(to_unsigned(31,8) ,
49838	 => std_logic_vector(to_unsigned(35,8) ,
49839	 => std_logic_vector(to_unsigned(35,8) ,
49840	 => std_logic_vector(to_unsigned(28,8) ,
49841	 => std_logic_vector(to_unsigned(19,8) ,
49842	 => std_logic_vector(to_unsigned(22,8) ,
49843	 => std_logic_vector(to_unsigned(30,8) ,
49844	 => std_logic_vector(to_unsigned(32,8) ,
49845	 => std_logic_vector(to_unsigned(37,8) ,
49846	 => std_logic_vector(to_unsigned(51,8) ,
49847	 => std_logic_vector(to_unsigned(62,8) ,
49848	 => std_logic_vector(to_unsigned(50,8) ,
49849	 => std_logic_vector(to_unsigned(28,8) ,
49850	 => std_logic_vector(to_unsigned(91,8) ,
49851	 => std_logic_vector(to_unsigned(79,8) ,
49852	 => std_logic_vector(to_unsigned(3,8) ,
49853	 => std_logic_vector(to_unsigned(0,8) ,
49854	 => std_logic_vector(to_unsigned(4,8) ,
49855	 => std_logic_vector(to_unsigned(56,8) ,
49856	 => std_logic_vector(to_unsigned(118,8) ,
49857	 => std_logic_vector(to_unsigned(71,8) ,
49858	 => std_logic_vector(to_unsigned(99,8) ,
49859	 => std_logic_vector(to_unsigned(63,8) ,
49860	 => std_logic_vector(to_unsigned(100,8) ,
49861	 => std_logic_vector(to_unsigned(86,8) ,
49862	 => std_logic_vector(to_unsigned(92,8) ,
49863	 => std_logic_vector(to_unsigned(78,8) ,
49864	 => std_logic_vector(to_unsigned(84,8) ,
49865	 => std_logic_vector(to_unsigned(56,8) ,
49866	 => std_logic_vector(to_unsigned(122,8) ,
49867	 => std_logic_vector(to_unsigned(127,8) ,
49868	 => std_logic_vector(to_unsigned(108,8) ,
49869	 => std_logic_vector(to_unsigned(41,8) ,
49870	 => std_logic_vector(to_unsigned(22,8) ,
49871	 => std_logic_vector(to_unsigned(33,8) ,
49872	 => std_logic_vector(to_unsigned(33,8) ,
49873	 => std_logic_vector(to_unsigned(30,8) ,
49874	 => std_logic_vector(to_unsigned(29,8) ,
49875	 => std_logic_vector(to_unsigned(23,8) ,
49876	 => std_logic_vector(to_unsigned(5,8) ,
49877	 => std_logic_vector(to_unsigned(1,8) ,
49878	 => std_logic_vector(to_unsigned(2,8) ,
49879	 => std_logic_vector(to_unsigned(3,8) ,
49880	 => std_logic_vector(to_unsigned(4,8) ,
49881	 => std_logic_vector(to_unsigned(2,8) ,
49882	 => std_logic_vector(to_unsigned(2,8) ,
49883	 => std_logic_vector(to_unsigned(5,8) ,
49884	 => std_logic_vector(to_unsigned(20,8) ,
49885	 => std_logic_vector(to_unsigned(36,8) ,
49886	 => std_logic_vector(to_unsigned(39,8) ,
49887	 => std_logic_vector(to_unsigned(38,8) ,
49888	 => std_logic_vector(to_unsigned(20,8) ,
49889	 => std_logic_vector(to_unsigned(16,8) ,
49890	 => std_logic_vector(to_unsigned(19,8) ,
49891	 => std_logic_vector(to_unsigned(22,8) ,
49892	 => std_logic_vector(to_unsigned(37,8) ,
49893	 => std_logic_vector(to_unsigned(50,8) ,
49894	 => std_logic_vector(to_unsigned(45,8) ,
49895	 => std_logic_vector(to_unsigned(26,8) ,
49896	 => std_logic_vector(to_unsigned(15,8) ,
49897	 => std_logic_vector(to_unsigned(13,8) ,
49898	 => std_logic_vector(to_unsigned(27,8) ,
49899	 => std_logic_vector(to_unsigned(26,8) ,
49900	 => std_logic_vector(to_unsigned(23,8) ,
49901	 => std_logic_vector(to_unsigned(29,8) ,
49902	 => std_logic_vector(to_unsigned(13,8) ,
49903	 => std_logic_vector(to_unsigned(11,8) ,
49904	 => std_logic_vector(to_unsigned(16,8) ,
49905	 => std_logic_vector(to_unsigned(32,8) ,
49906	 => std_logic_vector(to_unsigned(26,8) ,
49907	 => std_logic_vector(to_unsigned(18,8) ,
49908	 => std_logic_vector(to_unsigned(41,8) ,
49909	 => std_logic_vector(to_unsigned(32,8) ,
49910	 => std_logic_vector(to_unsigned(51,8) ,
49911	 => std_logic_vector(to_unsigned(72,8) ,
49912	 => std_logic_vector(to_unsigned(84,8) ,
49913	 => std_logic_vector(to_unsigned(61,8) ,
49914	 => std_logic_vector(to_unsigned(51,8) ,
49915	 => std_logic_vector(to_unsigned(27,8) ,
49916	 => std_logic_vector(to_unsigned(69,8) ,
49917	 => std_logic_vector(to_unsigned(163,8) ,
49918	 => std_logic_vector(to_unsigned(159,8) ,
49919	 => std_logic_vector(to_unsigned(104,8) ,
49920	 => std_logic_vector(to_unsigned(56,8) ,
49921	 => std_logic_vector(to_unsigned(104,8) ,
49922	 => std_logic_vector(to_unsigned(107,8) ,
49923	 => std_logic_vector(to_unsigned(116,8) ,
49924	 => std_logic_vector(to_unsigned(114,8) ,
49925	 => std_logic_vector(to_unsigned(93,8) ,
49926	 => std_logic_vector(to_unsigned(88,8) ,
49927	 => std_logic_vector(to_unsigned(103,8) ,
49928	 => std_logic_vector(to_unsigned(124,8) ,
49929	 => std_logic_vector(to_unsigned(134,8) ,
49930	 => std_logic_vector(to_unsigned(82,8) ,
49931	 => std_logic_vector(to_unsigned(48,8) ,
49932	 => std_logic_vector(to_unsigned(57,8) ,
49933	 => std_logic_vector(to_unsigned(54,8) ,
49934	 => std_logic_vector(to_unsigned(58,8) ,
49935	 => std_logic_vector(to_unsigned(77,8) ,
49936	 => std_logic_vector(to_unsigned(111,8) ,
49937	 => std_logic_vector(to_unsigned(122,8) ,
49938	 => std_logic_vector(to_unsigned(118,8) ,
49939	 => std_logic_vector(to_unsigned(127,8) ,
49940	 => std_logic_vector(to_unsigned(118,8) ,
49941	 => std_logic_vector(to_unsigned(121,8) ,
49942	 => std_logic_vector(to_unsigned(115,8) ,
49943	 => std_logic_vector(to_unsigned(88,8) ,
49944	 => std_logic_vector(to_unsigned(85,8) ,
49945	 => std_logic_vector(to_unsigned(90,8) ,
49946	 => std_logic_vector(to_unsigned(84,8) ,
49947	 => std_logic_vector(to_unsigned(92,8) ,
49948	 => std_logic_vector(to_unsigned(85,8) ,
49949	 => std_logic_vector(to_unsigned(77,8) ,
49950	 => std_logic_vector(to_unsigned(91,8) ,
49951	 => std_logic_vector(to_unsigned(87,8) ,
49952	 => std_logic_vector(to_unsigned(95,8) ,
49953	 => std_logic_vector(to_unsigned(101,8) ,
49954	 => std_logic_vector(to_unsigned(68,8) ,
49955	 => std_logic_vector(to_unsigned(33,8) ,
49956	 => std_logic_vector(to_unsigned(40,8) ,
49957	 => std_logic_vector(to_unsigned(44,8) ,
49958	 => std_logic_vector(to_unsigned(59,8) ,
49959	 => std_logic_vector(to_unsigned(47,8) ,
49960	 => std_logic_vector(to_unsigned(52,8) ,
49961	 => std_logic_vector(to_unsigned(96,8) ,
49962	 => std_logic_vector(to_unsigned(62,8) ,
49963	 => std_logic_vector(to_unsigned(55,8) ,
49964	 => std_logic_vector(to_unsigned(80,8) ,
49965	 => std_logic_vector(to_unsigned(100,8) ,
49966	 => std_logic_vector(to_unsigned(92,8) ,
49967	 => std_logic_vector(to_unsigned(58,8) ,
49968	 => std_logic_vector(to_unsigned(58,8) ,
49969	 => std_logic_vector(to_unsigned(86,8) ,
49970	 => std_logic_vector(to_unsigned(103,8) ,
49971	 => std_logic_vector(to_unsigned(73,8) ,
49972	 => std_logic_vector(to_unsigned(57,8) ,
49973	 => std_logic_vector(to_unsigned(67,8) ,
49974	 => std_logic_vector(to_unsigned(73,8) ,
49975	 => std_logic_vector(to_unsigned(68,8) ,
49976	 => std_logic_vector(to_unsigned(79,8) ,
49977	 => std_logic_vector(to_unsigned(90,8) ,
49978	 => std_logic_vector(to_unsigned(91,8) ,
49979	 => std_logic_vector(to_unsigned(92,8) ,
49980	 => std_logic_vector(to_unsigned(72,8) ,
49981	 => std_logic_vector(to_unsigned(76,8) ,
49982	 => std_logic_vector(to_unsigned(74,8) ,
49983	 => std_logic_vector(to_unsigned(68,8) ,
49984	 => std_logic_vector(to_unsigned(77,8) ,
49985	 => std_logic_vector(to_unsigned(77,8) ,
49986	 => std_logic_vector(to_unsigned(86,8) ,
49987	 => std_logic_vector(to_unsigned(79,8) ,
49988	 => std_logic_vector(to_unsigned(41,8) ,
49989	 => std_logic_vector(to_unsigned(56,8) ,
49990	 => std_logic_vector(to_unsigned(70,8) ,
49991	 => std_logic_vector(to_unsigned(53,8) ,
49992	 => std_logic_vector(to_unsigned(67,8) ,
49993	 => std_logic_vector(to_unsigned(65,8) ,
49994	 => std_logic_vector(to_unsigned(50,8) ,
49995	 => std_logic_vector(to_unsigned(36,8) ,
49996	 => std_logic_vector(to_unsigned(67,8) ,
49997	 => std_logic_vector(to_unsigned(124,8) ,
49998	 => std_logic_vector(to_unsigned(109,8) ,
49999	 => std_logic_vector(to_unsigned(63,8) ,
50000	 => std_logic_vector(to_unsigned(66,8) ,
50001	 => std_logic_vector(to_unsigned(63,8) ,
50002	 => std_logic_vector(to_unsigned(54,8) ,
50003	 => std_logic_vector(to_unsigned(62,8) ,
50004	 => std_logic_vector(to_unsigned(57,8) ,
50005	 => std_logic_vector(to_unsigned(58,8) ,
50006	 => std_logic_vector(to_unsigned(59,8) ,
50007	 => std_logic_vector(to_unsigned(53,8) ,
50008	 => std_logic_vector(to_unsigned(46,8) ,
50009	 => std_logic_vector(to_unsigned(49,8) ,
50010	 => std_logic_vector(to_unsigned(42,8) ,
50011	 => std_logic_vector(to_unsigned(36,8) ,
50012	 => std_logic_vector(to_unsigned(41,8) ,
50013	 => std_logic_vector(to_unsigned(45,8) ,
50014	 => std_logic_vector(to_unsigned(35,8) ,
50015	 => std_logic_vector(to_unsigned(34,8) ,
50016	 => std_logic_vector(to_unsigned(41,8) ,
50017	 => std_logic_vector(to_unsigned(38,8) ,
50018	 => std_logic_vector(to_unsigned(38,8) ,
50019	 => std_logic_vector(to_unsigned(41,8) ,
50020	 => std_logic_vector(to_unsigned(45,8) ,
50021	 => std_logic_vector(to_unsigned(51,8) ,
50022	 => std_logic_vector(to_unsigned(40,8) ,
50023	 => std_logic_vector(to_unsigned(45,8) ,
50024	 => std_logic_vector(to_unsigned(85,8) ,
50025	 => std_logic_vector(to_unsigned(76,8) ,
50026	 => std_logic_vector(to_unsigned(62,8) ,
50027	 => std_logic_vector(to_unsigned(61,8) ,
50028	 => std_logic_vector(to_unsigned(74,8) ,
50029	 => std_logic_vector(to_unsigned(69,8) ,
50030	 => std_logic_vector(to_unsigned(66,8) ,
50031	 => std_logic_vector(to_unsigned(71,8) ,
50032	 => std_logic_vector(to_unsigned(73,8) ,
50033	 => std_logic_vector(to_unsigned(86,8) ,
50034	 => std_logic_vector(to_unsigned(95,8) ,
50035	 => std_logic_vector(to_unsigned(105,8) ,
50036	 => std_logic_vector(to_unsigned(103,8) ,
50037	 => std_logic_vector(to_unsigned(105,8) ,
50038	 => std_logic_vector(to_unsigned(66,8) ,
50039	 => std_logic_vector(to_unsigned(25,8) ,
50040	 => std_logic_vector(to_unsigned(65,8) ,
50041	 => std_logic_vector(to_unsigned(82,8) ,
50042	 => std_logic_vector(to_unsigned(79,8) ,
50043	 => std_logic_vector(to_unsigned(77,8) ,
50044	 => std_logic_vector(to_unsigned(88,8) ,
50045	 => std_logic_vector(to_unsigned(111,8) ,
50046	 => std_logic_vector(to_unsigned(90,8) ,
50047	 => std_logic_vector(to_unsigned(59,8) ,
50048	 => std_logic_vector(to_unsigned(45,8) ,
50049	 => std_logic_vector(to_unsigned(58,8) ,
50050	 => std_logic_vector(to_unsigned(50,8) ,
50051	 => std_logic_vector(to_unsigned(45,8) ,
50052	 => std_logic_vector(to_unsigned(59,8) ,
50053	 => std_logic_vector(to_unsigned(37,8) ,
50054	 => std_logic_vector(to_unsigned(39,8) ,
50055	 => std_logic_vector(to_unsigned(41,8) ,
50056	 => std_logic_vector(to_unsigned(22,8) ,
50057	 => std_logic_vector(to_unsigned(16,8) ,
50058	 => std_logic_vector(to_unsigned(17,8) ,
50059	 => std_logic_vector(to_unsigned(17,8) ,
50060	 => std_logic_vector(to_unsigned(24,8) ,
50061	 => std_logic_vector(to_unsigned(58,8) ,
50062	 => std_logic_vector(to_unsigned(85,8) ,
50063	 => std_logic_vector(to_unsigned(35,8) ,
50064	 => std_logic_vector(to_unsigned(55,8) ,
50065	 => std_logic_vector(to_unsigned(103,8) ,
50066	 => std_logic_vector(to_unsigned(59,8) ,
50067	 => std_logic_vector(to_unsigned(23,8) ,
50068	 => std_logic_vector(to_unsigned(10,8) ,
50069	 => std_logic_vector(to_unsigned(33,8) ,
50070	 => std_logic_vector(to_unsigned(80,8) ,
50071	 => std_logic_vector(to_unsigned(60,8) ,
50072	 => std_logic_vector(to_unsigned(80,8) ,
50073	 => std_logic_vector(to_unsigned(56,8) ,
50074	 => std_logic_vector(to_unsigned(67,8) ,
50075	 => std_logic_vector(to_unsigned(46,8) ,
50076	 => std_logic_vector(to_unsigned(86,8) ,
50077	 => std_logic_vector(to_unsigned(71,8) ,
50078	 => std_logic_vector(to_unsigned(32,8) ,
50079	 => std_logic_vector(to_unsigned(24,8) ,
50080	 => std_logic_vector(to_unsigned(14,8) ,
50081	 => std_logic_vector(to_unsigned(39,8) ,
50082	 => std_logic_vector(to_unsigned(48,8) ,
50083	 => std_logic_vector(to_unsigned(35,8) ,
50084	 => std_logic_vector(to_unsigned(34,8) ,
50085	 => std_logic_vector(to_unsigned(30,8) ,
50086	 => std_logic_vector(to_unsigned(42,8) ,
50087	 => std_logic_vector(to_unsigned(36,8) ,
50088	 => std_logic_vector(to_unsigned(22,8) ,
50089	 => std_logic_vector(to_unsigned(45,8) ,
50090	 => std_logic_vector(to_unsigned(34,8) ,
50091	 => std_logic_vector(to_unsigned(22,8) ,
50092	 => std_logic_vector(to_unsigned(19,8) ,
50093	 => std_logic_vector(to_unsigned(20,8) ,
50094	 => std_logic_vector(to_unsigned(30,8) ,
50095	 => std_logic_vector(to_unsigned(35,8) ,
50096	 => std_logic_vector(to_unsigned(20,8) ,
50097	 => std_logic_vector(to_unsigned(30,8) ,
50098	 => std_logic_vector(to_unsigned(43,8) ,
50099	 => std_logic_vector(to_unsigned(69,8) ,
50100	 => std_logic_vector(to_unsigned(56,8) ,
50101	 => std_logic_vector(to_unsigned(57,8) ,
50102	 => std_logic_vector(to_unsigned(58,8) ,
50103	 => std_logic_vector(to_unsigned(45,8) ,
50104	 => std_logic_vector(to_unsigned(38,8) ,
50105	 => std_logic_vector(to_unsigned(46,8) ,
50106	 => std_logic_vector(to_unsigned(38,8) ,
50107	 => std_logic_vector(to_unsigned(31,8) ,
50108	 => std_logic_vector(to_unsigned(20,8) ,
50109	 => std_logic_vector(to_unsigned(24,8) ,
50110	 => std_logic_vector(to_unsigned(39,8) ,
50111	 => std_logic_vector(to_unsigned(31,8) ,
50112	 => std_logic_vector(to_unsigned(17,8) ,
50113	 => std_logic_vector(to_unsigned(16,8) ,
50114	 => std_logic_vector(to_unsigned(24,8) ,
50115	 => std_logic_vector(to_unsigned(23,8) ,
50116	 => std_logic_vector(to_unsigned(15,8) ,
50117	 => std_logic_vector(to_unsigned(25,8) ,
50118	 => std_logic_vector(to_unsigned(37,8) ,
50119	 => std_logic_vector(to_unsigned(53,8) ,
50120	 => std_logic_vector(to_unsigned(90,8) ,
50121	 => std_logic_vector(to_unsigned(77,8) ,
50122	 => std_logic_vector(to_unsigned(40,8) ,
50123	 => std_logic_vector(to_unsigned(37,8) ,
50124	 => std_logic_vector(to_unsigned(43,8) ,
50125	 => std_logic_vector(to_unsigned(33,8) ,
50126	 => std_logic_vector(to_unsigned(37,8) ,
50127	 => std_logic_vector(to_unsigned(33,8) ,
50128	 => std_logic_vector(to_unsigned(25,8) ,
50129	 => std_logic_vector(to_unsigned(31,8) ,
50130	 => std_logic_vector(to_unsigned(34,8) ,
50131	 => std_logic_vector(to_unsigned(40,8) ,
50132	 => std_logic_vector(to_unsigned(35,8) ,
50133	 => std_logic_vector(to_unsigned(32,8) ,
50134	 => std_logic_vector(to_unsigned(24,8) ,
50135	 => std_logic_vector(to_unsigned(22,8) ,
50136	 => std_logic_vector(to_unsigned(29,8) ,
50137	 => std_logic_vector(to_unsigned(32,8) ,
50138	 => std_logic_vector(to_unsigned(39,8) ,
50139	 => std_logic_vector(to_unsigned(27,8) ,
50140	 => std_logic_vector(to_unsigned(30,8) ,
50141	 => std_logic_vector(to_unsigned(41,8) ,
50142	 => std_logic_vector(to_unsigned(30,8) ,
50143	 => std_logic_vector(to_unsigned(25,8) ,
50144	 => std_logic_vector(to_unsigned(26,8) ,
50145	 => std_logic_vector(to_unsigned(37,8) ,
50146	 => std_logic_vector(to_unsigned(34,8) ,
50147	 => std_logic_vector(to_unsigned(32,8) ,
50148	 => std_logic_vector(to_unsigned(37,8) ,
50149	 => std_logic_vector(to_unsigned(30,8) ,
50150	 => std_logic_vector(to_unsigned(35,8) ,
50151	 => std_logic_vector(to_unsigned(38,8) ,
50152	 => std_logic_vector(to_unsigned(32,8) ,
50153	 => std_logic_vector(to_unsigned(32,8) ,
50154	 => std_logic_vector(to_unsigned(47,8) ,
50155	 => std_logic_vector(to_unsigned(44,8) ,
50156	 => std_logic_vector(to_unsigned(29,8) ,
50157	 => std_logic_vector(to_unsigned(28,8) ,
50158	 => std_logic_vector(to_unsigned(25,8) ,
50159	 => std_logic_vector(to_unsigned(33,8) ,
50160	 => std_logic_vector(to_unsigned(42,8) ,
50161	 => std_logic_vector(to_unsigned(19,8) ,
50162	 => std_logic_vector(to_unsigned(14,8) ,
50163	 => std_logic_vector(to_unsigned(20,8) ,
50164	 => std_logic_vector(to_unsigned(36,8) ,
50165	 => std_logic_vector(to_unsigned(39,8) ,
50166	 => std_logic_vector(to_unsigned(42,8) ,
50167	 => std_logic_vector(to_unsigned(42,8) ,
50168	 => std_logic_vector(to_unsigned(24,8) ,
50169	 => std_logic_vector(to_unsigned(41,8) ,
50170	 => std_logic_vector(to_unsigned(87,8) ,
50171	 => std_logic_vector(to_unsigned(96,8) ,
50172	 => std_logic_vector(to_unsigned(37,8) ,
50173	 => std_logic_vector(to_unsigned(3,8) ,
50174	 => std_logic_vector(to_unsigned(0,8) ,
50175	 => std_logic_vector(to_unsigned(16,8) ,
50176	 => std_logic_vector(to_unsigned(119,8) ,
50177	 => std_logic_vector(to_unsigned(69,8) ,
50178	 => std_logic_vector(to_unsigned(100,8) ,
50179	 => std_logic_vector(to_unsigned(64,8) ,
50180	 => std_logic_vector(to_unsigned(85,8) ,
50181	 => std_logic_vector(to_unsigned(74,8) ,
50182	 => std_logic_vector(to_unsigned(86,8) ,
50183	 => std_logic_vector(to_unsigned(62,8) ,
50184	 => std_logic_vector(to_unsigned(97,8) ,
50185	 => std_logic_vector(to_unsigned(74,8) ,
50186	 => std_logic_vector(to_unsigned(122,8) ,
50187	 => std_logic_vector(to_unsigned(86,8) ,
50188	 => std_logic_vector(to_unsigned(41,8) ,
50189	 => std_logic_vector(to_unsigned(27,8) ,
50190	 => std_logic_vector(to_unsigned(23,8) ,
50191	 => std_logic_vector(to_unsigned(23,8) ,
50192	 => std_logic_vector(to_unsigned(28,8) ,
50193	 => std_logic_vector(to_unsigned(25,8) ,
50194	 => std_logic_vector(to_unsigned(17,8) ,
50195	 => std_logic_vector(to_unsigned(23,8) ,
50196	 => std_logic_vector(to_unsigned(12,8) ,
50197	 => std_logic_vector(to_unsigned(0,8) ,
50198	 => std_logic_vector(to_unsigned(0,8) ,
50199	 => std_logic_vector(to_unsigned(0,8) ,
50200	 => std_logic_vector(to_unsigned(0,8) ,
50201	 => std_logic_vector(to_unsigned(1,8) ,
50202	 => std_logic_vector(to_unsigned(6,8) ,
50203	 => std_logic_vector(to_unsigned(10,8) ,
50204	 => std_logic_vector(to_unsigned(16,8) ,
50205	 => std_logic_vector(to_unsigned(25,8) ,
50206	 => std_logic_vector(to_unsigned(30,8) ,
50207	 => std_logic_vector(to_unsigned(24,8) ,
50208	 => std_logic_vector(to_unsigned(25,8) ,
50209	 => std_logic_vector(to_unsigned(25,8) ,
50210	 => std_logic_vector(to_unsigned(27,8) ,
50211	 => std_logic_vector(to_unsigned(26,8) ,
50212	 => std_logic_vector(to_unsigned(30,8) ,
50213	 => std_logic_vector(to_unsigned(45,8) ,
50214	 => std_logic_vector(to_unsigned(39,8) ,
50215	 => std_logic_vector(to_unsigned(19,8) ,
50216	 => std_logic_vector(to_unsigned(13,8) ,
50217	 => std_logic_vector(to_unsigned(20,8) ,
50218	 => std_logic_vector(to_unsigned(29,8) ,
50219	 => std_logic_vector(to_unsigned(16,8) ,
50220	 => std_logic_vector(to_unsigned(20,8) ,
50221	 => std_logic_vector(to_unsigned(27,8) ,
50222	 => std_logic_vector(to_unsigned(25,8) ,
50223	 => std_logic_vector(to_unsigned(18,8) ,
50224	 => std_logic_vector(to_unsigned(10,8) ,
50225	 => std_logic_vector(to_unsigned(27,8) ,
50226	 => std_logic_vector(to_unsigned(22,8) ,
50227	 => std_logic_vector(to_unsigned(17,8) ,
50228	 => std_logic_vector(to_unsigned(50,8) ,
50229	 => std_logic_vector(to_unsigned(47,8) ,
50230	 => std_logic_vector(to_unsigned(45,8) ,
50231	 => std_logic_vector(to_unsigned(37,8) ,
50232	 => std_logic_vector(to_unsigned(49,8) ,
50233	 => std_logic_vector(to_unsigned(42,8) ,
50234	 => std_logic_vector(to_unsigned(47,8) ,
50235	 => std_logic_vector(to_unsigned(45,8) ,
50236	 => std_logic_vector(to_unsigned(60,8) ,
50237	 => std_logic_vector(to_unsigned(71,8) ,
50238	 => std_logic_vector(to_unsigned(78,8) ,
50239	 => std_logic_vector(to_unsigned(68,8) ,
50240	 => std_logic_vector(to_unsigned(20,8) ,
50241	 => std_logic_vector(to_unsigned(112,8) ,
50242	 => std_logic_vector(to_unsigned(108,8) ,
50243	 => std_logic_vector(to_unsigned(100,8) ,
50244	 => std_logic_vector(to_unsigned(87,8) ,
50245	 => std_logic_vector(to_unsigned(78,8) ,
50246	 => std_logic_vector(to_unsigned(86,8) ,
50247	 => std_logic_vector(to_unsigned(109,8) ,
50248	 => std_logic_vector(to_unsigned(131,8) ,
50249	 => std_logic_vector(to_unsigned(139,8) ,
50250	 => std_logic_vector(to_unsigned(81,8) ,
50251	 => std_logic_vector(to_unsigned(49,8) ,
50252	 => std_logic_vector(to_unsigned(58,8) ,
50253	 => std_logic_vector(to_unsigned(57,8) ,
50254	 => std_logic_vector(to_unsigned(71,8) ,
50255	 => std_logic_vector(to_unsigned(87,8) ,
50256	 => std_logic_vector(to_unsigned(96,8) ,
50257	 => std_logic_vector(to_unsigned(108,8) ,
50258	 => std_logic_vector(to_unsigned(125,8) ,
50259	 => std_logic_vector(to_unsigned(128,8) ,
50260	 => std_logic_vector(to_unsigned(124,8) ,
50261	 => std_logic_vector(to_unsigned(118,8) ,
50262	 => std_logic_vector(to_unsigned(105,8) ,
50263	 => std_logic_vector(to_unsigned(91,8) ,
50264	 => std_logic_vector(to_unsigned(87,8) ,
50265	 => std_logic_vector(to_unsigned(85,8) ,
50266	 => std_logic_vector(to_unsigned(86,8) ,
50267	 => std_logic_vector(to_unsigned(96,8) ,
50268	 => std_logic_vector(to_unsigned(86,8) ,
50269	 => std_logic_vector(to_unsigned(74,8) ,
50270	 => std_logic_vector(to_unsigned(90,8) ,
50271	 => std_logic_vector(to_unsigned(90,8) ,
50272	 => std_logic_vector(to_unsigned(88,8) ,
50273	 => std_logic_vector(to_unsigned(97,8) ,
50274	 => std_logic_vector(to_unsigned(73,8) ,
50275	 => std_logic_vector(to_unsigned(35,8) ,
50276	 => std_logic_vector(to_unsigned(33,8) ,
50277	 => std_logic_vector(to_unsigned(25,8) ,
50278	 => std_logic_vector(to_unsigned(24,8) ,
50279	 => std_logic_vector(to_unsigned(53,8) ,
50280	 => std_logic_vector(to_unsigned(80,8) ,
50281	 => std_logic_vector(to_unsigned(70,8) ,
50282	 => std_logic_vector(to_unsigned(43,8) ,
50283	 => std_logic_vector(to_unsigned(45,8) ,
50284	 => std_logic_vector(to_unsigned(64,8) ,
50285	 => std_logic_vector(to_unsigned(92,8) ,
50286	 => std_logic_vector(to_unsigned(130,8) ,
50287	 => std_logic_vector(to_unsigned(125,8) ,
50288	 => std_logic_vector(to_unsigned(134,8) ,
50289	 => std_logic_vector(to_unsigned(159,8) ,
50290	 => std_logic_vector(to_unsigned(130,8) ,
50291	 => std_logic_vector(to_unsigned(79,8) ,
50292	 => std_logic_vector(to_unsigned(78,8) ,
50293	 => std_logic_vector(to_unsigned(88,8) ,
50294	 => std_logic_vector(to_unsigned(85,8) ,
50295	 => std_logic_vector(to_unsigned(76,8) ,
50296	 => std_logic_vector(to_unsigned(77,8) ,
50297	 => std_logic_vector(to_unsigned(63,8) ,
50298	 => std_logic_vector(to_unsigned(70,8) ,
50299	 => std_logic_vector(to_unsigned(82,8) ,
50300	 => std_logic_vector(to_unsigned(70,8) ,
50301	 => std_logic_vector(to_unsigned(60,8) ,
50302	 => std_logic_vector(to_unsigned(66,8) ,
50303	 => std_logic_vector(to_unsigned(63,8) ,
50304	 => std_logic_vector(to_unsigned(77,8) ,
50305	 => std_logic_vector(to_unsigned(73,8) ,
50306	 => std_logic_vector(to_unsigned(79,8) ,
50307	 => std_logic_vector(to_unsigned(82,8) ,
50308	 => std_logic_vector(to_unsigned(80,8) ,
50309	 => std_logic_vector(to_unsigned(104,8) ,
50310	 => std_logic_vector(to_unsigned(101,8) ,
50311	 => std_logic_vector(to_unsigned(67,8) ,
50312	 => std_logic_vector(to_unsigned(100,8) ,
50313	 => std_logic_vector(to_unsigned(105,8) ,
50314	 => std_logic_vector(to_unsigned(96,8) ,
50315	 => std_logic_vector(to_unsigned(108,8) ,
50316	 => std_logic_vector(to_unsigned(111,8) ,
50317	 => std_logic_vector(to_unsigned(112,8) ,
50318	 => std_logic_vector(to_unsigned(96,8) ,
50319	 => std_logic_vector(to_unsigned(59,8) ,
50320	 => std_logic_vector(to_unsigned(56,8) ,
50321	 => std_logic_vector(to_unsigned(67,8) ,
50322	 => std_logic_vector(to_unsigned(74,8) ,
50323	 => std_logic_vector(to_unsigned(62,8) ,
50324	 => std_logic_vector(to_unsigned(56,8) ,
50325	 => std_logic_vector(to_unsigned(55,8) ,
50326	 => std_logic_vector(to_unsigned(54,8) ,
50327	 => std_logic_vector(to_unsigned(48,8) ,
50328	 => std_logic_vector(to_unsigned(45,8) ,
50329	 => std_logic_vector(to_unsigned(41,8) ,
50330	 => std_logic_vector(to_unsigned(47,8) ,
50331	 => std_logic_vector(to_unsigned(40,8) ,
50332	 => std_logic_vector(to_unsigned(38,8) ,
50333	 => std_logic_vector(to_unsigned(40,8) ,
50334	 => std_logic_vector(to_unsigned(31,8) ,
50335	 => std_logic_vector(to_unsigned(35,8) ,
50336	 => std_logic_vector(to_unsigned(36,8) ,
50337	 => std_logic_vector(to_unsigned(35,8) ,
50338	 => std_logic_vector(to_unsigned(32,8) ,
50339	 => std_logic_vector(to_unsigned(37,8) ,
50340	 => std_logic_vector(to_unsigned(35,8) ,
50341	 => std_logic_vector(to_unsigned(42,8) ,
50342	 => std_logic_vector(to_unsigned(40,8) ,
50343	 => std_logic_vector(to_unsigned(44,8) ,
50344	 => std_logic_vector(to_unsigned(87,8) ,
50345	 => std_logic_vector(to_unsigned(78,8) ,
50346	 => std_logic_vector(to_unsigned(55,8) ,
50347	 => std_logic_vector(to_unsigned(58,8) ,
50348	 => std_logic_vector(to_unsigned(68,8) ,
50349	 => std_logic_vector(to_unsigned(60,8) ,
50350	 => std_logic_vector(to_unsigned(45,8) ,
50351	 => std_logic_vector(to_unsigned(51,8) ,
50352	 => std_logic_vector(to_unsigned(41,8) ,
50353	 => std_logic_vector(to_unsigned(43,8) ,
50354	 => std_logic_vector(to_unsigned(40,8) ,
50355	 => std_logic_vector(to_unsigned(55,8) ,
50356	 => std_logic_vector(to_unsigned(53,8) ,
50357	 => std_logic_vector(to_unsigned(65,8) ,
50358	 => std_logic_vector(to_unsigned(43,8) ,
50359	 => std_logic_vector(to_unsigned(22,8) ,
50360	 => std_logic_vector(to_unsigned(37,8) ,
50361	 => std_logic_vector(to_unsigned(50,8) ,
50362	 => std_logic_vector(to_unsigned(43,8) ,
50363	 => std_logic_vector(to_unsigned(41,8) ,
50364	 => std_logic_vector(to_unsigned(79,8) ,
50365	 => std_logic_vector(to_unsigned(85,8) ,
50366	 => std_logic_vector(to_unsigned(52,8) ,
50367	 => std_logic_vector(to_unsigned(45,8) ,
50368	 => std_logic_vector(to_unsigned(53,8) ,
50369	 => std_logic_vector(to_unsigned(57,8) ,
50370	 => std_logic_vector(to_unsigned(32,8) ,
50371	 => std_logic_vector(to_unsigned(36,8) ,
50372	 => std_logic_vector(to_unsigned(61,8) ,
50373	 => std_logic_vector(to_unsigned(43,8) ,
50374	 => std_logic_vector(to_unsigned(43,8) ,
50375	 => std_logic_vector(to_unsigned(35,8) ,
50376	 => std_logic_vector(to_unsigned(20,8) ,
50377	 => std_logic_vector(to_unsigned(14,8) ,
50378	 => std_logic_vector(to_unsigned(16,8) ,
50379	 => std_logic_vector(to_unsigned(18,8) ,
50380	 => std_logic_vector(to_unsigned(25,8) ,
50381	 => std_logic_vector(to_unsigned(58,8) ,
50382	 => std_logic_vector(to_unsigned(90,8) ,
50383	 => std_logic_vector(to_unsigned(45,8) ,
50384	 => std_logic_vector(to_unsigned(67,8) ,
50385	 => std_logic_vector(to_unsigned(103,8) ,
50386	 => std_logic_vector(to_unsigned(49,8) ,
50387	 => std_logic_vector(to_unsigned(17,8) ,
50388	 => std_logic_vector(to_unsigned(7,8) ,
50389	 => std_logic_vector(to_unsigned(30,8) ,
50390	 => std_logic_vector(to_unsigned(79,8) ,
50391	 => std_logic_vector(to_unsigned(50,8) ,
50392	 => std_logic_vector(to_unsigned(76,8) ,
50393	 => std_logic_vector(to_unsigned(49,8) ,
50394	 => std_logic_vector(to_unsigned(68,8) ,
50395	 => std_logic_vector(to_unsigned(58,8) ,
50396	 => std_logic_vector(to_unsigned(87,8) ,
50397	 => std_logic_vector(to_unsigned(65,8) ,
50398	 => std_logic_vector(to_unsigned(29,8) ,
50399	 => std_logic_vector(to_unsigned(15,8) ,
50400	 => std_logic_vector(to_unsigned(13,8) ,
50401	 => std_logic_vector(to_unsigned(60,8) ,
50402	 => std_logic_vector(to_unsigned(50,8) ,
50403	 => std_logic_vector(to_unsigned(42,8) ,
50404	 => std_logic_vector(to_unsigned(45,8) ,
50405	 => std_logic_vector(to_unsigned(41,8) ,
50406	 => std_logic_vector(to_unsigned(28,8) ,
50407	 => std_logic_vector(to_unsigned(30,8) ,
50408	 => std_logic_vector(to_unsigned(47,8) ,
50409	 => std_logic_vector(to_unsigned(37,8) ,
50410	 => std_logic_vector(to_unsigned(20,8) ,
50411	 => std_logic_vector(to_unsigned(12,8) ,
50412	 => std_logic_vector(to_unsigned(14,8) ,
50413	 => std_logic_vector(to_unsigned(28,8) ,
50414	 => std_logic_vector(to_unsigned(32,8) ,
50415	 => std_logic_vector(to_unsigned(35,8) ,
50416	 => std_logic_vector(to_unsigned(25,8) ,
50417	 => std_logic_vector(to_unsigned(29,8) ,
50418	 => std_logic_vector(to_unsigned(41,8) ,
50419	 => std_logic_vector(to_unsigned(63,8) ,
50420	 => std_logic_vector(to_unsigned(63,8) ,
50421	 => std_logic_vector(to_unsigned(65,8) ,
50422	 => std_logic_vector(to_unsigned(69,8) ,
50423	 => std_logic_vector(to_unsigned(47,8) ,
50424	 => std_logic_vector(to_unsigned(30,8) ,
50425	 => std_logic_vector(to_unsigned(34,8) ,
50426	 => std_logic_vector(to_unsigned(32,8) ,
50427	 => std_logic_vector(to_unsigned(25,8) ,
50428	 => std_logic_vector(to_unsigned(17,8) ,
50429	 => std_logic_vector(to_unsigned(28,8) ,
50430	 => std_logic_vector(to_unsigned(40,8) ,
50431	 => std_logic_vector(to_unsigned(35,8) ,
50432	 => std_logic_vector(to_unsigned(32,8) ,
50433	 => std_logic_vector(to_unsigned(32,8) ,
50434	 => std_logic_vector(to_unsigned(33,8) ,
50435	 => std_logic_vector(to_unsigned(24,8) ,
50436	 => std_logic_vector(to_unsigned(24,8) ,
50437	 => std_logic_vector(to_unsigned(23,8) ,
50438	 => std_logic_vector(to_unsigned(29,8) ,
50439	 => std_logic_vector(to_unsigned(32,8) ,
50440	 => std_logic_vector(to_unsigned(43,8) ,
50441	 => std_logic_vector(to_unsigned(47,8) ,
50442	 => std_logic_vector(to_unsigned(37,8) ,
50443	 => std_logic_vector(to_unsigned(37,8) ,
50444	 => std_logic_vector(to_unsigned(41,8) ,
50445	 => std_logic_vector(to_unsigned(32,8) ,
50446	 => std_logic_vector(to_unsigned(56,8) ,
50447	 => std_logic_vector(to_unsigned(56,8) ,
50448	 => std_logic_vector(to_unsigned(70,8) ,
50449	 => std_logic_vector(to_unsigned(71,8) ,
50450	 => std_logic_vector(to_unsigned(25,8) ,
50451	 => std_logic_vector(to_unsigned(34,8) ,
50452	 => std_logic_vector(to_unsigned(29,8) ,
50453	 => std_logic_vector(to_unsigned(30,8) ,
50454	 => std_logic_vector(to_unsigned(53,8) ,
50455	 => std_logic_vector(to_unsigned(49,8) ,
50456	 => std_logic_vector(to_unsigned(35,8) ,
50457	 => std_logic_vector(to_unsigned(27,8) ,
50458	 => std_logic_vector(to_unsigned(36,8) ,
50459	 => std_logic_vector(to_unsigned(25,8) ,
50460	 => std_logic_vector(to_unsigned(29,8) ,
50461	 => std_logic_vector(to_unsigned(31,8) ,
50462	 => std_logic_vector(to_unsigned(25,8) ,
50463	 => std_logic_vector(to_unsigned(39,8) ,
50464	 => std_logic_vector(to_unsigned(29,8) ,
50465	 => std_logic_vector(to_unsigned(30,8) ,
50466	 => std_logic_vector(to_unsigned(27,8) ,
50467	 => std_logic_vector(to_unsigned(22,8) ,
50468	 => std_logic_vector(to_unsigned(26,8) ,
50469	 => std_logic_vector(to_unsigned(25,8) ,
50470	 => std_logic_vector(to_unsigned(30,8) ,
50471	 => std_logic_vector(to_unsigned(29,8) ,
50472	 => std_logic_vector(to_unsigned(28,8) ,
50473	 => std_logic_vector(to_unsigned(33,8) ,
50474	 => std_logic_vector(to_unsigned(45,8) ,
50475	 => std_logic_vector(to_unsigned(35,8) ,
50476	 => std_logic_vector(to_unsigned(25,8) ,
50477	 => std_logic_vector(to_unsigned(24,8) ,
50478	 => std_logic_vector(to_unsigned(19,8) ,
50479	 => std_logic_vector(to_unsigned(36,8) ,
50480	 => std_logic_vector(to_unsigned(49,8) ,
50481	 => std_logic_vector(to_unsigned(21,8) ,
50482	 => std_logic_vector(to_unsigned(17,8) ,
50483	 => std_logic_vector(to_unsigned(20,8) ,
50484	 => std_logic_vector(to_unsigned(41,8) ,
50485	 => std_logic_vector(to_unsigned(48,8) ,
50486	 => std_logic_vector(to_unsigned(30,8) ,
50487	 => std_logic_vector(to_unsigned(23,8) ,
50488	 => std_logic_vector(to_unsigned(25,8) ,
50489	 => std_logic_vector(to_unsigned(25,8) ,
50490	 => std_logic_vector(to_unsigned(81,8) ,
50491	 => std_logic_vector(to_unsigned(90,8) ,
50492	 => std_logic_vector(to_unsigned(90,8) ,
50493	 => std_logic_vector(to_unsigned(15,8) ,
50494	 => std_logic_vector(to_unsigned(0,8) ,
50495	 => std_logic_vector(to_unsigned(4,8) ,
50496	 => std_logic_vector(to_unsigned(63,8) ,
50497	 => std_logic_vector(to_unsigned(59,8) ,
50498	 => std_logic_vector(to_unsigned(88,8) ,
50499	 => std_logic_vector(to_unsigned(84,8) ,
50500	 => std_logic_vector(to_unsigned(91,8) ,
50501	 => std_logic_vector(to_unsigned(67,8) ,
50502	 => std_logic_vector(to_unsigned(92,8) ,
50503	 => std_logic_vector(to_unsigned(81,8) ,
50504	 => std_logic_vector(to_unsigned(95,8) ,
50505	 => std_logic_vector(to_unsigned(76,8) ,
50506	 => std_logic_vector(to_unsigned(101,8) ,
50507	 => std_logic_vector(to_unsigned(45,8) ,
50508	 => std_logic_vector(to_unsigned(30,8) ,
50509	 => std_logic_vector(to_unsigned(37,8) ,
50510	 => std_logic_vector(to_unsigned(23,8) ,
50511	 => std_logic_vector(to_unsigned(19,8) ,
50512	 => std_logic_vector(to_unsigned(42,8) ,
50513	 => std_logic_vector(to_unsigned(36,8) ,
50514	 => std_logic_vector(to_unsigned(19,8) ,
50515	 => std_logic_vector(to_unsigned(22,8) ,
50516	 => std_logic_vector(to_unsigned(12,8) ,
50517	 => std_logic_vector(to_unsigned(1,8) ,
50518	 => std_logic_vector(to_unsigned(0,8) ,
50519	 => std_logic_vector(to_unsigned(0,8) ,
50520	 => std_logic_vector(to_unsigned(0,8) ,
50521	 => std_logic_vector(to_unsigned(3,8) ,
50522	 => std_logic_vector(to_unsigned(42,8) ,
50523	 => std_logic_vector(to_unsigned(48,8) ,
50524	 => std_logic_vector(to_unsigned(23,8) ,
50525	 => std_logic_vector(to_unsigned(15,8) ,
50526	 => std_logic_vector(to_unsigned(24,8) ,
50527	 => std_logic_vector(to_unsigned(18,8) ,
50528	 => std_logic_vector(to_unsigned(13,8) ,
50529	 => std_logic_vector(to_unsigned(5,8) ,
50530	 => std_logic_vector(to_unsigned(7,8) ,
50531	 => std_logic_vector(to_unsigned(27,8) ,
50532	 => std_logic_vector(to_unsigned(30,8) ,
50533	 => std_logic_vector(to_unsigned(45,8) ,
50534	 => std_logic_vector(to_unsigned(35,8) ,
50535	 => std_logic_vector(to_unsigned(38,8) ,
50536	 => std_logic_vector(to_unsigned(27,8) ,
50537	 => std_logic_vector(to_unsigned(18,8) ,
50538	 => std_logic_vector(to_unsigned(23,8) ,
50539	 => std_logic_vector(to_unsigned(12,8) ,
50540	 => std_logic_vector(to_unsigned(24,8) ,
50541	 => std_logic_vector(to_unsigned(46,8) ,
50542	 => std_logic_vector(to_unsigned(44,8) ,
50543	 => std_logic_vector(to_unsigned(26,8) ,
50544	 => std_logic_vector(to_unsigned(12,8) ,
50545	 => std_logic_vector(to_unsigned(24,8) ,
50546	 => std_logic_vector(to_unsigned(17,8) ,
50547	 => std_logic_vector(to_unsigned(18,8) ,
50548	 => std_logic_vector(to_unsigned(35,8) ,
50549	 => std_logic_vector(to_unsigned(24,8) ,
50550	 => std_logic_vector(to_unsigned(31,8) ,
50551	 => std_logic_vector(to_unsigned(12,8) ,
50552	 => std_logic_vector(to_unsigned(17,8) ,
50553	 => std_logic_vector(to_unsigned(30,8) ,
50554	 => std_logic_vector(to_unsigned(36,8) ,
50555	 => std_logic_vector(to_unsigned(37,8) ,
50556	 => std_logic_vector(to_unsigned(55,8) ,
50557	 => std_logic_vector(to_unsigned(45,8) ,
50558	 => std_logic_vector(to_unsigned(45,8) ,
50559	 => std_logic_vector(to_unsigned(63,8) ,
50560	 => std_logic_vector(to_unsigned(43,8) ,
50561	 => std_logic_vector(to_unsigned(95,8) ,
50562	 => std_logic_vector(to_unsigned(91,8) ,
50563	 => std_logic_vector(to_unsigned(88,8) ,
50564	 => std_logic_vector(to_unsigned(108,8) ,
50565	 => std_logic_vector(to_unsigned(127,8) ,
50566	 => std_logic_vector(to_unsigned(130,8) ,
50567	 => std_logic_vector(to_unsigned(130,8) ,
50568	 => std_logic_vector(to_unsigned(104,8) ,
50569	 => std_logic_vector(to_unsigned(111,8) ,
50570	 => std_logic_vector(to_unsigned(97,8) ,
50571	 => std_logic_vector(to_unsigned(67,8) ,
50572	 => std_logic_vector(to_unsigned(71,8) ,
50573	 => std_logic_vector(to_unsigned(84,8) ,
50574	 => std_logic_vector(to_unsigned(92,8) ,
50575	 => std_logic_vector(to_unsigned(105,8) ,
50576	 => std_logic_vector(to_unsigned(112,8) ,
50577	 => std_logic_vector(to_unsigned(121,8) ,
50578	 => std_logic_vector(to_unsigned(122,8) ,
50579	 => std_logic_vector(to_unsigned(128,8) ,
50580	 => std_logic_vector(to_unsigned(121,8) ,
50581	 => std_logic_vector(to_unsigned(112,8) ,
50582	 => std_logic_vector(to_unsigned(109,8) ,
50583	 => std_logic_vector(to_unsigned(91,8) ,
50584	 => std_logic_vector(to_unsigned(67,8) ,
50585	 => std_logic_vector(to_unsigned(66,8) ,
50586	 => std_logic_vector(to_unsigned(69,8) ,
50587	 => std_logic_vector(to_unsigned(80,8) ,
50588	 => std_logic_vector(to_unsigned(81,8) ,
50589	 => std_logic_vector(to_unsigned(72,8) ,
50590	 => std_logic_vector(to_unsigned(84,8) ,
50591	 => std_logic_vector(to_unsigned(74,8) ,
50592	 => std_logic_vector(to_unsigned(87,8) ,
50593	 => std_logic_vector(to_unsigned(93,8) ,
50594	 => std_logic_vector(to_unsigned(68,8) ,
50595	 => std_logic_vector(to_unsigned(46,8) ,
50596	 => std_logic_vector(to_unsigned(50,8) ,
50597	 => std_logic_vector(to_unsigned(43,8) ,
50598	 => std_logic_vector(to_unsigned(41,8) ,
50599	 => std_logic_vector(to_unsigned(101,8) ,
50600	 => std_logic_vector(to_unsigned(127,8) ,
50601	 => std_logic_vector(to_unsigned(108,8) ,
50602	 => std_logic_vector(to_unsigned(112,8) ,
50603	 => std_logic_vector(to_unsigned(96,8) ,
50604	 => std_logic_vector(to_unsigned(92,8) ,
50605	 => std_logic_vector(to_unsigned(96,8) ,
50606	 => std_logic_vector(to_unsigned(108,8) ,
50607	 => std_logic_vector(to_unsigned(122,8) ,
50608	 => std_logic_vector(to_unsigned(114,8) ,
50609	 => std_logic_vector(to_unsigned(112,8) ,
50610	 => std_logic_vector(to_unsigned(124,8) ,
50611	 => std_logic_vector(to_unsigned(121,8) ,
50612	 => std_logic_vector(to_unsigned(125,8) ,
50613	 => std_logic_vector(to_unsigned(133,8) ,
50614	 => std_logic_vector(to_unsigned(141,8) ,
50615	 => std_logic_vector(to_unsigned(116,8) ,
50616	 => std_logic_vector(to_unsigned(97,8) ,
50617	 => std_logic_vector(to_unsigned(90,8) ,
50618	 => std_logic_vector(to_unsigned(88,8) ,
50619	 => std_logic_vector(to_unsigned(97,8) ,
50620	 => std_logic_vector(to_unsigned(97,8) ,
50621	 => std_logic_vector(to_unsigned(49,8) ,
50622	 => std_logic_vector(to_unsigned(48,8) ,
50623	 => std_logic_vector(to_unsigned(55,8) ,
50624	 => std_logic_vector(to_unsigned(71,8) ,
50625	 => std_logic_vector(to_unsigned(65,8) ,
50626	 => std_logic_vector(to_unsigned(57,8) ,
50627	 => std_logic_vector(to_unsigned(67,8) ,
50628	 => std_logic_vector(to_unsigned(124,8) ,
50629	 => std_logic_vector(to_unsigned(118,8) ,
50630	 => std_logic_vector(to_unsigned(87,8) ,
50631	 => std_logic_vector(to_unsigned(67,8) ,
50632	 => std_logic_vector(to_unsigned(88,8) ,
50633	 => std_logic_vector(to_unsigned(104,8) ,
50634	 => std_logic_vector(to_unsigned(78,8) ,
50635	 => std_logic_vector(to_unsigned(90,8) ,
50636	 => std_logic_vector(to_unsigned(92,8) ,
50637	 => std_logic_vector(to_unsigned(112,8) ,
50638	 => std_logic_vector(to_unsigned(97,8) ,
50639	 => std_logic_vector(to_unsigned(59,8) ,
50640	 => std_logic_vector(to_unsigned(49,8) ,
50641	 => std_logic_vector(to_unsigned(55,8) ,
50642	 => std_logic_vector(to_unsigned(61,8) ,
50643	 => std_logic_vector(to_unsigned(55,8) ,
50644	 => std_logic_vector(to_unsigned(52,8) ,
50645	 => std_logic_vector(to_unsigned(54,8) ,
50646	 => std_logic_vector(to_unsigned(49,8) ,
50647	 => std_logic_vector(to_unsigned(29,8) ,
50648	 => std_logic_vector(to_unsigned(24,8) ,
50649	 => std_logic_vector(to_unsigned(36,8) ,
50650	 => std_logic_vector(to_unsigned(45,8) ,
50651	 => std_logic_vector(to_unsigned(52,8) ,
50652	 => std_logic_vector(to_unsigned(52,8) ,
50653	 => std_logic_vector(to_unsigned(52,8) ,
50654	 => std_logic_vector(to_unsigned(54,8) ,
50655	 => std_logic_vector(to_unsigned(52,8) ,
50656	 => std_logic_vector(to_unsigned(47,8) ,
50657	 => std_logic_vector(to_unsigned(35,8) ,
50658	 => std_logic_vector(to_unsigned(32,8) ,
50659	 => std_logic_vector(to_unsigned(44,8) ,
50660	 => std_logic_vector(to_unsigned(49,8) ,
50661	 => std_logic_vector(to_unsigned(45,8) ,
50662	 => std_logic_vector(to_unsigned(44,8) ,
50663	 => std_logic_vector(to_unsigned(56,8) ,
50664	 => std_logic_vector(to_unsigned(81,8) ,
50665	 => std_logic_vector(to_unsigned(68,8) ,
50666	 => std_logic_vector(to_unsigned(56,8) ,
50667	 => std_logic_vector(to_unsigned(61,8) ,
50668	 => std_logic_vector(to_unsigned(59,8) ,
50669	 => std_logic_vector(to_unsigned(56,8) ,
50670	 => std_logic_vector(to_unsigned(57,8) ,
50671	 => std_logic_vector(to_unsigned(63,8) ,
50672	 => std_logic_vector(to_unsigned(58,8) ,
50673	 => std_logic_vector(to_unsigned(49,8) ,
50674	 => std_logic_vector(to_unsigned(41,8) ,
50675	 => std_logic_vector(to_unsigned(49,8) ,
50676	 => std_logic_vector(to_unsigned(47,8) ,
50677	 => std_logic_vector(to_unsigned(57,8) ,
50678	 => std_logic_vector(to_unsigned(34,8) ,
50679	 => std_logic_vector(to_unsigned(20,8) ,
50680	 => std_logic_vector(to_unsigned(30,8) ,
50681	 => std_logic_vector(to_unsigned(30,8) ,
50682	 => std_logic_vector(to_unsigned(29,8) ,
50683	 => std_logic_vector(to_unsigned(33,8) ,
50684	 => std_logic_vector(to_unsigned(74,8) ,
50685	 => std_logic_vector(to_unsigned(69,8) ,
50686	 => std_logic_vector(to_unsigned(59,8) ,
50687	 => std_logic_vector(to_unsigned(60,8) ,
50688	 => std_logic_vector(to_unsigned(47,8) ,
50689	 => std_logic_vector(to_unsigned(48,8) ,
50690	 => std_logic_vector(to_unsigned(37,8) ,
50691	 => std_logic_vector(to_unsigned(34,8) ,
50692	 => std_logic_vector(to_unsigned(51,8) ,
50693	 => std_logic_vector(to_unsigned(35,8) ,
50694	 => std_logic_vector(to_unsigned(36,8) ,
50695	 => std_logic_vector(to_unsigned(36,8) ,
50696	 => std_logic_vector(to_unsigned(14,8) ,
50697	 => std_logic_vector(to_unsigned(11,8) ,
50698	 => std_logic_vector(to_unsigned(12,8) ,
50699	 => std_logic_vector(to_unsigned(12,8) ,
50700	 => std_logic_vector(to_unsigned(26,8) ,
50701	 => std_logic_vector(to_unsigned(46,8) ,
50702	 => std_logic_vector(to_unsigned(63,8) ,
50703	 => std_logic_vector(to_unsigned(54,8) ,
50704	 => std_logic_vector(to_unsigned(72,8) ,
50705	 => std_logic_vector(to_unsigned(96,8) ,
50706	 => std_logic_vector(to_unsigned(62,8) ,
50707	 => std_logic_vector(to_unsigned(27,8) ,
50708	 => std_logic_vector(to_unsigned(6,8) ,
50709	 => std_logic_vector(to_unsigned(31,8) ,
50710	 => std_logic_vector(to_unsigned(80,8) ,
50711	 => std_logic_vector(to_unsigned(41,8) ,
50712	 => std_logic_vector(to_unsigned(72,8) ,
50713	 => std_logic_vector(to_unsigned(52,8) ,
50714	 => std_logic_vector(to_unsigned(56,8) ,
50715	 => std_logic_vector(to_unsigned(35,8) ,
50716	 => std_logic_vector(to_unsigned(81,8) ,
50717	 => std_logic_vector(to_unsigned(67,8) ,
50718	 => std_logic_vector(to_unsigned(23,8) ,
50719	 => std_logic_vector(to_unsigned(9,8) ,
50720	 => std_logic_vector(to_unsigned(12,8) ,
50721	 => std_logic_vector(to_unsigned(63,8) ,
50722	 => std_logic_vector(to_unsigned(60,8) ,
50723	 => std_logic_vector(to_unsigned(61,8) ,
50724	 => std_logic_vector(to_unsigned(59,8) ,
50725	 => std_logic_vector(to_unsigned(62,8) ,
50726	 => std_logic_vector(to_unsigned(19,8) ,
50727	 => std_logic_vector(to_unsigned(13,8) ,
50728	 => std_logic_vector(to_unsigned(79,8) ,
50729	 => std_logic_vector(to_unsigned(43,8) ,
50730	 => std_logic_vector(to_unsigned(19,8) ,
50731	 => std_logic_vector(to_unsigned(6,8) ,
50732	 => std_logic_vector(to_unsigned(14,8) ,
50733	 => std_logic_vector(to_unsigned(66,8) ,
50734	 => std_logic_vector(to_unsigned(31,8) ,
50735	 => std_logic_vector(to_unsigned(29,8) ,
50736	 => std_logic_vector(to_unsigned(47,8) ,
50737	 => std_logic_vector(to_unsigned(31,8) ,
50738	 => std_logic_vector(to_unsigned(34,8) ,
50739	 => std_logic_vector(to_unsigned(60,8) ,
50740	 => std_logic_vector(to_unsigned(66,8) ,
50741	 => std_logic_vector(to_unsigned(63,8) ,
50742	 => std_logic_vector(to_unsigned(43,8) ,
50743	 => std_logic_vector(to_unsigned(17,8) ,
50744	 => std_logic_vector(to_unsigned(24,8) ,
50745	 => std_logic_vector(to_unsigned(61,8) ,
50746	 => std_logic_vector(to_unsigned(44,8) ,
50747	 => std_logic_vector(to_unsigned(30,8) ,
50748	 => std_logic_vector(to_unsigned(25,8) ,
50749	 => std_logic_vector(to_unsigned(27,8) ,
50750	 => std_logic_vector(to_unsigned(35,8) ,
50751	 => std_logic_vector(to_unsigned(26,8) ,
50752	 => std_logic_vector(to_unsigned(24,8) ,
50753	 => std_logic_vector(to_unsigned(18,8) ,
50754	 => std_logic_vector(to_unsigned(16,8) ,
50755	 => std_logic_vector(to_unsigned(32,8) ,
50756	 => std_logic_vector(to_unsigned(45,8) ,
50757	 => std_logic_vector(to_unsigned(32,8) ,
50758	 => std_logic_vector(to_unsigned(23,8) ,
50759	 => std_logic_vector(to_unsigned(26,8) ,
50760	 => std_logic_vector(to_unsigned(19,8) ,
50761	 => std_logic_vector(to_unsigned(30,8) ,
50762	 => std_logic_vector(to_unsigned(33,8) ,
50763	 => std_logic_vector(to_unsigned(28,8) ,
50764	 => std_logic_vector(to_unsigned(29,8) ,
50765	 => std_logic_vector(to_unsigned(52,8) ,
50766	 => std_logic_vector(to_unsigned(78,8) ,
50767	 => std_logic_vector(to_unsigned(56,8) ,
50768	 => std_logic_vector(to_unsigned(65,8) ,
50769	 => std_logic_vector(to_unsigned(60,8) ,
50770	 => std_logic_vector(to_unsigned(27,8) ,
50771	 => std_logic_vector(to_unsigned(30,8) ,
50772	 => std_logic_vector(to_unsigned(27,8) ,
50773	 => std_logic_vector(to_unsigned(27,8) ,
50774	 => std_logic_vector(to_unsigned(73,8) ,
50775	 => std_logic_vector(to_unsigned(85,8) ,
50776	 => std_logic_vector(to_unsigned(37,8) ,
50777	 => std_logic_vector(to_unsigned(26,8) ,
50778	 => std_logic_vector(to_unsigned(35,8) ,
50779	 => std_logic_vector(to_unsigned(14,8) ,
50780	 => std_logic_vector(to_unsigned(22,8) ,
50781	 => std_logic_vector(to_unsigned(30,8) ,
50782	 => std_logic_vector(to_unsigned(22,8) ,
50783	 => std_logic_vector(to_unsigned(41,8) ,
50784	 => std_logic_vector(to_unsigned(30,8) ,
50785	 => std_logic_vector(to_unsigned(29,8) ,
50786	 => std_logic_vector(to_unsigned(27,8) ,
50787	 => std_logic_vector(to_unsigned(20,8) ,
50788	 => std_logic_vector(to_unsigned(20,8) ,
50789	 => std_logic_vector(to_unsigned(19,8) ,
50790	 => std_logic_vector(to_unsigned(22,8) ,
50791	 => std_logic_vector(to_unsigned(22,8) ,
50792	 => std_logic_vector(to_unsigned(23,8) ,
50793	 => std_logic_vector(to_unsigned(28,8) ,
50794	 => std_logic_vector(to_unsigned(22,8) ,
50795	 => std_logic_vector(to_unsigned(16,8) ,
50796	 => std_logic_vector(to_unsigned(20,8) ,
50797	 => std_logic_vector(to_unsigned(18,8) ,
50798	 => std_logic_vector(to_unsigned(27,8) ,
50799	 => std_logic_vector(to_unsigned(53,8) ,
50800	 => std_logic_vector(to_unsigned(35,8) ,
50801	 => std_logic_vector(to_unsigned(15,8) ,
50802	 => std_logic_vector(to_unsigned(16,8) ,
50803	 => std_logic_vector(to_unsigned(16,8) ,
50804	 => std_logic_vector(to_unsigned(17,8) ,
50805	 => std_logic_vector(to_unsigned(19,8) ,
50806	 => std_logic_vector(to_unsigned(24,8) ,
50807	 => std_logic_vector(to_unsigned(31,8) ,
50808	 => std_logic_vector(to_unsigned(42,8) ,
50809	 => std_logic_vector(to_unsigned(30,8) ,
50810	 => std_logic_vector(to_unsigned(72,8) ,
50811	 => std_logic_vector(to_unsigned(74,8) ,
50812	 => std_logic_vector(to_unsigned(82,8) ,
50813	 => std_logic_vector(to_unsigned(43,8) ,
50814	 => std_logic_vector(to_unsigned(1,8) ,
50815	 => std_logic_vector(to_unsigned(1,8) ,
50816	 => std_logic_vector(to_unsigned(13,8) ,
50817	 => std_logic_vector(to_unsigned(66,8) ,
50818	 => std_logic_vector(to_unsigned(91,8) ,
50819	 => std_logic_vector(to_unsigned(52,8) ,
50820	 => std_logic_vector(to_unsigned(87,8) ,
50821	 => std_logic_vector(to_unsigned(76,8) ,
50822	 => std_logic_vector(to_unsigned(81,8) ,
50823	 => std_logic_vector(to_unsigned(65,8) ,
50824	 => std_logic_vector(to_unsigned(97,8) ,
50825	 => std_logic_vector(to_unsigned(100,8) ,
50826	 => std_logic_vector(to_unsigned(68,8) ,
50827	 => std_logic_vector(to_unsigned(35,8) ,
50828	 => std_logic_vector(to_unsigned(53,8) ,
50829	 => std_logic_vector(to_unsigned(45,8) ,
50830	 => std_logic_vector(to_unsigned(35,8) ,
50831	 => std_logic_vector(to_unsigned(32,8) ,
50832	 => std_logic_vector(to_unsigned(35,8) ,
50833	 => std_logic_vector(to_unsigned(23,8) ,
50834	 => std_logic_vector(to_unsigned(22,8) ,
50835	 => std_logic_vector(to_unsigned(33,8) ,
50836	 => std_logic_vector(to_unsigned(22,8) ,
50837	 => std_logic_vector(to_unsigned(3,8) ,
50838	 => std_logic_vector(to_unsigned(0,8) ,
50839	 => std_logic_vector(to_unsigned(0,8) ,
50840	 => std_logic_vector(to_unsigned(0,8) ,
50841	 => std_logic_vector(to_unsigned(1,8) ,
50842	 => std_logic_vector(to_unsigned(25,8) ,
50843	 => std_logic_vector(to_unsigned(33,8) ,
50844	 => std_logic_vector(to_unsigned(29,8) ,
50845	 => std_logic_vector(to_unsigned(32,8) ,
50846	 => std_logic_vector(to_unsigned(29,8) ,
50847	 => std_logic_vector(to_unsigned(22,8) ,
50848	 => std_logic_vector(to_unsigned(26,8) ,
50849	 => std_logic_vector(to_unsigned(19,8) ,
50850	 => std_logic_vector(to_unsigned(22,8) ,
50851	 => std_logic_vector(to_unsigned(29,8) ,
50852	 => std_logic_vector(to_unsigned(32,8) ,
50853	 => std_logic_vector(to_unsigned(41,8) ,
50854	 => std_logic_vector(to_unsigned(38,8) ,
50855	 => std_logic_vector(to_unsigned(61,8) ,
50856	 => std_logic_vector(to_unsigned(38,8) ,
50857	 => std_logic_vector(to_unsigned(16,8) ,
50858	 => std_logic_vector(to_unsigned(17,8) ,
50859	 => std_logic_vector(to_unsigned(11,8) ,
50860	 => std_logic_vector(to_unsigned(23,8) ,
50861	 => std_logic_vector(to_unsigned(56,8) ,
50862	 => std_logic_vector(to_unsigned(52,8) ,
50863	 => std_logic_vector(to_unsigned(25,8) ,
50864	 => std_logic_vector(to_unsigned(9,8) ,
50865	 => std_logic_vector(to_unsigned(15,8) ,
50866	 => std_logic_vector(to_unsigned(13,8) ,
50867	 => std_logic_vector(to_unsigned(17,8) ,
50868	 => std_logic_vector(to_unsigned(42,8) ,
50869	 => std_logic_vector(to_unsigned(35,8) ,
50870	 => std_logic_vector(to_unsigned(44,8) ,
50871	 => std_logic_vector(to_unsigned(25,8) ,
50872	 => std_logic_vector(to_unsigned(25,8) ,
50873	 => std_logic_vector(to_unsigned(27,8) ,
50874	 => std_logic_vector(to_unsigned(26,8) ,
50875	 => std_logic_vector(to_unsigned(21,8) ,
50876	 => std_logic_vector(to_unsigned(34,8) ,
50877	 => std_logic_vector(to_unsigned(30,8) ,
50878	 => std_logic_vector(to_unsigned(34,8) ,
50879	 => std_logic_vector(to_unsigned(44,8) ,
50880	 => std_logic_vector(to_unsigned(13,8) ,
50881	 => std_logic_vector(to_unsigned(111,8) ,
50882	 => std_logic_vector(to_unsigned(104,8) ,
50883	 => std_logic_vector(to_unsigned(104,8) ,
50884	 => std_logic_vector(to_unsigned(111,8) ,
50885	 => std_logic_vector(to_unsigned(112,8) ,
50886	 => std_logic_vector(to_unsigned(118,8) ,
50887	 => std_logic_vector(to_unsigned(125,8) ,
50888	 => std_logic_vector(to_unsigned(101,8) ,
50889	 => std_logic_vector(to_unsigned(112,8) ,
50890	 => std_logic_vector(to_unsigned(103,8) ,
50891	 => std_logic_vector(to_unsigned(96,8) ,
50892	 => std_logic_vector(to_unsigned(100,8) ,
50893	 => std_logic_vector(to_unsigned(101,8) ,
50894	 => std_logic_vector(to_unsigned(108,8) ,
50895	 => std_logic_vector(to_unsigned(100,8) ,
50896	 => std_logic_vector(to_unsigned(103,8) ,
50897	 => std_logic_vector(to_unsigned(114,8) ,
50898	 => std_logic_vector(to_unsigned(96,8) ,
50899	 => std_logic_vector(to_unsigned(121,8) ,
50900	 => std_logic_vector(to_unsigned(116,8) ,
50901	 => std_logic_vector(to_unsigned(128,8) ,
50902	 => std_logic_vector(to_unsigned(130,8) ,
50903	 => std_logic_vector(to_unsigned(103,8) ,
50904	 => std_logic_vector(to_unsigned(88,8) ,
50905	 => std_logic_vector(to_unsigned(74,8) ,
50906	 => std_logic_vector(to_unsigned(74,8) ,
50907	 => std_logic_vector(to_unsigned(66,8) ,
50908	 => std_logic_vector(to_unsigned(78,8) ,
50909	 => std_logic_vector(to_unsigned(88,8) ,
50910	 => std_logic_vector(to_unsigned(87,8) ,
50911	 => std_logic_vector(to_unsigned(76,8) ,
50912	 => std_logic_vector(to_unsigned(79,8) ,
50913	 => std_logic_vector(to_unsigned(88,8) ,
50914	 => std_logic_vector(to_unsigned(65,8) ,
50915	 => std_logic_vector(to_unsigned(35,8) ,
50916	 => std_logic_vector(to_unsigned(41,8) ,
50917	 => std_logic_vector(to_unsigned(45,8) ,
50918	 => std_logic_vector(to_unsigned(45,8) ,
50919	 => std_logic_vector(to_unsigned(79,8) ,
50920	 => std_logic_vector(to_unsigned(114,8) ,
50921	 => std_logic_vector(to_unsigned(114,8) ,
50922	 => std_logic_vector(to_unsigned(121,8) ,
50923	 => std_logic_vector(to_unsigned(119,8) ,
50924	 => std_logic_vector(to_unsigned(125,8) ,
50925	 => std_logic_vector(to_unsigned(130,8) ,
50926	 => std_logic_vector(to_unsigned(122,8) ,
50927	 => std_logic_vector(to_unsigned(125,8) ,
50928	 => std_logic_vector(to_unsigned(116,8) ,
50929	 => std_logic_vector(to_unsigned(64,8) ,
50930	 => std_logic_vector(to_unsigned(82,8) ,
50931	 => std_logic_vector(to_unsigned(73,8) ,
50932	 => std_logic_vector(to_unsigned(95,8) ,
50933	 => std_logic_vector(to_unsigned(93,8) ,
50934	 => std_logic_vector(to_unsigned(99,8) ,
50935	 => std_logic_vector(to_unsigned(109,8) ,
50936	 => std_logic_vector(to_unsigned(125,8) ,
50937	 => std_logic_vector(to_unsigned(141,8) ,
50938	 => std_logic_vector(to_unsigned(136,8) ,
50939	 => std_logic_vector(to_unsigned(139,8) ,
50940	 => std_logic_vector(to_unsigned(147,8) ,
50941	 => std_logic_vector(to_unsigned(93,8) ,
50942	 => std_logic_vector(to_unsigned(86,8) ,
50943	 => std_logic_vector(to_unsigned(101,8) ,
50944	 => std_logic_vector(to_unsigned(92,8) ,
50945	 => std_logic_vector(to_unsigned(85,8) ,
50946	 => std_logic_vector(to_unsigned(90,8) ,
50947	 => std_logic_vector(to_unsigned(78,8) ,
50948	 => std_logic_vector(to_unsigned(88,8) ,
50949	 => std_logic_vector(to_unsigned(84,8) ,
50950	 => std_logic_vector(to_unsigned(93,8) ,
50951	 => std_logic_vector(to_unsigned(127,8) ,
50952	 => std_logic_vector(to_unsigned(99,8) ,
50953	 => std_logic_vector(to_unsigned(81,8) ,
50954	 => std_logic_vector(to_unsigned(68,8) ,
50955	 => std_logic_vector(to_unsigned(73,8) ,
50956	 => std_logic_vector(to_unsigned(88,8) ,
50957	 => std_logic_vector(to_unsigned(108,8) ,
50958	 => std_logic_vector(to_unsigned(93,8) ,
50959	 => std_logic_vector(to_unsigned(58,8) ,
50960	 => std_logic_vector(to_unsigned(53,8) ,
50961	 => std_logic_vector(to_unsigned(61,8) ,
50962	 => std_logic_vector(to_unsigned(61,8) ,
50963	 => std_logic_vector(to_unsigned(59,8) ,
50964	 => std_logic_vector(to_unsigned(56,8) ,
50965	 => std_logic_vector(to_unsigned(65,8) ,
50966	 => std_logic_vector(to_unsigned(55,8) ,
50967	 => std_logic_vector(to_unsigned(39,8) ,
50968	 => std_logic_vector(to_unsigned(36,8) ,
50969	 => std_logic_vector(to_unsigned(43,8) ,
50970	 => std_logic_vector(to_unsigned(53,8) ,
50971	 => std_logic_vector(to_unsigned(50,8) ,
50972	 => std_logic_vector(to_unsigned(58,8) ,
50973	 => std_logic_vector(to_unsigned(67,8) ,
50974	 => std_logic_vector(to_unsigned(57,8) ,
50975	 => std_logic_vector(to_unsigned(51,8) ,
50976	 => std_logic_vector(to_unsigned(44,8) ,
50977	 => std_logic_vector(to_unsigned(29,8) ,
50978	 => std_logic_vector(to_unsigned(25,8) ,
50979	 => std_logic_vector(to_unsigned(35,8) ,
50980	 => std_logic_vector(to_unsigned(35,8) ,
50981	 => std_logic_vector(to_unsigned(32,8) ,
50982	 => std_logic_vector(to_unsigned(35,8) ,
50983	 => std_logic_vector(to_unsigned(45,8) ,
50984	 => std_logic_vector(to_unsigned(71,8) ,
50985	 => std_logic_vector(to_unsigned(66,8) ,
50986	 => std_logic_vector(to_unsigned(52,8) ,
50987	 => std_logic_vector(to_unsigned(48,8) ,
50988	 => std_logic_vector(to_unsigned(56,8) ,
50989	 => std_logic_vector(to_unsigned(58,8) ,
50990	 => std_logic_vector(to_unsigned(40,8) ,
50991	 => std_logic_vector(to_unsigned(47,8) ,
50992	 => std_logic_vector(to_unsigned(55,8) ,
50993	 => std_logic_vector(to_unsigned(53,8) ,
50994	 => std_logic_vector(to_unsigned(50,8) ,
50995	 => std_logic_vector(to_unsigned(51,8) ,
50996	 => std_logic_vector(to_unsigned(56,8) ,
50997	 => std_logic_vector(to_unsigned(52,8) ,
50998	 => std_logic_vector(to_unsigned(41,8) ,
50999	 => std_logic_vector(to_unsigned(24,8) ,
51000	 => std_logic_vector(to_unsigned(22,8) ,
51001	 => std_logic_vector(to_unsigned(30,8) ,
51002	 => std_logic_vector(to_unsigned(37,8) ,
51003	 => std_logic_vector(to_unsigned(30,8) ,
51004	 => std_logic_vector(to_unsigned(74,8) ,
51005	 => std_logic_vector(to_unsigned(82,8) ,
51006	 => std_logic_vector(to_unsigned(60,8) ,
51007	 => std_logic_vector(to_unsigned(49,8) ,
51008	 => std_logic_vector(to_unsigned(46,8) ,
51009	 => std_logic_vector(to_unsigned(51,8) ,
51010	 => std_logic_vector(to_unsigned(35,8) ,
51011	 => std_logic_vector(to_unsigned(35,8) ,
51012	 => std_logic_vector(to_unsigned(45,8) ,
51013	 => std_logic_vector(to_unsigned(37,8) ,
51014	 => std_logic_vector(to_unsigned(40,8) ,
51015	 => std_logic_vector(to_unsigned(35,8) ,
51016	 => std_logic_vector(to_unsigned(14,8) ,
51017	 => std_logic_vector(to_unsigned(9,8) ,
51018	 => std_logic_vector(to_unsigned(22,8) ,
51019	 => std_logic_vector(to_unsigned(51,8) ,
51020	 => std_logic_vector(to_unsigned(28,8) ,
51021	 => std_logic_vector(to_unsigned(23,8) ,
51022	 => std_logic_vector(to_unsigned(29,8) ,
51023	 => std_logic_vector(to_unsigned(24,8) ,
51024	 => std_logic_vector(to_unsigned(25,8) ,
51025	 => std_logic_vector(to_unsigned(31,8) ,
51026	 => std_logic_vector(to_unsigned(43,8) ,
51027	 => std_logic_vector(to_unsigned(46,8) ,
51028	 => std_logic_vector(to_unsigned(30,8) ,
51029	 => std_logic_vector(to_unsigned(42,8) ,
51030	 => std_logic_vector(to_unsigned(62,8) ,
51031	 => std_logic_vector(to_unsigned(60,8) ,
51032	 => std_logic_vector(to_unsigned(81,8) ,
51033	 => std_logic_vector(to_unsigned(69,8) ,
51034	 => std_logic_vector(to_unsigned(64,8) ,
51035	 => std_logic_vector(to_unsigned(20,8) ,
51036	 => std_logic_vector(to_unsigned(79,8) ,
51037	 => std_logic_vector(to_unsigned(72,8) ,
51038	 => std_logic_vector(to_unsigned(18,8) ,
51039	 => std_logic_vector(to_unsigned(8,8) ,
51040	 => std_logic_vector(to_unsigned(8,8) ,
51041	 => std_logic_vector(to_unsigned(56,8) ,
51042	 => std_logic_vector(to_unsigned(31,8) ,
51043	 => std_logic_vector(to_unsigned(35,8) ,
51044	 => std_logic_vector(to_unsigned(48,8) ,
51045	 => std_logic_vector(to_unsigned(41,8) ,
51046	 => std_logic_vector(to_unsigned(29,8) ,
51047	 => std_logic_vector(to_unsigned(24,8) ,
51048	 => std_logic_vector(to_unsigned(77,8) ,
51049	 => std_logic_vector(to_unsigned(41,8) ,
51050	 => std_logic_vector(to_unsigned(17,8) ,
51051	 => std_logic_vector(to_unsigned(6,8) ,
51052	 => std_logic_vector(to_unsigned(15,8) ,
51053	 => std_logic_vector(to_unsigned(79,8) ,
51054	 => std_logic_vector(to_unsigned(45,8) ,
51055	 => std_logic_vector(to_unsigned(41,8) ,
51056	 => std_logic_vector(to_unsigned(64,8) ,
51057	 => std_logic_vector(to_unsigned(41,8) ,
51058	 => std_logic_vector(to_unsigned(30,8) ,
51059	 => std_logic_vector(to_unsigned(54,8) ,
51060	 => std_logic_vector(to_unsigned(35,8) ,
51061	 => std_logic_vector(to_unsigned(54,8) ,
51062	 => std_logic_vector(to_unsigned(35,8) ,
51063	 => std_logic_vector(to_unsigned(35,8) ,
51064	 => std_logic_vector(to_unsigned(53,8) ,
51065	 => std_logic_vector(to_unsigned(44,8) ,
51066	 => std_logic_vector(to_unsigned(19,8) ,
51067	 => std_logic_vector(to_unsigned(10,8) ,
51068	 => std_logic_vector(to_unsigned(24,8) ,
51069	 => std_logic_vector(to_unsigned(29,8) ,
51070	 => std_logic_vector(to_unsigned(27,8) ,
51071	 => std_logic_vector(to_unsigned(24,8) ,
51072	 => std_logic_vector(to_unsigned(31,8) ,
51073	 => std_logic_vector(to_unsigned(37,8) ,
51074	 => std_logic_vector(to_unsigned(37,8) ,
51075	 => std_logic_vector(to_unsigned(43,8) ,
51076	 => std_logic_vector(to_unsigned(37,8) ,
51077	 => std_logic_vector(to_unsigned(12,8) ,
51078	 => std_logic_vector(to_unsigned(23,8) ,
51079	 => std_logic_vector(to_unsigned(17,8) ,
51080	 => std_logic_vector(to_unsigned(6,8) ,
51081	 => std_logic_vector(to_unsigned(12,8) ,
51082	 => std_logic_vector(to_unsigned(31,8) ,
51083	 => std_logic_vector(to_unsigned(30,8) ,
51084	 => std_logic_vector(to_unsigned(23,8) ,
51085	 => std_logic_vector(to_unsigned(35,8) ,
51086	 => std_logic_vector(to_unsigned(39,8) ,
51087	 => std_logic_vector(to_unsigned(45,8) ,
51088	 => std_logic_vector(to_unsigned(59,8) ,
51089	 => std_logic_vector(to_unsigned(63,8) ,
51090	 => std_logic_vector(to_unsigned(28,8) ,
51091	 => std_logic_vector(to_unsigned(23,8) ,
51092	 => std_logic_vector(to_unsigned(24,8) ,
51093	 => std_logic_vector(to_unsigned(21,8) ,
51094	 => std_logic_vector(to_unsigned(27,8) ,
51095	 => std_logic_vector(to_unsigned(29,8) ,
51096	 => std_logic_vector(to_unsigned(22,8) ,
51097	 => std_logic_vector(to_unsigned(22,8) ,
51098	 => std_logic_vector(to_unsigned(26,8) ,
51099	 => std_logic_vector(to_unsigned(12,8) ,
51100	 => std_logic_vector(to_unsigned(17,8) ,
51101	 => std_logic_vector(to_unsigned(17,8) ,
51102	 => std_logic_vector(to_unsigned(23,8) ,
51103	 => std_logic_vector(to_unsigned(27,8) ,
51104	 => std_logic_vector(to_unsigned(15,8) ,
51105	 => std_logic_vector(to_unsigned(15,8) ,
51106	 => std_logic_vector(to_unsigned(15,8) ,
51107	 => std_logic_vector(to_unsigned(17,8) ,
51108	 => std_logic_vector(to_unsigned(19,8) ,
51109	 => std_logic_vector(to_unsigned(16,8) ,
51110	 => std_logic_vector(to_unsigned(21,8) ,
51111	 => std_logic_vector(to_unsigned(24,8) ,
51112	 => std_logic_vector(to_unsigned(24,8) ,
51113	 => std_logic_vector(to_unsigned(23,8) ,
51114	 => std_logic_vector(to_unsigned(14,8) ,
51115	 => std_logic_vector(to_unsigned(11,8) ,
51116	 => std_logic_vector(to_unsigned(14,8) ,
51117	 => std_logic_vector(to_unsigned(24,8) ,
51118	 => std_logic_vector(to_unsigned(29,8) ,
51119	 => std_logic_vector(to_unsigned(28,8) ,
51120	 => std_logic_vector(to_unsigned(24,8) ,
51121	 => std_logic_vector(to_unsigned(22,8) ,
51122	 => std_logic_vector(to_unsigned(32,8) ,
51123	 => std_logic_vector(to_unsigned(21,8) ,
51124	 => std_logic_vector(to_unsigned(15,8) ,
51125	 => std_logic_vector(to_unsigned(12,8) ,
51126	 => std_logic_vector(to_unsigned(18,8) ,
51127	 => std_logic_vector(to_unsigned(33,8) ,
51128	 => std_logic_vector(to_unsigned(43,8) ,
51129	 => std_logic_vector(to_unsigned(28,8) ,
51130	 => std_logic_vector(to_unsigned(62,8) ,
51131	 => std_logic_vector(to_unsigned(93,8) ,
51132	 => std_logic_vector(to_unsigned(90,8) ,
51133	 => std_logic_vector(to_unsigned(67,8) ,
51134	 => std_logic_vector(to_unsigned(13,8) ,
51135	 => std_logic_vector(to_unsigned(1,8) ,
51136	 => std_logic_vector(to_unsigned(2,8) ,
51137	 => std_logic_vector(to_unsigned(37,8) ,
51138	 => std_logic_vector(to_unsigned(91,8) ,
51139	 => std_logic_vector(to_unsigned(51,8) ,
51140	 => std_logic_vector(to_unsigned(85,8) ,
51141	 => std_logic_vector(to_unsigned(68,8) ,
51142	 => std_logic_vector(to_unsigned(78,8) ,
51143	 => std_logic_vector(to_unsigned(65,8) ,
51144	 => std_logic_vector(to_unsigned(85,8) ,
51145	 => std_logic_vector(to_unsigned(78,8) ,
51146	 => std_logic_vector(to_unsigned(55,8) ,
51147	 => std_logic_vector(to_unsigned(22,8) ,
51148	 => std_logic_vector(to_unsigned(30,8) ,
51149	 => std_logic_vector(to_unsigned(32,8) ,
51150	 => std_logic_vector(to_unsigned(19,8) ,
51151	 => std_logic_vector(to_unsigned(17,8) ,
51152	 => std_logic_vector(to_unsigned(13,8) ,
51153	 => std_logic_vector(to_unsigned(9,8) ,
51154	 => std_logic_vector(to_unsigned(9,8) ,
51155	 => std_logic_vector(to_unsigned(13,8) ,
51156	 => std_logic_vector(to_unsigned(20,8) ,
51157	 => std_logic_vector(to_unsigned(6,8) ,
51158	 => std_logic_vector(to_unsigned(0,8) ,
51159	 => std_logic_vector(to_unsigned(0,8) ,
51160	 => std_logic_vector(to_unsigned(0,8) ,
51161	 => std_logic_vector(to_unsigned(0,8) ,
51162	 => std_logic_vector(to_unsigned(14,8) ,
51163	 => std_logic_vector(to_unsigned(29,8) ,
51164	 => std_logic_vector(to_unsigned(9,8) ,
51165	 => std_logic_vector(to_unsigned(17,8) ,
51166	 => std_logic_vector(to_unsigned(26,8) ,
51167	 => std_logic_vector(to_unsigned(15,8) ,
51168	 => std_logic_vector(to_unsigned(14,8) ,
51169	 => std_logic_vector(to_unsigned(13,8) ,
51170	 => std_logic_vector(to_unsigned(23,8) ,
51171	 => std_logic_vector(to_unsigned(29,8) ,
51172	 => std_logic_vector(to_unsigned(34,8) ,
51173	 => std_logic_vector(to_unsigned(42,8) ,
51174	 => std_logic_vector(to_unsigned(35,8) ,
51175	 => std_logic_vector(to_unsigned(37,8) ,
51176	 => std_logic_vector(to_unsigned(29,8) ,
51177	 => std_logic_vector(to_unsigned(23,8) ,
51178	 => std_logic_vector(to_unsigned(17,8) ,
51179	 => std_logic_vector(to_unsigned(38,8) ,
51180	 => std_logic_vector(to_unsigned(53,8) ,
51181	 => std_logic_vector(to_unsigned(41,8) ,
51182	 => std_logic_vector(to_unsigned(42,8) ,
51183	 => std_logic_vector(to_unsigned(23,8) ,
51184	 => std_logic_vector(to_unsigned(11,8) ,
51185	 => std_logic_vector(to_unsigned(10,8) ,
51186	 => std_logic_vector(to_unsigned(7,8) ,
51187	 => std_logic_vector(to_unsigned(13,8) ,
51188	 => std_logic_vector(to_unsigned(48,8) ,
51189	 => std_logic_vector(to_unsigned(41,8) ,
51190	 => std_logic_vector(to_unsigned(41,8) ,
51191	 => std_logic_vector(to_unsigned(32,8) ,
51192	 => std_logic_vector(to_unsigned(46,8) ,
51193	 => std_logic_vector(to_unsigned(47,8) ,
51194	 => std_logic_vector(to_unsigned(47,8) ,
51195	 => std_logic_vector(to_unsigned(51,8) ,
51196	 => std_logic_vector(to_unsigned(57,8) ,
51197	 => std_logic_vector(to_unsigned(51,8) ,
51198	 => std_logic_vector(to_unsigned(45,8) ,
51199	 => std_logic_vector(to_unsigned(45,8) ,
51200	 => std_logic_vector(to_unsigned(17,8) ,
51201	 => std_logic_vector(to_unsigned(119,8) ,
51202	 => std_logic_vector(to_unsigned(107,8) ,
51203	 => std_logic_vector(to_unsigned(104,8) ,
51204	 => std_logic_vector(to_unsigned(95,8) ,
51205	 => std_logic_vector(to_unsigned(71,8) ,
51206	 => std_logic_vector(to_unsigned(76,8) ,
51207	 => std_logic_vector(to_unsigned(88,8) ,
51208	 => std_logic_vector(to_unsigned(95,8) ,
51209	 => std_logic_vector(to_unsigned(116,8) ,
51210	 => std_logic_vector(to_unsigned(115,8) ,
51211	 => std_logic_vector(to_unsigned(127,8) ,
51212	 => std_logic_vector(to_unsigned(124,8) ,
51213	 => std_logic_vector(to_unsigned(122,8) ,
51214	 => std_logic_vector(to_unsigned(122,8) ,
51215	 => std_logic_vector(to_unsigned(99,8) ,
51216	 => std_logic_vector(to_unsigned(87,8) ,
51217	 => std_logic_vector(to_unsigned(99,8) ,
51218	 => std_logic_vector(to_unsigned(99,8) ,
51219	 => std_logic_vector(to_unsigned(119,8) ,
51220	 => std_logic_vector(to_unsigned(130,8) ,
51221	 => std_logic_vector(to_unsigned(118,8) ,
51222	 => std_logic_vector(to_unsigned(79,8) ,
51223	 => std_logic_vector(to_unsigned(68,8) ,
51224	 => std_logic_vector(to_unsigned(84,8) ,
51225	 => std_logic_vector(to_unsigned(90,8) ,
51226	 => std_logic_vector(to_unsigned(122,8) ,
51227	 => std_logic_vector(to_unsigned(108,8) ,
51228	 => std_logic_vector(to_unsigned(84,8) ,
51229	 => std_logic_vector(to_unsigned(78,8) ,
51230	 => std_logic_vector(to_unsigned(77,8) ,
51231	 => std_logic_vector(to_unsigned(76,8) ,
51232	 => std_logic_vector(to_unsigned(79,8) ,
51233	 => std_logic_vector(to_unsigned(85,8) ,
51234	 => std_logic_vector(to_unsigned(61,8) ,
51235	 => std_logic_vector(to_unsigned(35,8) ,
51236	 => std_logic_vector(to_unsigned(39,8) ,
51237	 => std_logic_vector(to_unsigned(41,8) ,
51238	 => std_logic_vector(to_unsigned(36,8) ,
51239	 => std_logic_vector(to_unsigned(62,8) ,
51240	 => std_logic_vector(to_unsigned(99,8) ,
51241	 => std_logic_vector(to_unsigned(87,8) ,
51242	 => std_logic_vector(to_unsigned(95,8) ,
51243	 => std_logic_vector(to_unsigned(105,8) ,
51244	 => std_logic_vector(to_unsigned(119,8) ,
51245	 => std_logic_vector(to_unsigned(124,8) ,
51246	 => std_logic_vector(to_unsigned(111,8) ,
51247	 => std_logic_vector(to_unsigned(115,8) ,
51248	 => std_logic_vector(to_unsigned(131,8) ,
51249	 => std_logic_vector(to_unsigned(62,8) ,
51250	 => std_logic_vector(to_unsigned(62,8) ,
51251	 => std_logic_vector(to_unsigned(68,8) ,
51252	 => std_logic_vector(to_unsigned(86,8) ,
51253	 => std_logic_vector(to_unsigned(73,8) ,
51254	 => std_logic_vector(to_unsigned(61,8) ,
51255	 => std_logic_vector(to_unsigned(66,8) ,
51256	 => std_logic_vector(to_unsigned(114,8) ,
51257	 => std_logic_vector(to_unsigned(144,8) ,
51258	 => std_logic_vector(to_unsigned(142,8) ,
51259	 => std_logic_vector(to_unsigned(133,8) ,
51260	 => std_logic_vector(to_unsigned(139,8) ,
51261	 => std_logic_vector(to_unsigned(131,8) ,
51262	 => std_logic_vector(to_unsigned(88,8) ,
51263	 => std_logic_vector(to_unsigned(104,8) ,
51264	 => std_logic_vector(to_unsigned(122,8) ,
51265	 => std_logic_vector(to_unsigned(124,8) ,
51266	 => std_logic_vector(to_unsigned(141,8) ,
51267	 => std_logic_vector(to_unsigned(147,8) ,
51268	 => std_logic_vector(to_unsigned(131,8) ,
51269	 => std_logic_vector(to_unsigned(125,8) ,
51270	 => std_logic_vector(to_unsigned(136,8) ,
51271	 => std_logic_vector(to_unsigned(154,8) ,
51272	 => std_logic_vector(to_unsigned(87,8) ,
51273	 => std_logic_vector(to_unsigned(60,8) ,
51274	 => std_logic_vector(to_unsigned(60,8) ,
51275	 => std_logic_vector(to_unsigned(63,8) ,
51276	 => std_logic_vector(to_unsigned(76,8) ,
51277	 => std_logic_vector(to_unsigned(93,8) ,
51278	 => std_logic_vector(to_unsigned(81,8) ,
51279	 => std_logic_vector(to_unsigned(58,8) ,
51280	 => std_logic_vector(to_unsigned(51,8) ,
51281	 => std_logic_vector(to_unsigned(57,8) ,
51282	 => std_logic_vector(to_unsigned(59,8) ,
51283	 => std_logic_vector(to_unsigned(64,8) ,
51284	 => std_logic_vector(to_unsigned(70,8) ,
51285	 => std_logic_vector(to_unsigned(71,8) ,
51286	 => std_logic_vector(to_unsigned(60,8) ,
51287	 => std_logic_vector(to_unsigned(51,8) ,
51288	 => std_logic_vector(to_unsigned(36,8) ,
51289	 => std_logic_vector(to_unsigned(42,8) ,
51290	 => std_logic_vector(to_unsigned(71,8) ,
51291	 => std_logic_vector(to_unsigned(50,8) ,
51292	 => std_logic_vector(to_unsigned(51,8) ,
51293	 => std_logic_vector(to_unsigned(48,8) ,
51294	 => std_logic_vector(to_unsigned(39,8) ,
51295	 => std_logic_vector(to_unsigned(37,8) ,
51296	 => std_logic_vector(to_unsigned(32,8) ,
51297	 => std_logic_vector(to_unsigned(31,8) ,
51298	 => std_logic_vector(to_unsigned(34,8) ,
51299	 => std_logic_vector(to_unsigned(38,8) ,
51300	 => std_logic_vector(to_unsigned(36,8) ,
51301	 => std_logic_vector(to_unsigned(34,8) ,
51302	 => std_logic_vector(to_unsigned(33,8) ,
51303	 => std_logic_vector(to_unsigned(28,8) ,
51304	 => std_logic_vector(to_unsigned(57,8) ,
51305	 => std_logic_vector(to_unsigned(88,8) ,
51306	 => std_logic_vector(to_unsigned(77,8) ,
51307	 => std_logic_vector(to_unsigned(71,8) ,
51308	 => std_logic_vector(to_unsigned(69,8) ,
51309	 => std_logic_vector(to_unsigned(65,8) ,
51310	 => std_logic_vector(to_unsigned(42,8) ,
51311	 => std_logic_vector(to_unsigned(45,8) ,
51312	 => std_logic_vector(to_unsigned(41,8) ,
51313	 => std_logic_vector(to_unsigned(37,8) ,
51314	 => std_logic_vector(to_unsigned(33,8) ,
51315	 => std_logic_vector(to_unsigned(41,8) ,
51316	 => std_logic_vector(to_unsigned(42,8) ,
51317	 => std_logic_vector(to_unsigned(45,8) ,
51318	 => std_logic_vector(to_unsigned(42,8) ,
51319	 => std_logic_vector(to_unsigned(23,8) ,
51320	 => std_logic_vector(to_unsigned(24,8) ,
51321	 => std_logic_vector(to_unsigned(33,8) ,
51322	 => std_logic_vector(to_unsigned(30,8) ,
51323	 => std_logic_vector(to_unsigned(26,8) ,
51324	 => std_logic_vector(to_unsigned(69,8) ,
51325	 => std_logic_vector(to_unsigned(77,8) ,
51326	 => std_logic_vector(to_unsigned(43,8) ,
51327	 => std_logic_vector(to_unsigned(37,8) ,
51328	 => std_logic_vector(to_unsigned(68,8) ,
51329	 => std_logic_vector(to_unsigned(73,8) ,
51330	 => std_logic_vector(to_unsigned(23,8) ,
51331	 => std_logic_vector(to_unsigned(12,8) ,
51332	 => std_logic_vector(to_unsigned(34,8) ,
51333	 => std_logic_vector(to_unsigned(37,8) ,
51334	 => std_logic_vector(to_unsigned(23,8) ,
51335	 => std_logic_vector(to_unsigned(24,8) ,
51336	 => std_logic_vector(to_unsigned(25,8) ,
51337	 => std_logic_vector(to_unsigned(15,8) ,
51338	 => std_logic_vector(to_unsigned(15,8) ,
51339	 => std_logic_vector(to_unsigned(39,8) ,
51340	 => std_logic_vector(to_unsigned(32,8) ,
51341	 => std_logic_vector(to_unsigned(42,8) ,
51342	 => std_logic_vector(to_unsigned(56,8) ,
51343	 => std_logic_vector(to_unsigned(40,8) ,
51344	 => std_logic_vector(to_unsigned(47,8) ,
51345	 => std_logic_vector(to_unsigned(47,8) ,
51346	 => std_logic_vector(to_unsigned(22,8) ,
51347	 => std_logic_vector(to_unsigned(12,8) ,
51348	 => std_logic_vector(to_unsigned(12,8) ,
51349	 => std_logic_vector(to_unsigned(19,8) ,
51350	 => std_logic_vector(to_unsigned(19,8) ,
51351	 => std_logic_vector(to_unsigned(20,8) ,
51352	 => std_logic_vector(to_unsigned(26,8) ,
51353	 => std_logic_vector(to_unsigned(30,8) ,
51354	 => std_logic_vector(to_unsigned(35,8) ,
51355	 => std_logic_vector(to_unsigned(31,8) ,
51356	 => std_logic_vector(to_unsigned(48,8) ,
51357	 => std_logic_vector(to_unsigned(61,8) ,
51358	 => std_logic_vector(to_unsigned(39,8) ,
51359	 => std_logic_vector(to_unsigned(19,8) ,
51360	 => std_logic_vector(to_unsigned(17,8) ,
51361	 => std_logic_vector(to_unsigned(61,8) ,
51362	 => std_logic_vector(to_unsigned(31,8) ,
51363	 => std_logic_vector(to_unsigned(37,8) ,
51364	 => std_logic_vector(to_unsigned(54,8) ,
51365	 => std_logic_vector(to_unsigned(37,8) ,
51366	 => std_logic_vector(to_unsigned(30,8) ,
51367	 => std_logic_vector(to_unsigned(27,8) ,
51368	 => std_logic_vector(to_unsigned(71,8) ,
51369	 => std_logic_vector(to_unsigned(38,8) ,
51370	 => std_logic_vector(to_unsigned(17,8) ,
51371	 => std_logic_vector(to_unsigned(5,8) ,
51372	 => std_logic_vector(to_unsigned(12,8) ,
51373	 => std_logic_vector(to_unsigned(74,8) ,
51374	 => std_logic_vector(to_unsigned(33,8) ,
51375	 => std_logic_vector(to_unsigned(33,8) ,
51376	 => std_logic_vector(to_unsigned(71,8) ,
51377	 => std_logic_vector(to_unsigned(39,8) ,
51378	 => std_logic_vector(to_unsigned(35,8) ,
51379	 => std_logic_vector(to_unsigned(54,8) ,
51380	 => std_logic_vector(to_unsigned(37,8) ,
51381	 => std_logic_vector(to_unsigned(55,8) ,
51382	 => std_logic_vector(to_unsigned(37,8) ,
51383	 => std_logic_vector(to_unsigned(51,8) ,
51384	 => std_logic_vector(to_unsigned(63,8) ,
51385	 => std_logic_vector(to_unsigned(17,8) ,
51386	 => std_logic_vector(to_unsigned(8,8) ,
51387	 => std_logic_vector(to_unsigned(16,8) ,
51388	 => std_logic_vector(to_unsigned(20,8) ,
51389	 => std_logic_vector(to_unsigned(20,8) ,
51390	 => std_logic_vector(to_unsigned(29,8) ,
51391	 => std_logic_vector(to_unsigned(16,8) ,
51392	 => std_logic_vector(to_unsigned(20,8) ,
51393	 => std_logic_vector(to_unsigned(29,8) ,
51394	 => std_logic_vector(to_unsigned(32,8) ,
51395	 => std_logic_vector(to_unsigned(30,8) ,
51396	 => std_logic_vector(to_unsigned(35,8) ,
51397	 => std_logic_vector(to_unsigned(12,8) ,
51398	 => std_logic_vector(to_unsigned(24,8) ,
51399	 => std_logic_vector(to_unsigned(23,8) ,
51400	 => std_logic_vector(to_unsigned(17,8) ,
51401	 => std_logic_vector(to_unsigned(17,8) ,
51402	 => std_logic_vector(to_unsigned(29,8) ,
51403	 => std_logic_vector(to_unsigned(32,8) ,
51404	 => std_logic_vector(to_unsigned(43,8) ,
51405	 => std_logic_vector(to_unsigned(17,8) ,
51406	 => std_logic_vector(to_unsigned(3,8) ,
51407	 => std_logic_vector(to_unsigned(5,8) ,
51408	 => std_logic_vector(to_unsigned(5,8) ,
51409	 => std_logic_vector(to_unsigned(9,8) ,
51410	 => std_logic_vector(to_unsigned(17,8) ,
51411	 => std_logic_vector(to_unsigned(19,8) ,
51412	 => std_logic_vector(to_unsigned(17,8) ,
51413	 => std_logic_vector(to_unsigned(16,8) ,
51414	 => std_logic_vector(to_unsigned(12,8) ,
51415	 => std_logic_vector(to_unsigned(10,8) ,
51416	 => std_logic_vector(to_unsigned(14,8) ,
51417	 => std_logic_vector(to_unsigned(17,8) ,
51418	 => std_logic_vector(to_unsigned(17,8) ,
51419	 => std_logic_vector(to_unsigned(10,8) ,
51420	 => std_logic_vector(to_unsigned(25,8) ,
51421	 => std_logic_vector(to_unsigned(22,8) ,
51422	 => std_logic_vector(to_unsigned(20,8) ,
51423	 => std_logic_vector(to_unsigned(28,8) ,
51424	 => std_logic_vector(to_unsigned(15,8) ,
51425	 => std_logic_vector(to_unsigned(15,8) ,
51426	 => std_logic_vector(to_unsigned(18,8) ,
51427	 => std_logic_vector(to_unsigned(17,8) ,
51428	 => std_logic_vector(to_unsigned(15,8) ,
51429	 => std_logic_vector(to_unsigned(17,8) ,
51430	 => std_logic_vector(to_unsigned(20,8) ,
51431	 => std_logic_vector(to_unsigned(22,8) ,
51432	 => std_logic_vector(to_unsigned(22,8) ,
51433	 => std_logic_vector(to_unsigned(19,8) ,
51434	 => std_logic_vector(to_unsigned(12,8) ,
51435	 => std_logic_vector(to_unsigned(11,8) ,
51436	 => std_logic_vector(to_unsigned(20,8) ,
51437	 => std_logic_vector(to_unsigned(30,8) ,
51438	 => std_logic_vector(to_unsigned(29,8) ,
51439	 => std_logic_vector(to_unsigned(9,8) ,
51440	 => std_logic_vector(to_unsigned(12,8) ,
51441	 => std_logic_vector(to_unsigned(22,8) ,
51442	 => std_logic_vector(to_unsigned(30,8) ,
51443	 => std_logic_vector(to_unsigned(23,8) ,
51444	 => std_logic_vector(to_unsigned(27,8) ,
51445	 => std_logic_vector(to_unsigned(30,8) ,
51446	 => std_logic_vector(to_unsigned(30,8) ,
51447	 => std_logic_vector(to_unsigned(35,8) ,
51448	 => std_logic_vector(to_unsigned(37,8) ,
51449	 => std_logic_vector(to_unsigned(36,8) ,
51450	 => std_logic_vector(to_unsigned(79,8) ,
51451	 => std_logic_vector(to_unsigned(81,8) ,
51452	 => std_logic_vector(to_unsigned(77,8) ,
51453	 => std_logic_vector(to_unsigned(64,8) ,
51454	 => std_logic_vector(to_unsigned(64,8) ,
51455	 => std_logic_vector(to_unsigned(4,8) ,
51456	 => std_logic_vector(to_unsigned(0,8) ,
51457	 => std_logic_vector(to_unsigned(11,8) ,
51458	 => std_logic_vector(to_unsigned(77,8) ,
51459	 => std_logic_vector(to_unsigned(45,8) ,
51460	 => std_logic_vector(to_unsigned(67,8) ,
51461	 => std_logic_vector(to_unsigned(49,8) ,
51462	 => std_logic_vector(to_unsigned(68,8) ,
51463	 => std_logic_vector(to_unsigned(68,8) ,
51464	 => std_logic_vector(to_unsigned(73,8) ,
51465	 => std_logic_vector(to_unsigned(57,8) ,
51466	 => std_logic_vector(to_unsigned(45,8) ,
51467	 => std_logic_vector(to_unsigned(18,8) ,
51468	 => std_logic_vector(to_unsigned(17,8) ,
51469	 => std_logic_vector(to_unsigned(22,8) ,
51470	 => std_logic_vector(to_unsigned(15,8) ,
51471	 => std_logic_vector(to_unsigned(11,8) ,
51472	 => std_logic_vector(to_unsigned(14,8) ,
51473	 => std_logic_vector(to_unsigned(14,8) ,
51474	 => std_logic_vector(to_unsigned(14,8) ,
51475	 => std_logic_vector(to_unsigned(9,8) ,
51476	 => std_logic_vector(to_unsigned(9,8) ,
51477	 => std_logic_vector(to_unsigned(5,8) ,
51478	 => std_logic_vector(to_unsigned(0,8) ,
51479	 => std_logic_vector(to_unsigned(0,8) ,
51480	 => std_logic_vector(to_unsigned(0,8) ,
51481	 => std_logic_vector(to_unsigned(0,8) ,
51482	 => std_logic_vector(to_unsigned(8,8) ,
51483	 => std_logic_vector(to_unsigned(37,8) ,
51484	 => std_logic_vector(to_unsigned(19,8) ,
51485	 => std_logic_vector(to_unsigned(25,8) ,
51486	 => std_logic_vector(to_unsigned(29,8) ,
51487	 => std_logic_vector(to_unsigned(14,8) ,
51488	 => std_logic_vector(to_unsigned(11,8) ,
51489	 => std_logic_vector(to_unsigned(4,8) ,
51490	 => std_logic_vector(to_unsigned(9,8) ,
51491	 => std_logic_vector(to_unsigned(23,8) ,
51492	 => std_logic_vector(to_unsigned(34,8) ,
51493	 => std_logic_vector(to_unsigned(41,8) ,
51494	 => std_logic_vector(to_unsigned(31,8) ,
51495	 => std_logic_vector(to_unsigned(24,8) ,
51496	 => std_logic_vector(to_unsigned(28,8) ,
51497	 => std_logic_vector(to_unsigned(37,8) ,
51498	 => std_logic_vector(to_unsigned(30,8) ,
51499	 => std_logic_vector(to_unsigned(39,8) ,
51500	 => std_logic_vector(to_unsigned(61,8) ,
51501	 => std_logic_vector(to_unsigned(56,8) ,
51502	 => std_logic_vector(to_unsigned(52,8) ,
51503	 => std_logic_vector(to_unsigned(44,8) ,
51504	 => std_logic_vector(to_unsigned(39,8) ,
51505	 => std_logic_vector(to_unsigned(34,8) ,
51506	 => std_logic_vector(to_unsigned(23,8) ,
51507	 => std_logic_vector(to_unsigned(35,8) ,
51508	 => std_logic_vector(to_unsigned(37,8) ,
51509	 => std_logic_vector(to_unsigned(23,8) ,
51510	 => std_logic_vector(to_unsigned(16,8) ,
51511	 => std_logic_vector(to_unsigned(2,8) ,
51512	 => std_logic_vector(to_unsigned(11,8) ,
51513	 => std_logic_vector(to_unsigned(26,8) ,
51514	 => std_logic_vector(to_unsigned(28,8) ,
51515	 => std_logic_vector(to_unsigned(40,8) ,
51516	 => std_logic_vector(to_unsigned(45,8) ,
51517	 => std_logic_vector(to_unsigned(24,8) ,
51518	 => std_logic_vector(to_unsigned(39,8) ,
51519	 => std_logic_vector(to_unsigned(67,8) ,
51520	 => std_logic_vector(to_unsigned(45,8) ,
51521	 => std_logic_vector(to_unsigned(103,8) ,
51522	 => std_logic_vector(to_unsigned(103,8) ,
51523	 => std_logic_vector(to_unsigned(101,8) ,
51524	 => std_logic_vector(to_unsigned(108,8) ,
51525	 => std_logic_vector(to_unsigned(107,8) ,
51526	 => std_logic_vector(to_unsigned(86,8) ,
51527	 => std_logic_vector(to_unsigned(79,8) ,
51528	 => std_logic_vector(to_unsigned(87,8) ,
51529	 => std_logic_vector(to_unsigned(96,8) ,
51530	 => std_logic_vector(to_unsigned(97,8) ,
51531	 => std_logic_vector(to_unsigned(111,8) ,
51532	 => std_logic_vector(to_unsigned(107,8) ,
51533	 => std_logic_vector(to_unsigned(119,8) ,
51534	 => std_logic_vector(to_unsigned(115,8) ,
51535	 => std_logic_vector(to_unsigned(111,8) ,
51536	 => std_logic_vector(to_unsigned(115,8) ,
51537	 => std_logic_vector(to_unsigned(114,8) ,
51538	 => std_logic_vector(to_unsigned(125,8) ,
51539	 => std_logic_vector(to_unsigned(124,8) ,
51540	 => std_logic_vector(to_unsigned(101,8) ,
51541	 => std_logic_vector(to_unsigned(76,8) ,
51542	 => std_logic_vector(to_unsigned(91,8) ,
51543	 => std_logic_vector(to_unsigned(104,8) ,
51544	 => std_logic_vector(to_unsigned(118,8) ,
51545	 => std_logic_vector(to_unsigned(122,8) ,
51546	 => std_logic_vector(to_unsigned(96,8) ,
51547	 => std_logic_vector(to_unsigned(65,8) ,
51548	 => std_logic_vector(to_unsigned(62,8) ,
51549	 => std_logic_vector(to_unsigned(50,8) ,
51550	 => std_logic_vector(to_unsigned(62,8) ,
51551	 => std_logic_vector(to_unsigned(64,8) ,
51552	 => std_logic_vector(to_unsigned(69,8) ,
51553	 => std_logic_vector(to_unsigned(60,8) ,
51554	 => std_logic_vector(to_unsigned(55,8) ,
51555	 => std_logic_vector(to_unsigned(46,8) ,
51556	 => std_logic_vector(to_unsigned(43,8) ,
51557	 => std_logic_vector(to_unsigned(51,8) ,
51558	 => std_logic_vector(to_unsigned(47,8) ,
51559	 => std_logic_vector(to_unsigned(68,8) ,
51560	 => std_logic_vector(to_unsigned(107,8) ,
51561	 => std_logic_vector(to_unsigned(71,8) ,
51562	 => std_logic_vector(to_unsigned(97,8) ,
51563	 => std_logic_vector(to_unsigned(87,8) ,
51564	 => std_logic_vector(to_unsigned(85,8) ,
51565	 => std_logic_vector(to_unsigned(100,8) ,
51566	 => std_logic_vector(to_unsigned(128,8) ,
51567	 => std_logic_vector(to_unsigned(134,8) ,
51568	 => std_logic_vector(to_unsigned(125,8) ,
51569	 => std_logic_vector(to_unsigned(64,8) ,
51570	 => std_logic_vector(to_unsigned(64,8) ,
51571	 => std_logic_vector(to_unsigned(86,8) ,
51572	 => std_logic_vector(to_unsigned(87,8) ,
51573	 => std_logic_vector(to_unsigned(92,8) ,
51574	 => std_logic_vector(to_unsigned(92,8) ,
51575	 => std_logic_vector(to_unsigned(104,8) ,
51576	 => std_logic_vector(to_unsigned(103,8) ,
51577	 => std_logic_vector(to_unsigned(107,8) ,
51578	 => std_logic_vector(to_unsigned(92,8) ,
51579	 => std_logic_vector(to_unsigned(91,8) ,
51580	 => std_logic_vector(to_unsigned(95,8) ,
51581	 => std_logic_vector(to_unsigned(100,8) ,
51582	 => std_logic_vector(to_unsigned(60,8) ,
51583	 => std_logic_vector(to_unsigned(62,8) ,
51584	 => std_logic_vector(to_unsigned(87,8) ,
51585	 => std_logic_vector(to_unsigned(93,8) ,
51586	 => std_logic_vector(to_unsigned(81,8) ,
51587	 => std_logic_vector(to_unsigned(114,8) ,
51588	 => std_logic_vector(to_unsigned(101,8) ,
51589	 => std_logic_vector(to_unsigned(122,8) ,
51590	 => std_logic_vector(to_unsigned(152,8) ,
51591	 => std_logic_vector(to_unsigned(144,8) ,
51592	 => std_logic_vector(to_unsigned(74,8) ,
51593	 => std_logic_vector(to_unsigned(51,8) ,
51594	 => std_logic_vector(to_unsigned(43,8) ,
51595	 => std_logic_vector(to_unsigned(50,8) ,
51596	 => std_logic_vector(to_unsigned(65,8) ,
51597	 => std_logic_vector(to_unsigned(96,8) ,
51598	 => std_logic_vector(to_unsigned(91,8) ,
51599	 => std_logic_vector(to_unsigned(40,8) ,
51600	 => std_logic_vector(to_unsigned(27,8) ,
51601	 => std_logic_vector(to_unsigned(32,8) ,
51602	 => std_logic_vector(to_unsigned(30,8) ,
51603	 => std_logic_vector(to_unsigned(35,8) ,
51604	 => std_logic_vector(to_unsigned(39,8) ,
51605	 => std_logic_vector(to_unsigned(40,8) ,
51606	 => std_logic_vector(to_unsigned(37,8) ,
51607	 => std_logic_vector(to_unsigned(34,8) ,
51608	 => std_logic_vector(to_unsigned(29,8) ,
51609	 => std_logic_vector(to_unsigned(37,8) ,
51610	 => std_logic_vector(to_unsigned(56,8) ,
51611	 => std_logic_vector(to_unsigned(45,8) ,
51612	 => std_logic_vector(to_unsigned(40,8) ,
51613	 => std_logic_vector(to_unsigned(37,8) ,
51614	 => std_logic_vector(to_unsigned(37,8) ,
51615	 => std_logic_vector(to_unsigned(35,8) ,
51616	 => std_logic_vector(to_unsigned(33,8) ,
51617	 => std_logic_vector(to_unsigned(30,8) ,
51618	 => std_logic_vector(to_unsigned(18,8) ,
51619	 => std_logic_vector(to_unsigned(25,8) ,
51620	 => std_logic_vector(to_unsigned(29,8) ,
51621	 => std_logic_vector(to_unsigned(30,8) ,
51622	 => std_logic_vector(to_unsigned(34,8) ,
51623	 => std_logic_vector(to_unsigned(30,8) ,
51624	 => std_logic_vector(to_unsigned(57,8) ,
51625	 => std_logic_vector(to_unsigned(86,8) ,
51626	 => std_logic_vector(to_unsigned(76,8) ,
51627	 => std_logic_vector(to_unsigned(72,8) ,
51628	 => std_logic_vector(to_unsigned(80,8) ,
51629	 => std_logic_vector(to_unsigned(77,8) ,
51630	 => std_logic_vector(to_unsigned(77,8) ,
51631	 => std_logic_vector(to_unsigned(77,8) ,
51632	 => std_logic_vector(to_unsigned(73,8) ,
51633	 => std_logic_vector(to_unsigned(63,8) ,
51634	 => std_logic_vector(to_unsigned(51,8) ,
51635	 => std_logic_vector(to_unsigned(53,8) ,
51636	 => std_logic_vector(to_unsigned(48,8) ,
51637	 => std_logic_vector(to_unsigned(55,8) ,
51638	 => std_logic_vector(to_unsigned(41,8) ,
51639	 => std_logic_vector(to_unsigned(22,8) ,
51640	 => std_logic_vector(to_unsigned(20,8) ,
51641	 => std_logic_vector(to_unsigned(22,8) ,
51642	 => std_logic_vector(to_unsigned(20,8) ,
51643	 => std_logic_vector(to_unsigned(22,8) ,
51644	 => std_logic_vector(to_unsigned(69,8) ,
51645	 => std_logic_vector(to_unsigned(64,8) ,
51646	 => std_logic_vector(to_unsigned(62,8) ,
51647	 => std_logic_vector(to_unsigned(80,8) ,
51648	 => std_logic_vector(to_unsigned(57,8) ,
51649	 => std_logic_vector(to_unsigned(63,8) ,
51650	 => std_logic_vector(to_unsigned(30,8) ,
51651	 => std_logic_vector(to_unsigned(24,8) ,
51652	 => std_logic_vector(to_unsigned(47,8) ,
51653	 => std_logic_vector(to_unsigned(49,8) ,
51654	 => std_logic_vector(to_unsigned(16,8) ,
51655	 => std_logic_vector(to_unsigned(11,8) ,
51656	 => std_logic_vector(to_unsigned(25,8) ,
51657	 => std_logic_vector(to_unsigned(25,8) ,
51658	 => std_logic_vector(to_unsigned(14,8) ,
51659	 => std_logic_vector(to_unsigned(14,8) ,
51660	 => std_logic_vector(to_unsigned(11,8) ,
51661	 => std_logic_vector(to_unsigned(32,8) ,
51662	 => std_logic_vector(to_unsigned(62,8) ,
51663	 => std_logic_vector(to_unsigned(27,8) ,
51664	 => std_logic_vector(to_unsigned(52,8) ,
51665	 => std_logic_vector(to_unsigned(82,8) ,
51666	 => std_logic_vector(to_unsigned(33,8) ,
51667	 => std_logic_vector(to_unsigned(13,8) ,
51668	 => std_logic_vector(to_unsigned(5,8) ,
51669	 => std_logic_vector(to_unsigned(18,8) ,
51670	 => std_logic_vector(to_unsigned(36,8) ,
51671	 => std_logic_vector(to_unsigned(7,8) ,
51672	 => std_logic_vector(to_unsigned(22,8) ,
51673	 => std_logic_vector(to_unsigned(25,8) ,
51674	 => std_logic_vector(to_unsigned(22,8) ,
51675	 => std_logic_vector(to_unsigned(18,8) ,
51676	 => std_logic_vector(to_unsigned(21,8) ,
51677	 => std_logic_vector(to_unsigned(23,8) ,
51678	 => std_logic_vector(to_unsigned(29,8) ,
51679	 => std_logic_vector(to_unsigned(30,8) ,
51680	 => std_logic_vector(to_unsigned(32,8) ,
51681	 => std_logic_vector(to_unsigned(33,8) ,
51682	 => std_logic_vector(to_unsigned(28,8) ,
51683	 => std_logic_vector(to_unsigned(34,8) ,
51684	 => std_logic_vector(to_unsigned(38,8) ,
51685	 => std_logic_vector(to_unsigned(39,8) ,
51686	 => std_logic_vector(to_unsigned(44,8) ,
51687	 => std_logic_vector(to_unsigned(42,8) ,
51688	 => std_logic_vector(to_unsigned(64,8) ,
51689	 => std_logic_vector(to_unsigned(36,8) ,
51690	 => std_logic_vector(to_unsigned(10,8) ,
51691	 => std_logic_vector(to_unsigned(3,8) ,
51692	 => std_logic_vector(to_unsigned(13,8) ,
51693	 => std_logic_vector(to_unsigned(77,8) ,
51694	 => std_logic_vector(to_unsigned(29,8) ,
51695	 => std_logic_vector(to_unsigned(21,8) ,
51696	 => std_logic_vector(to_unsigned(62,8) ,
51697	 => std_logic_vector(to_unsigned(48,8) ,
51698	 => std_logic_vector(to_unsigned(40,8) ,
51699	 => std_logic_vector(to_unsigned(38,8) ,
51700	 => std_logic_vector(to_unsigned(32,8) ,
51701	 => std_logic_vector(to_unsigned(52,8) ,
51702	 => std_logic_vector(to_unsigned(32,8) ,
51703	 => std_logic_vector(to_unsigned(20,8) ,
51704	 => std_logic_vector(to_unsigned(30,8) ,
51705	 => std_logic_vector(to_unsigned(20,8) ,
51706	 => std_logic_vector(to_unsigned(18,8) ,
51707	 => std_logic_vector(to_unsigned(50,8) ,
51708	 => std_logic_vector(to_unsigned(27,8) ,
51709	 => std_logic_vector(to_unsigned(16,8) ,
51710	 => std_logic_vector(to_unsigned(40,8) ,
51711	 => std_logic_vector(to_unsigned(39,8) ,
51712	 => std_logic_vector(to_unsigned(21,8) ,
51713	 => std_logic_vector(to_unsigned(9,8) ,
51714	 => std_logic_vector(to_unsigned(19,8) ,
51715	 => std_logic_vector(to_unsigned(30,8) ,
51716	 => std_logic_vector(to_unsigned(24,8) ,
51717	 => std_logic_vector(to_unsigned(25,8) ,
51718	 => std_logic_vector(to_unsigned(29,8) ,
51719	 => std_logic_vector(to_unsigned(28,8) ,
51720	 => std_logic_vector(to_unsigned(32,8) ,
51721	 => std_logic_vector(to_unsigned(35,8) ,
51722	 => std_logic_vector(to_unsigned(29,8) ,
51723	 => std_logic_vector(to_unsigned(27,8) ,
51724	 => std_logic_vector(to_unsigned(45,8) ,
51725	 => std_logic_vector(to_unsigned(33,8) ,
51726	 => std_logic_vector(to_unsigned(26,8) ,
51727	 => std_logic_vector(to_unsigned(19,8) ,
51728	 => std_logic_vector(to_unsigned(12,8) ,
51729	 => std_logic_vector(to_unsigned(10,8) ,
51730	 => std_logic_vector(to_unsigned(30,8) ,
51731	 => std_logic_vector(to_unsigned(33,8) ,
51732	 => std_logic_vector(to_unsigned(18,8) ,
51733	 => std_logic_vector(to_unsigned(13,8) ,
51734	 => std_logic_vector(to_unsigned(6,8) ,
51735	 => std_logic_vector(to_unsigned(5,8) ,
51736	 => std_logic_vector(to_unsigned(10,8) ,
51737	 => std_logic_vector(to_unsigned(21,8) ,
51738	 => std_logic_vector(to_unsigned(18,8) ,
51739	 => std_logic_vector(to_unsigned(7,8) ,
51740	 => std_logic_vector(to_unsigned(27,8) ,
51741	 => std_logic_vector(to_unsigned(23,8) ,
51742	 => std_logic_vector(to_unsigned(23,8) ,
51743	 => std_logic_vector(to_unsigned(32,8) ,
51744	 => std_logic_vector(to_unsigned(16,8) ,
51745	 => std_logic_vector(to_unsigned(15,8) ,
51746	 => std_logic_vector(to_unsigned(14,8) ,
51747	 => std_logic_vector(to_unsigned(15,8) ,
51748	 => std_logic_vector(to_unsigned(14,8) ,
51749	 => std_logic_vector(to_unsigned(14,8) ,
51750	 => std_logic_vector(to_unsigned(18,8) ,
51751	 => std_logic_vector(to_unsigned(20,8) ,
51752	 => std_logic_vector(to_unsigned(17,8) ,
51753	 => std_logic_vector(to_unsigned(15,8) ,
51754	 => std_logic_vector(to_unsigned(10,8) ,
51755	 => std_logic_vector(to_unsigned(14,8) ,
51756	 => std_logic_vector(to_unsigned(29,8) ,
51757	 => std_logic_vector(to_unsigned(26,8) ,
51758	 => std_logic_vector(to_unsigned(25,8) ,
51759	 => std_logic_vector(to_unsigned(20,8) ,
51760	 => std_logic_vector(to_unsigned(16,8) ,
51761	 => std_logic_vector(to_unsigned(27,8) ,
51762	 => std_logic_vector(to_unsigned(38,8) ,
51763	 => std_logic_vector(to_unsigned(27,8) ,
51764	 => std_logic_vector(to_unsigned(25,8) ,
51765	 => std_logic_vector(to_unsigned(37,8) ,
51766	 => std_logic_vector(to_unsigned(41,8) ,
51767	 => std_logic_vector(to_unsigned(38,8) ,
51768	 => std_logic_vector(to_unsigned(34,8) ,
51769	 => std_logic_vector(to_unsigned(30,8) ,
51770	 => std_logic_vector(to_unsigned(57,8) ,
51771	 => std_logic_vector(to_unsigned(67,8) ,
51772	 => std_logic_vector(to_unsigned(67,8) ,
51773	 => std_logic_vector(to_unsigned(56,8) ,
51774	 => std_logic_vector(to_unsigned(79,8) ,
51775	 => std_logic_vector(to_unsigned(10,8) ,
51776	 => std_logic_vector(to_unsigned(0,8) ,
51777	 => std_logic_vector(to_unsigned(2,8) ,
51778	 => std_logic_vector(to_unsigned(32,8) ,
51779	 => std_logic_vector(to_unsigned(42,8) ,
51780	 => std_logic_vector(to_unsigned(64,8) ,
51781	 => std_logic_vector(to_unsigned(51,8) ,
51782	 => std_logic_vector(to_unsigned(57,8) ,
51783	 => std_logic_vector(to_unsigned(50,8) ,
51784	 => std_logic_vector(to_unsigned(51,8) ,
51785	 => std_logic_vector(to_unsigned(38,8) ,
51786	 => std_logic_vector(to_unsigned(31,8) ,
51787	 => std_logic_vector(to_unsigned(17,8) ,
51788	 => std_logic_vector(to_unsigned(25,8) ,
51789	 => std_logic_vector(to_unsigned(22,8) ,
51790	 => std_logic_vector(to_unsigned(14,8) ,
51791	 => std_logic_vector(to_unsigned(15,8) ,
51792	 => std_logic_vector(to_unsigned(17,8) ,
51793	 => std_logic_vector(to_unsigned(14,8) ,
51794	 => std_logic_vector(to_unsigned(14,8) ,
51795	 => std_logic_vector(to_unsigned(15,8) ,
51796	 => std_logic_vector(to_unsigned(12,8) ,
51797	 => std_logic_vector(to_unsigned(6,8) ,
51798	 => std_logic_vector(to_unsigned(0,8) ,
51799	 => std_logic_vector(to_unsigned(0,8) ,
51800	 => std_logic_vector(to_unsigned(0,8) ,
51801	 => std_logic_vector(to_unsigned(0,8) ,
51802	 => std_logic_vector(to_unsigned(4,8) ,
51803	 => std_logic_vector(to_unsigned(31,8) ,
51804	 => std_logic_vector(to_unsigned(37,8) ,
51805	 => std_logic_vector(to_unsigned(30,8) ,
51806	 => std_logic_vector(to_unsigned(24,8) ,
51807	 => std_logic_vector(to_unsigned(22,8) ,
51808	 => std_logic_vector(to_unsigned(27,8) ,
51809	 => std_logic_vector(to_unsigned(22,8) ,
51810	 => std_logic_vector(to_unsigned(21,8) ,
51811	 => std_logic_vector(to_unsigned(23,8) ,
51812	 => std_logic_vector(to_unsigned(32,8) ,
51813	 => std_logic_vector(to_unsigned(37,8) ,
51814	 => std_logic_vector(to_unsigned(27,8) ,
51815	 => std_logic_vector(to_unsigned(8,8) ,
51816	 => std_logic_vector(to_unsigned(8,8) ,
51817	 => std_logic_vector(to_unsigned(9,8) ,
51818	 => std_logic_vector(to_unsigned(10,8) ,
51819	 => std_logic_vector(to_unsigned(17,8) ,
51820	 => std_logic_vector(to_unsigned(34,8) ,
51821	 => std_logic_vector(to_unsigned(40,8) ,
51822	 => std_logic_vector(to_unsigned(47,8) ,
51823	 => std_logic_vector(to_unsigned(47,8) ,
51824	 => std_logic_vector(to_unsigned(52,8) ,
51825	 => std_logic_vector(to_unsigned(58,8) ,
51826	 => std_logic_vector(to_unsigned(50,8) ,
51827	 => std_logic_vector(to_unsigned(51,8) ,
51828	 => std_logic_vector(to_unsigned(45,8) ,
51829	 => std_logic_vector(to_unsigned(37,8) ,
51830	 => std_logic_vector(to_unsigned(39,8) ,
51831	 => std_logic_vector(to_unsigned(22,8) ,
51832	 => std_logic_vector(to_unsigned(30,8) ,
51833	 => std_logic_vector(to_unsigned(36,8) ,
51834	 => std_logic_vector(to_unsigned(37,8) ,
51835	 => std_logic_vector(to_unsigned(36,8) ,
51836	 => std_logic_vector(to_unsigned(23,8) ,
51837	 => std_logic_vector(to_unsigned(2,8) ,
51838	 => std_logic_vector(to_unsigned(7,8) ,
51839	 => std_logic_vector(to_unsigned(45,8) ,
51840	 => std_logic_vector(to_unsigned(17,8) ,
51841	 => std_logic_vector(to_unsigned(104,8) ,
51842	 => std_logic_vector(to_unsigned(108,8) ,
51843	 => std_logic_vector(to_unsigned(122,8) ,
51844	 => std_logic_vector(to_unsigned(133,8) ,
51845	 => std_logic_vector(to_unsigned(125,8) ,
51846	 => std_logic_vector(to_unsigned(99,8) ,
51847	 => std_logic_vector(to_unsigned(103,8) ,
51848	 => std_logic_vector(to_unsigned(108,8) ,
51849	 => std_logic_vector(to_unsigned(108,8) ,
51850	 => std_logic_vector(to_unsigned(103,8) ,
51851	 => std_logic_vector(to_unsigned(105,8) ,
51852	 => std_logic_vector(to_unsigned(90,8) ,
51853	 => std_logic_vector(to_unsigned(93,8) ,
51854	 => std_logic_vector(to_unsigned(121,8) ,
51855	 => std_logic_vector(to_unsigned(136,8) ,
51856	 => std_logic_vector(to_unsigned(130,8) ,
51857	 => std_logic_vector(to_unsigned(97,8) ,
51858	 => std_logic_vector(to_unsigned(103,8) ,
51859	 => std_logic_vector(to_unsigned(114,8) ,
51860	 => std_logic_vector(to_unsigned(91,8) ,
51861	 => std_logic_vector(to_unsigned(90,8) ,
51862	 => std_logic_vector(to_unsigned(125,8) ,
51863	 => std_logic_vector(to_unsigned(141,8) ,
51864	 => std_logic_vector(to_unsigned(116,8) ,
51865	 => std_logic_vector(to_unsigned(73,8) ,
51866	 => std_logic_vector(to_unsigned(45,8) ,
51867	 => std_logic_vector(to_unsigned(37,8) ,
51868	 => std_logic_vector(to_unsigned(59,8) ,
51869	 => std_logic_vector(to_unsigned(86,8) ,
51870	 => std_logic_vector(to_unsigned(68,8) ,
51871	 => std_logic_vector(to_unsigned(58,8) ,
51872	 => std_logic_vector(to_unsigned(69,8) ,
51873	 => std_logic_vector(to_unsigned(76,8) ,
51874	 => std_logic_vector(to_unsigned(61,8) ,
51875	 => std_logic_vector(to_unsigned(28,8) ,
51876	 => std_logic_vector(to_unsigned(24,8) ,
51877	 => std_logic_vector(to_unsigned(32,8) ,
51878	 => std_logic_vector(to_unsigned(40,8) ,
51879	 => std_logic_vector(to_unsigned(63,8) ,
51880	 => std_logic_vector(to_unsigned(116,8) ,
51881	 => std_logic_vector(to_unsigned(115,8) ,
51882	 => std_logic_vector(to_unsigned(128,8) ,
51883	 => std_logic_vector(to_unsigned(111,8) ,
51884	 => std_logic_vector(to_unsigned(100,8) ,
51885	 => std_logic_vector(to_unsigned(108,8) ,
51886	 => std_logic_vector(to_unsigned(151,8) ,
51887	 => std_logic_vector(to_unsigned(154,8) ,
51888	 => std_logic_vector(to_unsigned(141,8) ,
51889	 => std_logic_vector(to_unsigned(68,8) ,
51890	 => std_logic_vector(to_unsigned(61,8) ,
51891	 => std_logic_vector(to_unsigned(76,8) ,
51892	 => std_logic_vector(to_unsigned(77,8) ,
51893	 => std_logic_vector(to_unsigned(74,8) ,
51894	 => std_logic_vector(to_unsigned(87,8) ,
51895	 => std_logic_vector(to_unsigned(125,8) ,
51896	 => std_logic_vector(to_unsigned(109,8) ,
51897	 => std_logic_vector(to_unsigned(97,8) ,
51898	 => std_logic_vector(to_unsigned(81,8) ,
51899	 => std_logic_vector(to_unsigned(95,8) ,
51900	 => std_logic_vector(to_unsigned(95,8) ,
51901	 => std_logic_vector(to_unsigned(109,8) ,
51902	 => std_logic_vector(to_unsigned(109,8) ,
51903	 => std_logic_vector(to_unsigned(91,8) ,
51904	 => std_logic_vector(to_unsigned(82,8) ,
51905	 => std_logic_vector(to_unsigned(92,8) ,
51906	 => std_logic_vector(to_unsigned(80,8) ,
51907	 => std_logic_vector(to_unsigned(91,8) ,
51908	 => std_logic_vector(to_unsigned(70,8) ,
51909	 => std_logic_vector(to_unsigned(90,8) ,
51910	 => std_logic_vector(to_unsigned(138,8) ,
51911	 => std_logic_vector(to_unsigned(138,8) ,
51912	 => std_logic_vector(to_unsigned(70,8) ,
51913	 => std_logic_vector(to_unsigned(43,8) ,
51914	 => std_logic_vector(to_unsigned(48,8) ,
51915	 => std_logic_vector(to_unsigned(63,8) ,
51916	 => std_logic_vector(to_unsigned(86,8) ,
51917	 => std_logic_vector(to_unsigned(101,8) ,
51918	 => std_logic_vector(to_unsigned(82,8) ,
51919	 => std_logic_vector(to_unsigned(65,8) ,
51920	 => std_logic_vector(to_unsigned(38,8) ,
51921	 => std_logic_vector(to_unsigned(21,8) ,
51922	 => std_logic_vector(to_unsigned(22,8) ,
51923	 => std_logic_vector(to_unsigned(23,8) ,
51924	 => std_logic_vector(to_unsigned(22,8) ,
51925	 => std_logic_vector(to_unsigned(26,8) ,
51926	 => std_logic_vector(to_unsigned(39,8) ,
51927	 => std_logic_vector(to_unsigned(36,8) ,
51928	 => std_logic_vector(to_unsigned(34,8) ,
51929	 => std_logic_vector(to_unsigned(30,8) ,
51930	 => std_logic_vector(to_unsigned(32,8) ,
51931	 => std_logic_vector(to_unsigned(37,8) ,
51932	 => std_logic_vector(to_unsigned(33,8) ,
51933	 => std_logic_vector(to_unsigned(37,8) ,
51934	 => std_logic_vector(to_unsigned(36,8) ,
51935	 => std_logic_vector(to_unsigned(41,8) ,
51936	 => std_logic_vector(to_unsigned(45,8) ,
51937	 => std_logic_vector(to_unsigned(45,8) ,
51938	 => std_logic_vector(to_unsigned(33,8) ,
51939	 => std_logic_vector(to_unsigned(36,8) ,
51940	 => std_logic_vector(to_unsigned(29,8) ,
51941	 => std_logic_vector(to_unsigned(29,8) ,
51942	 => std_logic_vector(to_unsigned(30,8) ,
51943	 => std_logic_vector(to_unsigned(27,8) ,
51944	 => std_logic_vector(to_unsigned(59,8) ,
51945	 => std_logic_vector(to_unsigned(68,8) ,
51946	 => std_logic_vector(to_unsigned(45,8) ,
51947	 => std_logic_vector(to_unsigned(46,8) ,
51948	 => std_logic_vector(to_unsigned(51,8) ,
51949	 => std_logic_vector(to_unsigned(58,8) ,
51950	 => std_logic_vector(to_unsigned(44,8) ,
51951	 => std_logic_vector(to_unsigned(49,8) ,
51952	 => std_logic_vector(to_unsigned(63,8) ,
51953	 => std_logic_vector(to_unsigned(71,8) ,
51954	 => std_logic_vector(to_unsigned(64,8) ,
51955	 => std_logic_vector(to_unsigned(73,8) ,
51956	 => std_logic_vector(to_unsigned(76,8) ,
51957	 => std_logic_vector(to_unsigned(80,8) ,
51958	 => std_logic_vector(to_unsigned(53,8) ,
51959	 => std_logic_vector(to_unsigned(22,8) ,
51960	 => std_logic_vector(to_unsigned(18,8) ,
51961	 => std_logic_vector(to_unsigned(20,8) ,
51962	 => std_logic_vector(to_unsigned(23,8) ,
51963	 => std_logic_vector(to_unsigned(20,8) ,
51964	 => std_logic_vector(to_unsigned(67,8) ,
51965	 => std_logic_vector(to_unsigned(88,8) ,
51966	 => std_logic_vector(to_unsigned(74,8) ,
51967	 => std_logic_vector(to_unsigned(53,8) ,
51968	 => std_logic_vector(to_unsigned(31,8) ,
51969	 => std_logic_vector(to_unsigned(65,8) ,
51970	 => std_logic_vector(to_unsigned(84,8) ,
51971	 => std_logic_vector(to_unsigned(51,8) ,
51972	 => std_logic_vector(to_unsigned(55,8) ,
51973	 => std_logic_vector(to_unsigned(54,8) ,
51974	 => std_logic_vector(to_unsigned(27,8) ,
51975	 => std_logic_vector(to_unsigned(16,8) ,
51976	 => std_logic_vector(to_unsigned(22,8) ,
51977	 => std_logic_vector(to_unsigned(27,8) ,
51978	 => std_logic_vector(to_unsigned(14,8) ,
51979	 => std_logic_vector(to_unsigned(9,8) ,
51980	 => std_logic_vector(to_unsigned(8,8) ,
51981	 => std_logic_vector(to_unsigned(41,8) ,
51982	 => std_logic_vector(to_unsigned(68,8) ,
51983	 => std_logic_vector(to_unsigned(22,8) ,
51984	 => std_logic_vector(to_unsigned(32,8) ,
51985	 => std_logic_vector(to_unsigned(73,8) ,
51986	 => std_logic_vector(to_unsigned(35,8) ,
51987	 => std_logic_vector(to_unsigned(13,8) ,
51988	 => std_logic_vector(to_unsigned(7,8) ,
51989	 => std_logic_vector(to_unsigned(18,8) ,
51990	 => std_logic_vector(to_unsigned(63,8) ,
51991	 => std_logic_vector(to_unsigned(33,8) ,
51992	 => std_logic_vector(to_unsigned(50,8) ,
51993	 => std_logic_vector(to_unsigned(51,8) ,
51994	 => std_logic_vector(to_unsigned(45,8) ,
51995	 => std_logic_vector(to_unsigned(29,8) ,
51996	 => std_logic_vector(to_unsigned(50,8) ,
51997	 => std_logic_vector(to_unsigned(30,8) ,
51998	 => std_logic_vector(to_unsigned(10,8) ,
51999	 => std_logic_vector(to_unsigned(8,8) ,
52000	 => std_logic_vector(to_unsigned(7,8) ,
52001	 => std_logic_vector(to_unsigned(22,8) ,
52002	 => std_logic_vector(to_unsigned(12,8) ,
52003	 => std_logic_vector(to_unsigned(9,8) ,
52004	 => std_logic_vector(to_unsigned(15,8) ,
52005	 => std_logic_vector(to_unsigned(16,8) ,
52006	 => std_logic_vector(to_unsigned(19,8) ,
52007	 => std_logic_vector(to_unsigned(24,8) ,
52008	 => std_logic_vector(to_unsigned(25,8) ,
52009	 => std_logic_vector(to_unsigned(29,8) ,
52010	 => std_logic_vector(to_unsigned(30,8) ,
52011	 => std_logic_vector(to_unsigned(18,8) ,
52012	 => std_logic_vector(to_unsigned(25,8) ,
52013	 => std_logic_vector(to_unsigned(66,8) ,
52014	 => std_logic_vector(to_unsigned(45,8) ,
52015	 => std_logic_vector(to_unsigned(45,8) ,
52016	 => std_logic_vector(to_unsigned(61,8) ,
52017	 => std_logic_vector(to_unsigned(49,8) ,
52018	 => std_logic_vector(to_unsigned(41,8) ,
52019	 => std_logic_vector(to_unsigned(23,8) ,
52020	 => std_logic_vector(to_unsigned(16,8) ,
52021	 => std_logic_vector(to_unsigned(24,8) ,
52022	 => std_logic_vector(to_unsigned(19,8) ,
52023	 => std_logic_vector(to_unsigned(27,8) ,
52024	 => std_logic_vector(to_unsigned(31,8) ,
52025	 => std_logic_vector(to_unsigned(31,8) ,
52026	 => std_logic_vector(to_unsigned(41,8) ,
52027	 => std_logic_vector(to_unsigned(37,8) ,
52028	 => std_logic_vector(to_unsigned(21,8) ,
52029	 => std_logic_vector(to_unsigned(23,8) ,
52030	 => std_logic_vector(to_unsigned(38,8) ,
52031	 => std_logic_vector(to_unsigned(45,8) ,
52032	 => std_logic_vector(to_unsigned(18,8) ,
52033	 => std_logic_vector(to_unsigned(6,8) ,
52034	 => std_logic_vector(to_unsigned(11,8) ,
52035	 => std_logic_vector(to_unsigned(22,8) ,
52036	 => std_logic_vector(to_unsigned(24,8) ,
52037	 => std_logic_vector(to_unsigned(23,8) ,
52038	 => std_logic_vector(to_unsigned(21,8) ,
52039	 => std_logic_vector(to_unsigned(19,8) ,
52040	 => std_logic_vector(to_unsigned(22,8) ,
52041	 => std_logic_vector(to_unsigned(22,8) ,
52042	 => std_logic_vector(to_unsigned(22,8) ,
52043	 => std_logic_vector(to_unsigned(19,8) ,
52044	 => std_logic_vector(to_unsigned(23,8) ,
52045	 => std_logic_vector(to_unsigned(31,8) ,
52046	 => std_logic_vector(to_unsigned(37,8) ,
52047	 => std_logic_vector(to_unsigned(35,8) ,
52048	 => std_logic_vector(to_unsigned(30,8) ,
52049	 => std_logic_vector(to_unsigned(29,8) ,
52050	 => std_logic_vector(to_unsigned(36,8) ,
52051	 => std_logic_vector(to_unsigned(29,8) ,
52052	 => std_logic_vector(to_unsigned(23,8) ,
52053	 => std_logic_vector(to_unsigned(26,8) ,
52054	 => std_logic_vector(to_unsigned(18,8) ,
52055	 => std_logic_vector(to_unsigned(14,8) ,
52056	 => std_logic_vector(to_unsigned(13,8) ,
52057	 => std_logic_vector(to_unsigned(17,8) ,
52058	 => std_logic_vector(to_unsigned(26,8) ,
52059	 => std_logic_vector(to_unsigned(17,8) ,
52060	 => std_logic_vector(to_unsigned(17,8) ,
52061	 => std_logic_vector(to_unsigned(13,8) ,
52062	 => std_logic_vector(to_unsigned(32,8) ,
52063	 => std_logic_vector(to_unsigned(33,8) ,
52064	 => std_logic_vector(to_unsigned(16,8) ,
52065	 => std_logic_vector(to_unsigned(14,8) ,
52066	 => std_logic_vector(to_unsigned(12,8) ,
52067	 => std_logic_vector(to_unsigned(13,8) ,
52068	 => std_logic_vector(to_unsigned(14,8) ,
52069	 => std_logic_vector(to_unsigned(15,8) ,
52070	 => std_logic_vector(to_unsigned(17,8) ,
52071	 => std_logic_vector(to_unsigned(18,8) ,
52072	 => std_logic_vector(to_unsigned(14,8) ,
52073	 => std_logic_vector(to_unsigned(13,8) ,
52074	 => std_logic_vector(to_unsigned(9,8) ,
52075	 => std_logic_vector(to_unsigned(13,8) ,
52076	 => std_logic_vector(to_unsigned(26,8) ,
52077	 => std_logic_vector(to_unsigned(17,8) ,
52078	 => std_logic_vector(to_unsigned(11,8) ,
52079	 => std_logic_vector(to_unsigned(21,8) ,
52080	 => std_logic_vector(to_unsigned(20,8) ,
52081	 => std_logic_vector(to_unsigned(24,8) ,
52082	 => std_logic_vector(to_unsigned(24,8) ,
52083	 => std_logic_vector(to_unsigned(20,8) ,
52084	 => std_logic_vector(to_unsigned(30,8) ,
52085	 => std_logic_vector(to_unsigned(39,8) ,
52086	 => std_logic_vector(to_unsigned(33,8) ,
52087	 => std_logic_vector(to_unsigned(31,8) ,
52088	 => std_logic_vector(to_unsigned(31,8) ,
52089	 => std_logic_vector(to_unsigned(25,8) ,
52090	 => std_logic_vector(to_unsigned(27,8) ,
52091	 => std_logic_vector(to_unsigned(37,8) ,
52092	 => std_logic_vector(to_unsigned(50,8) ,
52093	 => std_logic_vector(to_unsigned(38,8) ,
52094	 => std_logic_vector(to_unsigned(41,8) ,
52095	 => std_logic_vector(to_unsigned(18,8) ,
52096	 => std_logic_vector(to_unsigned(1,8) ,
52097	 => std_logic_vector(to_unsigned(0,8) ,
52098	 => std_logic_vector(to_unsigned(5,8) ,
52099	 => std_logic_vector(to_unsigned(32,8) ,
52100	 => std_logic_vector(to_unsigned(42,8) ,
52101	 => std_logic_vector(to_unsigned(50,8) ,
52102	 => std_logic_vector(to_unsigned(70,8) ,
52103	 => std_logic_vector(to_unsigned(63,8) ,
52104	 => std_logic_vector(to_unsigned(53,8) ,
52105	 => std_logic_vector(to_unsigned(39,8) ,
52106	 => std_logic_vector(to_unsigned(25,8) ,
52107	 => std_logic_vector(to_unsigned(14,8) ,
52108	 => std_logic_vector(to_unsigned(17,8) ,
52109	 => std_logic_vector(to_unsigned(19,8) ,
52110	 => std_logic_vector(to_unsigned(12,8) ,
52111	 => std_logic_vector(to_unsigned(12,8) ,
52112	 => std_logic_vector(to_unsigned(13,8) ,
52113	 => std_logic_vector(to_unsigned(13,8) ,
52114	 => std_logic_vector(to_unsigned(13,8) ,
52115	 => std_logic_vector(to_unsigned(15,8) ,
52116	 => std_logic_vector(to_unsigned(14,8) ,
52117	 => std_logic_vector(to_unsigned(7,8) ,
52118	 => std_logic_vector(to_unsigned(1,8) ,
52119	 => std_logic_vector(to_unsigned(0,8) ,
52120	 => std_logic_vector(to_unsigned(0,8) ,
52121	 => std_logic_vector(to_unsigned(0,8) ,
52122	 => std_logic_vector(to_unsigned(1,8) ,
52123	 => std_logic_vector(to_unsigned(13,8) ,
52124	 => std_logic_vector(to_unsigned(17,8) ,
52125	 => std_logic_vector(to_unsigned(12,8) ,
52126	 => std_logic_vector(to_unsigned(18,8) ,
52127	 => std_logic_vector(to_unsigned(15,8) ,
52128	 => std_logic_vector(to_unsigned(19,8) ,
52129	 => std_logic_vector(to_unsigned(20,8) ,
52130	 => std_logic_vector(to_unsigned(22,8) ,
52131	 => std_logic_vector(to_unsigned(28,8) ,
52132	 => std_logic_vector(to_unsigned(30,8) ,
52133	 => std_logic_vector(to_unsigned(30,8) ,
52134	 => std_logic_vector(to_unsigned(25,8) ,
52135	 => std_logic_vector(to_unsigned(13,8) ,
52136	 => std_logic_vector(to_unsigned(11,8) ,
52137	 => std_logic_vector(to_unsigned(9,8) ,
52138	 => std_logic_vector(to_unsigned(4,8) ,
52139	 => std_logic_vector(to_unsigned(28,8) ,
52140	 => std_logic_vector(to_unsigned(34,8) ,
52141	 => std_logic_vector(to_unsigned(17,8) ,
52142	 => std_logic_vector(to_unsigned(18,8) ,
52143	 => std_logic_vector(to_unsigned(16,8) ,
52144	 => std_logic_vector(to_unsigned(18,8) ,
52145	 => std_logic_vector(to_unsigned(24,8) ,
52146	 => std_logic_vector(to_unsigned(20,8) ,
52147	 => std_logic_vector(to_unsigned(41,8) ,
52148	 => std_logic_vector(to_unsigned(33,8) ,
52149	 => std_logic_vector(to_unsigned(20,8) ,
52150	 => std_logic_vector(to_unsigned(19,8) ,
52151	 => std_logic_vector(to_unsigned(19,8) ,
52152	 => std_logic_vector(to_unsigned(30,8) ,
52153	 => std_logic_vector(to_unsigned(40,8) ,
52154	 => std_logic_vector(to_unsigned(48,8) ,
52155	 => std_logic_vector(to_unsigned(51,8) ,
52156	 => std_logic_vector(to_unsigned(53,8) ,
52157	 => std_logic_vector(to_unsigned(41,8) ,
52158	 => std_logic_vector(to_unsigned(46,8) ,
52159	 => std_logic_vector(to_unsigned(60,8) ,
52160	 => std_logic_vector(to_unsigned(40,8) ,
52161	 => std_logic_vector(to_unsigned(114,8) ,
52162	 => std_logic_vector(to_unsigned(128,8) ,
52163	 => std_logic_vector(to_unsigned(146,8) ,
52164	 => std_logic_vector(to_unsigned(146,8) ,
52165	 => std_logic_vector(to_unsigned(124,8) ,
52166	 => std_logic_vector(to_unsigned(97,8) ,
52167	 => std_logic_vector(to_unsigned(114,8) ,
52168	 => std_logic_vector(to_unsigned(124,8) ,
52169	 => std_logic_vector(to_unsigned(127,8) ,
52170	 => std_logic_vector(to_unsigned(122,8) ,
52171	 => std_logic_vector(to_unsigned(109,8) ,
52172	 => std_logic_vector(to_unsigned(108,8) ,
52173	 => std_logic_vector(to_unsigned(103,8) ,
52174	 => std_logic_vector(to_unsigned(133,8) ,
52175	 => std_logic_vector(to_unsigned(147,8) ,
52176	 => std_logic_vector(to_unsigned(131,8) ,
52177	 => std_logic_vector(to_unsigned(92,8) ,
52178	 => std_logic_vector(to_unsigned(87,8) ,
52179	 => std_logic_vector(to_unsigned(109,8) ,
52180	 => std_logic_vector(to_unsigned(107,8) ,
52181	 => std_logic_vector(to_unsigned(96,8) ,
52182	 => std_logic_vector(to_unsigned(99,8) ,
52183	 => std_logic_vector(to_unsigned(97,8) ,
52184	 => std_logic_vector(to_unsigned(53,8) ,
52185	 => std_logic_vector(to_unsigned(41,8) ,
52186	 => std_logic_vector(to_unsigned(45,8) ,
52187	 => std_logic_vector(to_unsigned(52,8) ,
52188	 => std_logic_vector(to_unsigned(62,8) ,
52189	 => std_logic_vector(to_unsigned(78,8) ,
52190	 => std_logic_vector(to_unsigned(58,8) ,
52191	 => std_logic_vector(to_unsigned(36,8) ,
52192	 => std_logic_vector(to_unsigned(55,8) ,
52193	 => std_logic_vector(to_unsigned(70,8) ,
52194	 => std_logic_vector(to_unsigned(51,8) ,
52195	 => std_logic_vector(to_unsigned(23,8) ,
52196	 => std_logic_vector(to_unsigned(20,8) ,
52197	 => std_logic_vector(to_unsigned(26,8) ,
52198	 => std_logic_vector(to_unsigned(24,8) ,
52199	 => std_logic_vector(to_unsigned(32,8) ,
52200	 => std_logic_vector(to_unsigned(47,8) ,
52201	 => std_logic_vector(to_unsigned(65,8) ,
52202	 => std_logic_vector(to_unsigned(74,8) ,
52203	 => std_logic_vector(to_unsigned(85,8) ,
52204	 => std_logic_vector(to_unsigned(86,8) ,
52205	 => std_logic_vector(to_unsigned(105,8) ,
52206	 => std_logic_vector(to_unsigned(119,8) ,
52207	 => std_logic_vector(to_unsigned(124,8) ,
52208	 => std_logic_vector(to_unsigned(149,8) ,
52209	 => std_logic_vector(to_unsigned(74,8) ,
52210	 => std_logic_vector(to_unsigned(60,8) ,
52211	 => std_logic_vector(to_unsigned(81,8) ,
52212	 => std_logic_vector(to_unsigned(74,8) ,
52213	 => std_logic_vector(to_unsigned(64,8) ,
52214	 => std_logic_vector(to_unsigned(79,8) ,
52215	 => std_logic_vector(to_unsigned(95,8) ,
52216	 => std_logic_vector(to_unsigned(91,8) ,
52217	 => std_logic_vector(to_unsigned(95,8) ,
52218	 => std_logic_vector(to_unsigned(96,8) ,
52219	 => std_logic_vector(to_unsigned(115,8) ,
52220	 => std_logic_vector(to_unsigned(108,8) ,
52221	 => std_logic_vector(to_unsigned(111,8) ,
52222	 => std_logic_vector(to_unsigned(134,8) ,
52223	 => std_logic_vector(to_unsigned(91,8) ,
52224	 => std_logic_vector(to_unsigned(71,8) ,
52225	 => std_logic_vector(to_unsigned(105,8) ,
52226	 => std_logic_vector(to_unsigned(109,8) ,
52227	 => std_logic_vector(to_unsigned(99,8) ,
52228	 => std_logic_vector(to_unsigned(90,8) ,
52229	 => std_logic_vector(to_unsigned(97,8) ,
52230	 => std_logic_vector(to_unsigned(128,8) ,
52231	 => std_logic_vector(to_unsigned(133,8) ,
52232	 => std_logic_vector(to_unsigned(76,8) ,
52233	 => std_logic_vector(to_unsigned(43,8) ,
52234	 => std_logic_vector(to_unsigned(72,8) ,
52235	 => std_logic_vector(to_unsigned(86,8) ,
52236	 => std_logic_vector(to_unsigned(91,8) ,
52237	 => std_logic_vector(to_unsigned(92,8) ,
52238	 => std_logic_vector(to_unsigned(84,8) ,
52239	 => std_logic_vector(to_unsigned(88,8) ,
52240	 => std_logic_vector(to_unsigned(53,8) ,
52241	 => std_logic_vector(to_unsigned(23,8) ,
52242	 => std_logic_vector(to_unsigned(24,8) ,
52243	 => std_logic_vector(to_unsigned(22,8) ,
52244	 => std_logic_vector(to_unsigned(23,8) ,
52245	 => std_logic_vector(to_unsigned(23,8) ,
52246	 => std_logic_vector(to_unsigned(40,8) ,
52247	 => std_logic_vector(to_unsigned(37,8) ,
52248	 => std_logic_vector(to_unsigned(32,8) ,
52249	 => std_logic_vector(to_unsigned(34,8) ,
52250	 => std_logic_vector(to_unsigned(30,8) ,
52251	 => std_logic_vector(to_unsigned(32,8) ,
52252	 => std_logic_vector(to_unsigned(32,8) ,
52253	 => std_logic_vector(to_unsigned(38,8) ,
52254	 => std_logic_vector(to_unsigned(37,8) ,
52255	 => std_logic_vector(to_unsigned(43,8) ,
52256	 => std_logic_vector(to_unsigned(57,8) ,
52257	 => std_logic_vector(to_unsigned(72,8) ,
52258	 => std_logic_vector(to_unsigned(64,8) ,
52259	 => std_logic_vector(to_unsigned(49,8) ,
52260	 => std_logic_vector(to_unsigned(38,8) ,
52261	 => std_logic_vector(to_unsigned(34,8) ,
52262	 => std_logic_vector(to_unsigned(30,8) ,
52263	 => std_logic_vector(to_unsigned(29,8) ,
52264	 => std_logic_vector(to_unsigned(52,8) ,
52265	 => std_logic_vector(to_unsigned(62,8) ,
52266	 => std_logic_vector(to_unsigned(45,8) ,
52267	 => std_logic_vector(to_unsigned(50,8) ,
52268	 => std_logic_vector(to_unsigned(42,8) ,
52269	 => std_logic_vector(to_unsigned(48,8) ,
52270	 => std_logic_vector(to_unsigned(35,8) ,
52271	 => std_logic_vector(to_unsigned(35,8) ,
52272	 => std_logic_vector(to_unsigned(37,8) ,
52273	 => std_logic_vector(to_unsigned(36,8) ,
52274	 => std_logic_vector(to_unsigned(30,8) ,
52275	 => std_logic_vector(to_unsigned(34,8) ,
52276	 => std_logic_vector(to_unsigned(39,8) ,
52277	 => std_logic_vector(to_unsigned(54,8) ,
52278	 => std_logic_vector(to_unsigned(38,8) ,
52279	 => std_logic_vector(to_unsigned(17,8) ,
52280	 => std_logic_vector(to_unsigned(17,8) ,
52281	 => std_logic_vector(to_unsigned(22,8) ,
52282	 => std_logic_vector(to_unsigned(23,8) ,
52283	 => std_logic_vector(to_unsigned(25,8) ,
52284	 => std_logic_vector(to_unsigned(66,8) ,
52285	 => std_logic_vector(to_unsigned(84,8) ,
52286	 => std_logic_vector(to_unsigned(45,8) ,
52287	 => std_logic_vector(to_unsigned(35,8) ,
52288	 => std_logic_vector(to_unsigned(36,8) ,
52289	 => std_logic_vector(to_unsigned(63,8) ,
52290	 => std_logic_vector(to_unsigned(63,8) ,
52291	 => std_logic_vector(to_unsigned(35,8) ,
52292	 => std_logic_vector(to_unsigned(41,8) ,
52293	 => std_logic_vector(to_unsigned(51,8) ,
52294	 => std_logic_vector(to_unsigned(46,8) ,
52295	 => std_logic_vector(to_unsigned(32,8) ,
52296	 => std_logic_vector(to_unsigned(33,8) ,
52297	 => std_logic_vector(to_unsigned(26,8) ,
52298	 => std_logic_vector(to_unsigned(13,8) ,
52299	 => std_logic_vector(to_unsigned(14,8) ,
52300	 => std_logic_vector(to_unsigned(25,8) ,
52301	 => std_logic_vector(to_unsigned(44,8) ,
52302	 => std_logic_vector(to_unsigned(66,8) ,
52303	 => std_logic_vector(to_unsigned(37,8) ,
52304	 => std_logic_vector(to_unsigned(49,8) ,
52305	 => std_logic_vector(to_unsigned(84,8) ,
52306	 => std_logic_vector(to_unsigned(39,8) ,
52307	 => std_logic_vector(to_unsigned(11,8) ,
52308	 => std_logic_vector(to_unsigned(5,8) ,
52309	 => std_logic_vector(to_unsigned(17,8) ,
52310	 => std_logic_vector(to_unsigned(60,8) ,
52311	 => std_logic_vector(to_unsigned(42,8) ,
52312	 => std_logic_vector(to_unsigned(55,8) ,
52313	 => std_logic_vector(to_unsigned(51,8) ,
52314	 => std_logic_vector(to_unsigned(59,8) ,
52315	 => std_logic_vector(to_unsigned(51,8) ,
52316	 => std_logic_vector(to_unsigned(67,8) ,
52317	 => std_logic_vector(to_unsigned(44,8) ,
52318	 => std_logic_vector(to_unsigned(11,8) ,
52319	 => std_logic_vector(to_unsigned(6,8) ,
52320	 => std_logic_vector(to_unsigned(8,8) ,
52321	 => std_logic_vector(to_unsigned(48,8) ,
52322	 => std_logic_vector(to_unsigned(27,8) ,
52323	 => std_logic_vector(to_unsigned(17,8) ,
52324	 => std_logic_vector(to_unsigned(24,8) ,
52325	 => std_logic_vector(to_unsigned(19,8) ,
52326	 => std_logic_vector(to_unsigned(17,8) ,
52327	 => std_logic_vector(to_unsigned(16,8) ,
52328	 => std_logic_vector(to_unsigned(18,8) ,
52329	 => std_logic_vector(to_unsigned(13,8) ,
52330	 => std_logic_vector(to_unsigned(12,8) ,
52331	 => std_logic_vector(to_unsigned(13,8) ,
52332	 => std_logic_vector(to_unsigned(15,8) ,
52333	 => std_logic_vector(to_unsigned(17,8) ,
52334	 => std_logic_vector(to_unsigned(15,8) ,
52335	 => std_logic_vector(to_unsigned(23,8) ,
52336	 => std_logic_vector(to_unsigned(43,8) ,
52337	 => std_logic_vector(to_unsigned(43,8) ,
52338	 => std_logic_vector(to_unsigned(39,8) ,
52339	 => std_logic_vector(to_unsigned(31,8) ,
52340	 => std_logic_vector(to_unsigned(28,8) ,
52341	 => std_logic_vector(to_unsigned(33,8) ,
52342	 => std_logic_vector(to_unsigned(28,8) ,
52343	 => std_logic_vector(to_unsigned(28,8) ,
52344	 => std_logic_vector(to_unsigned(28,8) ,
52345	 => std_logic_vector(to_unsigned(35,8) ,
52346	 => std_logic_vector(to_unsigned(37,8) ,
52347	 => std_logic_vector(to_unsigned(35,8) ,
52348	 => std_logic_vector(to_unsigned(28,8) ,
52349	 => std_logic_vector(to_unsigned(23,8) ,
52350	 => std_logic_vector(to_unsigned(32,8) ,
52351	 => std_logic_vector(to_unsigned(30,8) ,
52352	 => std_logic_vector(to_unsigned(28,8) ,
52353	 => std_logic_vector(to_unsigned(25,8) ,
52354	 => std_logic_vector(to_unsigned(16,8) ,
52355	 => std_logic_vector(to_unsigned(17,8) ,
52356	 => std_logic_vector(to_unsigned(26,8) ,
52357	 => std_logic_vector(to_unsigned(49,8) ,
52358	 => std_logic_vector(to_unsigned(61,8) ,
52359	 => std_logic_vector(to_unsigned(35,8) ,
52360	 => std_logic_vector(to_unsigned(20,8) ,
52361	 => std_logic_vector(to_unsigned(32,8) ,
52362	 => std_logic_vector(to_unsigned(31,8) ,
52363	 => std_logic_vector(to_unsigned(22,8) ,
52364	 => std_logic_vector(to_unsigned(13,8) ,
52365	 => std_logic_vector(to_unsigned(12,8) ,
52366	 => std_logic_vector(to_unsigned(15,8) ,
52367	 => std_logic_vector(to_unsigned(14,8) ,
52368	 => std_logic_vector(to_unsigned(21,8) ,
52369	 => std_logic_vector(to_unsigned(22,8) ,
52370	 => std_logic_vector(to_unsigned(19,8) ,
52371	 => std_logic_vector(to_unsigned(22,8) ,
52372	 => std_logic_vector(to_unsigned(27,8) ,
52373	 => std_logic_vector(to_unsigned(28,8) ,
52374	 => std_logic_vector(to_unsigned(29,8) ,
52375	 => std_logic_vector(to_unsigned(27,8) ,
52376	 => std_logic_vector(to_unsigned(20,8) ,
52377	 => std_logic_vector(to_unsigned(15,8) ,
52378	 => std_logic_vector(to_unsigned(29,8) ,
52379	 => std_logic_vector(to_unsigned(41,8) ,
52380	 => std_logic_vector(to_unsigned(18,8) ,
52381	 => std_logic_vector(to_unsigned(18,8) ,
52382	 => std_logic_vector(to_unsigned(32,8) ,
52383	 => std_logic_vector(to_unsigned(25,8) ,
52384	 => std_logic_vector(to_unsigned(17,8) ,
52385	 => std_logic_vector(to_unsigned(16,8) ,
52386	 => std_logic_vector(to_unsigned(15,8) ,
52387	 => std_logic_vector(to_unsigned(14,8) ,
52388	 => std_logic_vector(to_unsigned(16,8) ,
52389	 => std_logic_vector(to_unsigned(12,8) ,
52390	 => std_logic_vector(to_unsigned(15,8) ,
52391	 => std_logic_vector(to_unsigned(18,8) ,
52392	 => std_logic_vector(to_unsigned(15,8) ,
52393	 => std_logic_vector(to_unsigned(25,8) ,
52394	 => std_logic_vector(to_unsigned(15,8) ,
52395	 => std_logic_vector(to_unsigned(10,8) ,
52396	 => std_logic_vector(to_unsigned(21,8) ,
52397	 => std_logic_vector(to_unsigned(12,8) ,
52398	 => std_logic_vector(to_unsigned(16,8) ,
52399	 => std_logic_vector(to_unsigned(32,8) ,
52400	 => std_logic_vector(to_unsigned(29,8) ,
52401	 => std_logic_vector(to_unsigned(16,8) ,
52402	 => std_logic_vector(to_unsigned(10,8) ,
52403	 => std_logic_vector(to_unsigned(25,8) ,
52404	 => std_logic_vector(to_unsigned(30,8) ,
52405	 => std_logic_vector(to_unsigned(30,8) ,
52406	 => std_logic_vector(to_unsigned(30,8) ,
52407	 => std_logic_vector(to_unsigned(27,8) ,
52408	 => std_logic_vector(to_unsigned(24,8) ,
52409	 => std_logic_vector(to_unsigned(32,8) ,
52410	 => std_logic_vector(to_unsigned(42,8) ,
52411	 => std_logic_vector(to_unsigned(54,8) ,
52412	 => std_logic_vector(to_unsigned(79,8) ,
52413	 => std_logic_vector(to_unsigned(71,8) ,
52414	 => std_logic_vector(to_unsigned(60,8) ,
52415	 => std_logic_vector(to_unsigned(35,8) ,
52416	 => std_logic_vector(to_unsigned(4,8) ,
52417	 => std_logic_vector(to_unsigned(0,8) ,
52418	 => std_logic_vector(to_unsigned(1,8) ,
52419	 => std_logic_vector(to_unsigned(18,8) ,
52420	 => std_logic_vector(to_unsigned(32,8) ,
52421	 => std_logic_vector(to_unsigned(32,8) ,
52422	 => std_logic_vector(to_unsigned(45,8) ,
52423	 => std_logic_vector(to_unsigned(51,8) ,
52424	 => std_logic_vector(to_unsigned(47,8) ,
52425	 => std_logic_vector(to_unsigned(55,8) ,
52426	 => std_logic_vector(to_unsigned(22,8) ,
52427	 => std_logic_vector(to_unsigned(12,8) ,
52428	 => std_logic_vector(to_unsigned(18,8) ,
52429	 => std_logic_vector(to_unsigned(19,8) ,
52430	 => std_logic_vector(to_unsigned(16,8) ,
52431	 => std_logic_vector(to_unsigned(12,8) ,
52432	 => std_logic_vector(to_unsigned(12,8) ,
52433	 => std_logic_vector(to_unsigned(13,8) ,
52434	 => std_logic_vector(to_unsigned(10,8) ,
52435	 => std_logic_vector(to_unsigned(8,8) ,
52436	 => std_logic_vector(to_unsigned(10,8) ,
52437	 => std_logic_vector(to_unsigned(8,8) ,
52438	 => std_logic_vector(to_unsigned(2,8) ,
52439	 => std_logic_vector(to_unsigned(0,8) ,
52440	 => std_logic_vector(to_unsigned(0,8) ,
52441	 => std_logic_vector(to_unsigned(0,8) ,
52442	 => std_logic_vector(to_unsigned(1,8) ,
52443	 => std_logic_vector(to_unsigned(9,8) ,
52444	 => std_logic_vector(to_unsigned(11,8) ,
52445	 => std_logic_vector(to_unsigned(10,8) ,
52446	 => std_logic_vector(to_unsigned(15,8) ,
52447	 => std_logic_vector(to_unsigned(10,8) ,
52448	 => std_logic_vector(to_unsigned(5,8) ,
52449	 => std_logic_vector(to_unsigned(4,8) ,
52450	 => std_logic_vector(to_unsigned(10,8) ,
52451	 => std_logic_vector(to_unsigned(25,8) ,
52452	 => std_logic_vector(to_unsigned(36,8) ,
52453	 => std_logic_vector(to_unsigned(33,8) ,
52454	 => std_logic_vector(to_unsigned(28,8) ,
52455	 => std_logic_vector(to_unsigned(20,8) ,
52456	 => std_logic_vector(to_unsigned(18,8) ,
52457	 => std_logic_vector(to_unsigned(23,8) ,
52458	 => std_logic_vector(to_unsigned(17,8) ,
52459	 => std_logic_vector(to_unsigned(29,8) ,
52460	 => std_logic_vector(to_unsigned(36,8) ,
52461	 => std_logic_vector(to_unsigned(37,8) ,
52462	 => std_logic_vector(to_unsigned(32,8) ,
52463	 => std_logic_vector(to_unsigned(36,8) ,
52464	 => std_logic_vector(to_unsigned(29,8) ,
52465	 => std_logic_vector(to_unsigned(23,8) ,
52466	 => std_logic_vector(to_unsigned(16,8) ,
52467	 => std_logic_vector(to_unsigned(41,8) ,
52468	 => std_logic_vector(to_unsigned(32,8) ,
52469	 => std_logic_vector(to_unsigned(17,8) ,
52470	 => std_logic_vector(to_unsigned(8,8) ,
52471	 => std_logic_vector(to_unsigned(3,8) ,
52472	 => std_logic_vector(to_unsigned(8,8) ,
52473	 => std_logic_vector(to_unsigned(16,8) ,
52474	 => std_logic_vector(to_unsigned(12,8) ,
52475	 => std_logic_vector(to_unsigned(23,8) ,
52476	 => std_logic_vector(to_unsigned(22,8) ,
52477	 => std_logic_vector(to_unsigned(9,8) ,
52478	 => std_logic_vector(to_unsigned(27,8) ,
52479	 => std_logic_vector(to_unsigned(36,8) ,
52480	 => std_logic_vector(to_unsigned(30,8) ,
52481	 => std_logic_vector(to_unsigned(116,8) ,
52482	 => std_logic_vector(to_unsigned(130,8) ,
52483	 => std_logic_vector(to_unsigned(133,8) ,
52484	 => std_logic_vector(to_unsigned(127,8) ,
52485	 => std_logic_vector(to_unsigned(108,8) ,
52486	 => std_logic_vector(to_unsigned(107,8) ,
52487	 => std_logic_vector(to_unsigned(114,8) ,
52488	 => std_logic_vector(to_unsigned(112,8) ,
52489	 => std_logic_vector(to_unsigned(112,8) ,
52490	 => std_logic_vector(to_unsigned(109,8) ,
52491	 => std_logic_vector(to_unsigned(107,8) ,
52492	 => std_logic_vector(to_unsigned(116,8) ,
52493	 => std_logic_vector(to_unsigned(114,8) ,
52494	 => std_logic_vector(to_unsigned(116,8) ,
52495	 => std_logic_vector(to_unsigned(121,8) ,
52496	 => std_logic_vector(to_unsigned(124,8) ,
52497	 => std_logic_vector(to_unsigned(107,8) ,
52498	 => std_logic_vector(to_unsigned(97,8) ,
52499	 => std_logic_vector(to_unsigned(99,8) ,
52500	 => std_logic_vector(to_unsigned(108,8) ,
52501	 => std_logic_vector(to_unsigned(108,8) ,
52502	 => std_logic_vector(to_unsigned(93,8) ,
52503	 => std_logic_vector(to_unsigned(86,8) ,
52504	 => std_logic_vector(to_unsigned(51,8) ,
52505	 => std_logic_vector(to_unsigned(59,8) ,
52506	 => std_logic_vector(to_unsigned(65,8) ,
52507	 => std_logic_vector(to_unsigned(47,8) ,
52508	 => std_logic_vector(to_unsigned(45,8) ,
52509	 => std_logic_vector(to_unsigned(53,8) ,
52510	 => std_logic_vector(to_unsigned(51,8) ,
52511	 => std_logic_vector(to_unsigned(45,8) ,
52512	 => std_logic_vector(to_unsigned(64,8) ,
52513	 => std_logic_vector(to_unsigned(55,8) ,
52514	 => std_logic_vector(to_unsigned(36,8) ,
52515	 => std_logic_vector(to_unsigned(26,8) ,
52516	 => std_logic_vector(to_unsigned(28,8) ,
52517	 => std_logic_vector(to_unsigned(30,8) ,
52518	 => std_logic_vector(to_unsigned(33,8) ,
52519	 => std_logic_vector(to_unsigned(32,8) ,
52520	 => std_logic_vector(to_unsigned(38,8) ,
52521	 => std_logic_vector(to_unsigned(44,8) ,
52522	 => std_logic_vector(to_unsigned(46,8) ,
52523	 => std_logic_vector(to_unsigned(57,8) ,
52524	 => std_logic_vector(to_unsigned(48,8) ,
52525	 => std_logic_vector(to_unsigned(47,8) ,
52526	 => std_logic_vector(to_unsigned(56,8) ,
52527	 => std_logic_vector(to_unsigned(58,8) ,
52528	 => std_logic_vector(to_unsigned(76,8) ,
52529	 => std_logic_vector(to_unsigned(57,8) ,
52530	 => std_logic_vector(to_unsigned(56,8) ,
52531	 => std_logic_vector(to_unsigned(68,8) ,
52532	 => std_logic_vector(to_unsigned(63,8) ,
52533	 => std_logic_vector(to_unsigned(71,8) ,
52534	 => std_logic_vector(to_unsigned(73,8) ,
52535	 => std_logic_vector(to_unsigned(96,8) ,
52536	 => std_logic_vector(to_unsigned(95,8) ,
52537	 => std_logic_vector(to_unsigned(101,8) ,
52538	 => std_logic_vector(to_unsigned(91,8) ,
52539	 => std_logic_vector(to_unsigned(101,8) ,
52540	 => std_logic_vector(to_unsigned(90,8) ,
52541	 => std_logic_vector(to_unsigned(77,8) ,
52542	 => std_logic_vector(to_unsigned(105,8) ,
52543	 => std_logic_vector(to_unsigned(78,8) ,
52544	 => std_logic_vector(to_unsigned(60,8) ,
52545	 => std_logic_vector(to_unsigned(85,8) ,
52546	 => std_logic_vector(to_unsigned(77,8) ,
52547	 => std_logic_vector(to_unsigned(97,8) ,
52548	 => std_logic_vector(to_unsigned(101,8) ,
52549	 => std_logic_vector(to_unsigned(96,8) ,
52550	 => std_logic_vector(to_unsigned(121,8) ,
52551	 => std_logic_vector(to_unsigned(141,8) ,
52552	 => std_logic_vector(to_unsigned(80,8) ,
52553	 => std_logic_vector(to_unsigned(65,8) ,
52554	 => std_logic_vector(to_unsigned(104,8) ,
52555	 => std_logic_vector(to_unsigned(91,8) ,
52556	 => std_logic_vector(to_unsigned(86,8) ,
52557	 => std_logic_vector(to_unsigned(80,8) ,
52558	 => std_logic_vector(to_unsigned(82,8) ,
52559	 => std_logic_vector(to_unsigned(85,8) ,
52560	 => std_logic_vector(to_unsigned(58,8) ,
52561	 => std_logic_vector(to_unsigned(32,8) ,
52562	 => std_logic_vector(to_unsigned(34,8) ,
52563	 => std_logic_vector(to_unsigned(30,8) ,
52564	 => std_logic_vector(to_unsigned(30,8) ,
52565	 => std_logic_vector(to_unsigned(30,8) ,
52566	 => std_logic_vector(to_unsigned(40,8) ,
52567	 => std_logic_vector(to_unsigned(37,8) ,
52568	 => std_logic_vector(to_unsigned(33,8) ,
52569	 => std_logic_vector(to_unsigned(30,8) ,
52570	 => std_logic_vector(to_unsigned(30,8) ,
52571	 => std_logic_vector(to_unsigned(32,8) ,
52572	 => std_logic_vector(to_unsigned(37,8) ,
52573	 => std_logic_vector(to_unsigned(45,8) ,
52574	 => std_logic_vector(to_unsigned(45,8) ,
52575	 => std_logic_vector(to_unsigned(42,8) ,
52576	 => std_logic_vector(to_unsigned(43,8) ,
52577	 => std_logic_vector(to_unsigned(54,8) ,
52578	 => std_logic_vector(to_unsigned(51,8) ,
52579	 => std_logic_vector(to_unsigned(47,8) ,
52580	 => std_logic_vector(to_unsigned(40,8) ,
52581	 => std_logic_vector(to_unsigned(24,8) ,
52582	 => std_logic_vector(to_unsigned(24,8) ,
52583	 => std_logic_vector(to_unsigned(25,8) ,
52584	 => std_logic_vector(to_unsigned(49,8) ,
52585	 => std_logic_vector(to_unsigned(58,8) ,
52586	 => std_logic_vector(to_unsigned(45,8) ,
52587	 => std_logic_vector(to_unsigned(48,8) ,
52588	 => std_logic_vector(to_unsigned(45,8) ,
52589	 => std_logic_vector(to_unsigned(45,8) ,
52590	 => std_logic_vector(to_unsigned(45,8) ,
52591	 => std_logic_vector(to_unsigned(43,8) ,
52592	 => std_logic_vector(to_unsigned(46,8) ,
52593	 => std_logic_vector(to_unsigned(43,8) ,
52594	 => std_logic_vector(to_unsigned(40,8) ,
52595	 => std_logic_vector(to_unsigned(41,8) ,
52596	 => std_logic_vector(to_unsigned(37,8) ,
52597	 => std_logic_vector(to_unsigned(43,8) ,
52598	 => std_logic_vector(to_unsigned(28,8) ,
52599	 => std_logic_vector(to_unsigned(17,8) ,
52600	 => std_logic_vector(to_unsigned(18,8) ,
52601	 => std_logic_vector(to_unsigned(17,8) ,
52602	 => std_logic_vector(to_unsigned(17,8) ,
52603	 => std_logic_vector(to_unsigned(16,8) ,
52604	 => std_logic_vector(to_unsigned(57,8) ,
52605	 => std_logic_vector(to_unsigned(66,8) ,
52606	 => std_logic_vector(to_unsigned(46,8) ,
52607	 => std_logic_vector(to_unsigned(51,8) ,
52608	 => std_logic_vector(to_unsigned(38,8) ,
52609	 => std_logic_vector(to_unsigned(63,8) ,
52610	 => std_logic_vector(to_unsigned(41,8) ,
52611	 => std_logic_vector(to_unsigned(23,8) ,
52612	 => std_logic_vector(to_unsigned(32,8) ,
52613	 => std_logic_vector(to_unsigned(32,8) ,
52614	 => std_logic_vector(to_unsigned(34,8) ,
52615	 => std_logic_vector(to_unsigned(36,8) ,
52616	 => std_logic_vector(to_unsigned(35,8) ,
52617	 => std_logic_vector(to_unsigned(20,8) ,
52618	 => std_logic_vector(to_unsigned(12,8) ,
52619	 => std_logic_vector(to_unsigned(22,8) ,
52620	 => std_logic_vector(to_unsigned(18,8) ,
52621	 => std_logic_vector(to_unsigned(26,8) ,
52622	 => std_logic_vector(to_unsigned(66,8) ,
52623	 => std_logic_vector(to_unsigned(18,8) ,
52624	 => std_logic_vector(to_unsigned(32,8) ,
52625	 => std_logic_vector(to_unsigned(82,8) ,
52626	 => std_logic_vector(to_unsigned(44,8) ,
52627	 => std_logic_vector(to_unsigned(14,8) ,
52628	 => std_logic_vector(to_unsigned(6,8) ,
52629	 => std_logic_vector(to_unsigned(15,8) ,
52630	 => std_logic_vector(to_unsigned(58,8) ,
52631	 => std_logic_vector(to_unsigned(37,8) ,
52632	 => std_logic_vector(to_unsigned(44,8) ,
52633	 => std_logic_vector(to_unsigned(35,8) ,
52634	 => std_logic_vector(to_unsigned(48,8) ,
52635	 => std_logic_vector(to_unsigned(26,8) ,
52636	 => std_logic_vector(to_unsigned(62,8) ,
52637	 => std_logic_vector(to_unsigned(46,8) ,
52638	 => std_logic_vector(to_unsigned(9,8) ,
52639	 => std_logic_vector(to_unsigned(6,8) ,
52640	 => std_logic_vector(to_unsigned(7,8) ,
52641	 => std_logic_vector(to_unsigned(52,8) ,
52642	 => std_logic_vector(to_unsigned(59,8) ,
52643	 => std_logic_vector(to_unsigned(42,8) ,
52644	 => std_logic_vector(to_unsigned(43,8) ,
52645	 => std_logic_vector(to_unsigned(39,8) ,
52646	 => std_logic_vector(to_unsigned(44,8) ,
52647	 => std_logic_vector(to_unsigned(38,8) ,
52648	 => std_logic_vector(to_unsigned(41,8) ,
52649	 => std_logic_vector(to_unsigned(15,8) ,
52650	 => std_logic_vector(to_unsigned(5,8) ,
52651	 => std_logic_vector(to_unsigned(3,8) ,
52652	 => std_logic_vector(to_unsigned(8,8) ,
52653	 => std_logic_vector(to_unsigned(35,8) ,
52654	 => std_logic_vector(to_unsigned(13,8) ,
52655	 => std_logic_vector(to_unsigned(14,8) ,
52656	 => std_logic_vector(to_unsigned(27,8) ,
52657	 => std_logic_vector(to_unsigned(30,8) ,
52658	 => std_logic_vector(to_unsigned(29,8) ,
52659	 => std_logic_vector(to_unsigned(28,8) ,
52660	 => std_logic_vector(to_unsigned(26,8) ,
52661	 => std_logic_vector(to_unsigned(27,8) ,
52662	 => std_logic_vector(to_unsigned(25,8) ,
52663	 => std_logic_vector(to_unsigned(29,8) ,
52664	 => std_logic_vector(to_unsigned(26,8) ,
52665	 => std_logic_vector(to_unsigned(24,8) ,
52666	 => std_logic_vector(to_unsigned(32,8) ,
52667	 => std_logic_vector(to_unsigned(40,8) ,
52668	 => std_logic_vector(to_unsigned(28,8) ,
52669	 => std_logic_vector(to_unsigned(17,8) ,
52670	 => std_logic_vector(to_unsigned(31,8) ,
52671	 => std_logic_vector(to_unsigned(24,8) ,
52672	 => std_logic_vector(to_unsigned(27,8) ,
52673	 => std_logic_vector(to_unsigned(35,8) ,
52674	 => std_logic_vector(to_unsigned(34,8) ,
52675	 => std_logic_vector(to_unsigned(28,8) ,
52676	 => std_logic_vector(to_unsigned(26,8) ,
52677	 => std_logic_vector(to_unsigned(45,8) ,
52678	 => std_logic_vector(to_unsigned(68,8) ,
52679	 => std_logic_vector(to_unsigned(40,8) ,
52680	 => std_logic_vector(to_unsigned(19,8) ,
52681	 => std_logic_vector(to_unsigned(67,8) ,
52682	 => std_logic_vector(to_unsigned(80,8) ,
52683	 => std_logic_vector(to_unsigned(47,8) ,
52684	 => std_logic_vector(to_unsigned(12,8) ,
52685	 => std_logic_vector(to_unsigned(8,8) ,
52686	 => std_logic_vector(to_unsigned(6,8) ,
52687	 => std_logic_vector(to_unsigned(2,8) ,
52688	 => std_logic_vector(to_unsigned(6,8) ,
52689	 => std_logic_vector(to_unsigned(6,8) ,
52690	 => std_logic_vector(to_unsigned(10,8) ,
52691	 => std_logic_vector(to_unsigned(17,8) ,
52692	 => std_logic_vector(to_unsigned(13,8) ,
52693	 => std_logic_vector(to_unsigned(16,8) ,
52694	 => std_logic_vector(to_unsigned(18,8) ,
52695	 => std_logic_vector(to_unsigned(13,8) ,
52696	 => std_logic_vector(to_unsigned(14,8) ,
52697	 => std_logic_vector(to_unsigned(14,8) ,
52698	 => std_logic_vector(to_unsigned(14,8) ,
52699	 => std_logic_vector(to_unsigned(27,8) ,
52700	 => std_logic_vector(to_unsigned(22,8) ,
52701	 => std_logic_vector(to_unsigned(23,8) ,
52702	 => std_logic_vector(to_unsigned(33,8) ,
52703	 => std_logic_vector(to_unsigned(22,8) ,
52704	 => std_logic_vector(to_unsigned(23,8) ,
52705	 => std_logic_vector(to_unsigned(23,8) ,
52706	 => std_logic_vector(to_unsigned(17,8) ,
52707	 => std_logic_vector(to_unsigned(18,8) ,
52708	 => std_logic_vector(to_unsigned(23,8) ,
52709	 => std_logic_vector(to_unsigned(9,8) ,
52710	 => std_logic_vector(to_unsigned(16,8) ,
52711	 => std_logic_vector(to_unsigned(17,8) ,
52712	 => std_logic_vector(to_unsigned(27,8) ,
52713	 => std_logic_vector(to_unsigned(31,8) ,
52714	 => std_logic_vector(to_unsigned(23,8) ,
52715	 => std_logic_vector(to_unsigned(16,8) ,
52716	 => std_logic_vector(to_unsigned(11,8) ,
52717	 => std_logic_vector(to_unsigned(12,8) ,
52718	 => std_logic_vector(to_unsigned(15,8) ,
52719	 => std_logic_vector(to_unsigned(22,8) ,
52720	 => std_logic_vector(to_unsigned(20,8) ,
52721	 => std_logic_vector(to_unsigned(12,8) ,
52722	 => std_logic_vector(to_unsigned(28,8) ,
52723	 => std_logic_vector(to_unsigned(27,8) ,
52724	 => std_logic_vector(to_unsigned(15,8) ,
52725	 => std_logic_vector(to_unsigned(25,8) ,
52726	 => std_logic_vector(to_unsigned(26,8) ,
52727	 => std_logic_vector(to_unsigned(27,8) ,
52728	 => std_logic_vector(to_unsigned(45,8) ,
52729	 => std_logic_vector(to_unsigned(59,8) ,
52730	 => std_logic_vector(to_unsigned(47,8) ,
52731	 => std_logic_vector(to_unsigned(34,8) ,
52732	 => std_logic_vector(to_unsigned(53,8) ,
52733	 => std_logic_vector(to_unsigned(60,8) ,
52734	 => std_logic_vector(to_unsigned(45,8) ,
52735	 => std_logic_vector(to_unsigned(36,8) ,
52736	 => std_logic_vector(to_unsigned(16,8) ,
52737	 => std_logic_vector(to_unsigned(1,8) ,
52738	 => std_logic_vector(to_unsigned(0,8) ,
52739	 => std_logic_vector(to_unsigned(5,8) ,
52740	 => std_logic_vector(to_unsigned(42,8) ,
52741	 => std_logic_vector(to_unsigned(35,8) ,
52742	 => std_logic_vector(to_unsigned(35,8) ,
52743	 => std_logic_vector(to_unsigned(41,8) ,
52744	 => std_logic_vector(to_unsigned(35,8) ,
52745	 => std_logic_vector(to_unsigned(37,8) ,
52746	 => std_logic_vector(to_unsigned(19,8) ,
52747	 => std_logic_vector(to_unsigned(10,8) ,
52748	 => std_logic_vector(to_unsigned(14,8) ,
52749	 => std_logic_vector(to_unsigned(13,8) ,
52750	 => std_logic_vector(to_unsigned(13,8) ,
52751	 => std_logic_vector(to_unsigned(13,8) ,
52752	 => std_logic_vector(to_unsigned(10,8) ,
52753	 => std_logic_vector(to_unsigned(13,8) ,
52754	 => std_logic_vector(to_unsigned(10,8) ,
52755	 => std_logic_vector(to_unsigned(8,8) ,
52756	 => std_logic_vector(to_unsigned(9,8) ,
52757	 => std_logic_vector(to_unsigned(8,8) ,
52758	 => std_logic_vector(to_unsigned(3,8) ,
52759	 => std_logic_vector(to_unsigned(0,8) ,
52760	 => std_logic_vector(to_unsigned(0,8) ,
52761	 => std_logic_vector(to_unsigned(0,8) ,
52762	 => std_logic_vector(to_unsigned(0,8) ,
52763	 => std_logic_vector(to_unsigned(5,8) ,
52764	 => std_logic_vector(to_unsigned(17,8) ,
52765	 => std_logic_vector(to_unsigned(17,8) ,
52766	 => std_logic_vector(to_unsigned(14,8) ,
52767	 => std_logic_vector(to_unsigned(11,8) ,
52768	 => std_logic_vector(to_unsigned(12,8) ,
52769	 => std_logic_vector(to_unsigned(9,8) ,
52770	 => std_logic_vector(to_unsigned(13,8) ,
52771	 => std_logic_vector(to_unsigned(25,8) ,
52772	 => std_logic_vector(to_unsigned(30,8) ,
52773	 => std_logic_vector(to_unsigned(29,8) ,
52774	 => std_logic_vector(to_unsigned(19,8) ,
52775	 => std_logic_vector(to_unsigned(6,8) ,
52776	 => std_logic_vector(to_unsigned(6,8) ,
52777	 => std_logic_vector(to_unsigned(11,8) ,
52778	 => std_logic_vector(to_unsigned(13,8) ,
52779	 => std_logic_vector(to_unsigned(17,8) ,
52780	 => std_logic_vector(to_unsigned(17,8) ,
52781	 => std_logic_vector(to_unsigned(16,8) ,
52782	 => std_logic_vector(to_unsigned(20,8) ,
52783	 => std_logic_vector(to_unsigned(17,8) ,
52784	 => std_logic_vector(to_unsigned(22,8) ,
52785	 => std_logic_vector(to_unsigned(23,8) ,
52786	 => std_logic_vector(to_unsigned(23,8) ,
52787	 => std_logic_vector(to_unsigned(36,8) ,
52788	 => std_logic_vector(to_unsigned(35,8) ,
52789	 => std_logic_vector(to_unsigned(32,8) ,
52790	 => std_logic_vector(to_unsigned(29,8) ,
52791	 => std_logic_vector(to_unsigned(23,8) ,
52792	 => std_logic_vector(to_unsigned(32,8) ,
52793	 => std_logic_vector(to_unsigned(35,8) ,
52794	 => std_logic_vector(to_unsigned(31,8) ,
52795	 => std_logic_vector(to_unsigned(39,8) ,
52796	 => std_logic_vector(to_unsigned(23,8) ,
52797	 => std_logic_vector(to_unsigned(3,8) ,
52798	 => std_logic_vector(to_unsigned(13,8) ,
52799	 => std_logic_vector(to_unsigned(19,8) ,
52800	 => std_logic_vector(to_unsigned(9,8) ,
52801	 => std_logic_vector(to_unsigned(118,8) ,
52802	 => std_logic_vector(to_unsigned(116,8) ,
52803	 => std_logic_vector(to_unsigned(114,8) ,
52804	 => std_logic_vector(to_unsigned(118,8) ,
52805	 => std_logic_vector(to_unsigned(122,8) ,
52806	 => std_logic_vector(to_unsigned(127,8) ,
52807	 => std_logic_vector(to_unsigned(116,8) ,
52808	 => std_logic_vector(to_unsigned(115,8) ,
52809	 => std_logic_vector(to_unsigned(122,8) ,
52810	 => std_logic_vector(to_unsigned(124,8) ,
52811	 => std_logic_vector(to_unsigned(118,8) ,
52812	 => std_logic_vector(to_unsigned(111,8) ,
52813	 => std_logic_vector(to_unsigned(103,8) ,
52814	 => std_logic_vector(to_unsigned(96,8) ,
52815	 => std_logic_vector(to_unsigned(108,8) ,
52816	 => std_logic_vector(to_unsigned(109,8) ,
52817	 => std_logic_vector(to_unsigned(105,8) ,
52818	 => std_logic_vector(to_unsigned(108,8) ,
52819	 => std_logic_vector(to_unsigned(109,8) ,
52820	 => std_logic_vector(to_unsigned(114,8) ,
52821	 => std_logic_vector(to_unsigned(121,8) ,
52822	 => std_logic_vector(to_unsigned(95,8) ,
52823	 => std_logic_vector(to_unsigned(74,8) ,
52824	 => std_logic_vector(to_unsigned(56,8) ,
52825	 => std_logic_vector(to_unsigned(51,8) ,
52826	 => std_logic_vector(to_unsigned(48,8) ,
52827	 => std_logic_vector(to_unsigned(39,8) ,
52828	 => std_logic_vector(to_unsigned(41,8) ,
52829	 => std_logic_vector(to_unsigned(41,8) ,
52830	 => std_logic_vector(to_unsigned(64,8) ,
52831	 => std_logic_vector(to_unsigned(97,8) ,
52832	 => std_logic_vector(to_unsigned(87,8) ,
52833	 => std_logic_vector(to_unsigned(61,8) ,
52834	 => std_logic_vector(to_unsigned(44,8) ,
52835	 => std_logic_vector(to_unsigned(21,8) ,
52836	 => std_logic_vector(to_unsigned(27,8) ,
52837	 => std_logic_vector(to_unsigned(24,8) ,
52838	 => std_logic_vector(to_unsigned(25,8) ,
52839	 => std_logic_vector(to_unsigned(32,8) ,
52840	 => std_logic_vector(to_unsigned(43,8) ,
52841	 => std_logic_vector(to_unsigned(46,8) ,
52842	 => std_logic_vector(to_unsigned(45,8) ,
52843	 => std_logic_vector(to_unsigned(54,8) ,
52844	 => std_logic_vector(to_unsigned(61,8) ,
52845	 => std_logic_vector(to_unsigned(55,8) ,
52846	 => std_logic_vector(to_unsigned(54,8) ,
52847	 => std_logic_vector(to_unsigned(62,8) ,
52848	 => std_logic_vector(to_unsigned(52,8) ,
52849	 => std_logic_vector(to_unsigned(51,8) ,
52850	 => std_logic_vector(to_unsigned(67,8) ,
52851	 => std_logic_vector(to_unsigned(67,8) ,
52852	 => std_logic_vector(to_unsigned(72,8) ,
52853	 => std_logic_vector(to_unsigned(70,8) ,
52854	 => std_logic_vector(to_unsigned(60,8) ,
52855	 => std_logic_vector(to_unsigned(88,8) ,
52856	 => std_logic_vector(to_unsigned(79,8) ,
52857	 => std_logic_vector(to_unsigned(73,8) ,
52858	 => std_logic_vector(to_unsigned(82,8) ,
52859	 => std_logic_vector(to_unsigned(95,8) ,
52860	 => std_logic_vector(to_unsigned(92,8) ,
52861	 => std_logic_vector(to_unsigned(80,8) ,
52862	 => std_logic_vector(to_unsigned(99,8) ,
52863	 => std_logic_vector(to_unsigned(86,8) ,
52864	 => std_logic_vector(to_unsigned(56,8) ,
52865	 => std_logic_vector(to_unsigned(64,8) ,
52866	 => std_logic_vector(to_unsigned(72,8) ,
52867	 => std_logic_vector(to_unsigned(88,8) ,
52868	 => std_logic_vector(to_unsigned(91,8) ,
52869	 => std_logic_vector(to_unsigned(96,8) ,
52870	 => std_logic_vector(to_unsigned(118,8) ,
52871	 => std_logic_vector(to_unsigned(142,8) ,
52872	 => std_logic_vector(to_unsigned(77,8) ,
52873	 => std_logic_vector(to_unsigned(57,8) ,
52874	 => std_logic_vector(to_unsigned(99,8) ,
52875	 => std_logic_vector(to_unsigned(91,8) ,
52876	 => std_logic_vector(to_unsigned(87,8) ,
52877	 => std_logic_vector(to_unsigned(87,8) ,
52878	 => std_logic_vector(to_unsigned(87,8) ,
52879	 => std_logic_vector(to_unsigned(97,8) ,
52880	 => std_logic_vector(to_unsigned(61,8) ,
52881	 => std_logic_vector(to_unsigned(25,8) ,
52882	 => std_logic_vector(to_unsigned(27,8) ,
52883	 => std_logic_vector(to_unsigned(27,8) ,
52884	 => std_logic_vector(to_unsigned(32,8) ,
52885	 => std_logic_vector(to_unsigned(43,8) ,
52886	 => std_logic_vector(to_unsigned(45,8) ,
52887	 => std_logic_vector(to_unsigned(25,8) ,
52888	 => std_logic_vector(to_unsigned(32,8) ,
52889	 => std_logic_vector(to_unsigned(40,8) ,
52890	 => std_logic_vector(to_unsigned(37,8) ,
52891	 => std_logic_vector(to_unsigned(44,8) ,
52892	 => std_logic_vector(to_unsigned(54,8) ,
52893	 => std_logic_vector(to_unsigned(53,8) ,
52894	 => std_logic_vector(to_unsigned(53,8) ,
52895	 => std_logic_vector(to_unsigned(55,8) ,
52896	 => std_logic_vector(to_unsigned(65,8) ,
52897	 => std_logic_vector(to_unsigned(70,8) ,
52898	 => std_logic_vector(to_unsigned(73,8) ,
52899	 => std_logic_vector(to_unsigned(87,8) ,
52900	 => std_logic_vector(to_unsigned(90,8) ,
52901	 => std_logic_vector(to_unsigned(67,8) ,
52902	 => std_logic_vector(to_unsigned(42,8) ,
52903	 => std_logic_vector(to_unsigned(22,8) ,
52904	 => std_logic_vector(to_unsigned(33,8) ,
52905	 => std_logic_vector(to_unsigned(52,8) ,
52906	 => std_logic_vector(to_unsigned(41,8) ,
52907	 => std_logic_vector(to_unsigned(43,8) ,
52908	 => std_logic_vector(to_unsigned(44,8) ,
52909	 => std_logic_vector(to_unsigned(42,8) ,
52910	 => std_logic_vector(to_unsigned(40,8) ,
52911	 => std_logic_vector(to_unsigned(41,8) ,
52912	 => std_logic_vector(to_unsigned(43,8) ,
52913	 => std_logic_vector(to_unsigned(43,8) ,
52914	 => std_logic_vector(to_unsigned(40,8) ,
52915	 => std_logic_vector(to_unsigned(42,8) ,
52916	 => std_logic_vector(to_unsigned(39,8) ,
52917	 => std_logic_vector(to_unsigned(42,8) ,
52918	 => std_logic_vector(to_unsigned(36,8) ,
52919	 => std_logic_vector(to_unsigned(19,8) ,
52920	 => std_logic_vector(to_unsigned(15,8) ,
52921	 => std_logic_vector(to_unsigned(23,8) ,
52922	 => std_logic_vector(to_unsigned(23,8) ,
52923	 => std_logic_vector(to_unsigned(18,8) ,
52924	 => std_logic_vector(to_unsigned(54,8) ,
52925	 => std_logic_vector(to_unsigned(68,8) ,
52926	 => std_logic_vector(to_unsigned(48,8) ,
52927	 => std_logic_vector(to_unsigned(45,8) ,
52928	 => std_logic_vector(to_unsigned(42,8) ,
52929	 => std_logic_vector(to_unsigned(65,8) ,
52930	 => std_logic_vector(to_unsigned(50,8) ,
52931	 => std_logic_vector(to_unsigned(32,8) ,
52932	 => std_logic_vector(to_unsigned(44,8) ,
52933	 => std_logic_vector(to_unsigned(39,8) ,
52934	 => std_logic_vector(to_unsigned(28,8) ,
52935	 => std_logic_vector(to_unsigned(21,8) ,
52936	 => std_logic_vector(to_unsigned(26,8) ,
52937	 => std_logic_vector(to_unsigned(31,8) ,
52938	 => std_logic_vector(to_unsigned(24,8) ,
52939	 => std_logic_vector(to_unsigned(16,8) ,
52940	 => std_logic_vector(to_unsigned(9,8) ,
52941	 => std_logic_vector(to_unsigned(20,8) ,
52942	 => std_logic_vector(to_unsigned(68,8) ,
52943	 => std_logic_vector(to_unsigned(25,8) ,
52944	 => std_logic_vector(to_unsigned(33,8) ,
52945	 => std_logic_vector(to_unsigned(78,8) ,
52946	 => std_logic_vector(to_unsigned(46,8) ,
52947	 => std_logic_vector(to_unsigned(13,8) ,
52948	 => std_logic_vector(to_unsigned(4,8) ,
52949	 => std_logic_vector(to_unsigned(13,8) ,
52950	 => std_logic_vector(to_unsigned(62,8) ,
52951	 => std_logic_vector(to_unsigned(41,8) ,
52952	 => std_logic_vector(to_unsigned(52,8) ,
52953	 => std_logic_vector(to_unsigned(63,8) ,
52954	 => std_logic_vector(to_unsigned(61,8) ,
52955	 => std_logic_vector(to_unsigned(38,8) ,
52956	 => std_logic_vector(to_unsigned(74,8) ,
52957	 => std_logic_vector(to_unsigned(51,8) ,
52958	 => std_logic_vector(to_unsigned(12,8) ,
52959	 => std_logic_vector(to_unsigned(6,8) ,
52960	 => std_logic_vector(to_unsigned(6,8) ,
52961	 => std_logic_vector(to_unsigned(49,8) ,
52962	 => std_logic_vector(to_unsigned(37,8) ,
52963	 => std_logic_vector(to_unsigned(28,8) ,
52964	 => std_logic_vector(to_unsigned(40,8) ,
52965	 => std_logic_vector(to_unsigned(35,8) ,
52966	 => std_logic_vector(to_unsigned(33,8) ,
52967	 => std_logic_vector(to_unsigned(34,8) ,
52968	 => std_logic_vector(to_unsigned(44,8) ,
52969	 => std_logic_vector(to_unsigned(17,8) ,
52970	 => std_logic_vector(to_unsigned(8,8) ,
52971	 => std_logic_vector(to_unsigned(3,8) ,
52972	 => std_logic_vector(to_unsigned(9,8) ,
52973	 => std_logic_vector(to_unsigned(68,8) ,
52974	 => std_logic_vector(to_unsigned(30,8) ,
52975	 => std_logic_vector(to_unsigned(25,8) ,
52976	 => std_logic_vector(to_unsigned(23,8) ,
52977	 => std_logic_vector(to_unsigned(19,8) ,
52978	 => std_logic_vector(to_unsigned(20,8) ,
52979	 => std_logic_vector(to_unsigned(21,8) ,
52980	 => std_logic_vector(to_unsigned(20,8) ,
52981	 => std_logic_vector(to_unsigned(17,8) ,
52982	 => std_logic_vector(to_unsigned(23,8) ,
52983	 => std_logic_vector(to_unsigned(28,8) ,
52984	 => std_logic_vector(to_unsigned(20,8) ,
52985	 => std_logic_vector(to_unsigned(29,8) ,
52986	 => std_logic_vector(to_unsigned(32,8) ,
52987	 => std_logic_vector(to_unsigned(35,8) ,
52988	 => std_logic_vector(to_unsigned(24,8) ,
52989	 => std_logic_vector(to_unsigned(17,8) ,
52990	 => std_logic_vector(to_unsigned(22,8) ,
52991	 => std_logic_vector(to_unsigned(15,8) ,
52992	 => std_logic_vector(to_unsigned(29,8) ,
52993	 => std_logic_vector(to_unsigned(33,8) ,
52994	 => std_logic_vector(to_unsigned(41,8) ,
52995	 => std_logic_vector(to_unsigned(32,8) ,
52996	 => std_logic_vector(to_unsigned(20,8) ,
52997	 => std_logic_vector(to_unsigned(27,8) ,
52998	 => std_logic_vector(to_unsigned(25,8) ,
52999	 => std_logic_vector(to_unsigned(22,8) ,
53000	 => std_logic_vector(to_unsigned(23,8) ,
53001	 => std_logic_vector(to_unsigned(34,8) ,
53002	 => std_logic_vector(to_unsigned(39,8) ,
53003	 => std_logic_vector(to_unsigned(35,8) ,
53004	 => std_logic_vector(to_unsigned(17,8) ,
53005	 => std_logic_vector(to_unsigned(10,8) ,
53006	 => std_logic_vector(to_unsigned(6,8) ,
53007	 => std_logic_vector(to_unsigned(16,8) ,
53008	 => std_logic_vector(to_unsigned(25,8) ,
53009	 => std_logic_vector(to_unsigned(5,8) ,
53010	 => std_logic_vector(to_unsigned(11,8) ,
53011	 => std_logic_vector(to_unsigned(18,8) ,
53012	 => std_logic_vector(to_unsigned(18,8) ,
53013	 => std_logic_vector(to_unsigned(19,8) ,
53014	 => std_logic_vector(to_unsigned(13,8) ,
53015	 => std_logic_vector(to_unsigned(13,8) ,
53016	 => std_logic_vector(to_unsigned(13,8) ,
53017	 => std_logic_vector(to_unsigned(11,8) ,
53018	 => std_logic_vector(to_unsigned(17,8) ,
53019	 => std_logic_vector(to_unsigned(24,8) ,
53020	 => std_logic_vector(to_unsigned(16,8) ,
53021	 => std_logic_vector(to_unsigned(17,8) ,
53022	 => std_logic_vector(to_unsigned(32,8) ,
53023	 => std_logic_vector(to_unsigned(28,8) ,
53024	 => std_logic_vector(to_unsigned(15,8) ,
53025	 => std_logic_vector(to_unsigned(12,8) ,
53026	 => std_logic_vector(to_unsigned(10,8) ,
53027	 => std_logic_vector(to_unsigned(11,8) ,
53028	 => std_logic_vector(to_unsigned(14,8) ,
53029	 => std_logic_vector(to_unsigned(8,8) ,
53030	 => std_logic_vector(to_unsigned(11,8) ,
53031	 => std_logic_vector(to_unsigned(23,8) ,
53032	 => std_logic_vector(to_unsigned(32,8) ,
53033	 => std_logic_vector(to_unsigned(33,8) ,
53034	 => std_logic_vector(to_unsigned(24,8) ,
53035	 => std_logic_vector(to_unsigned(16,8) ,
53036	 => std_logic_vector(to_unsigned(8,8) ,
53037	 => std_logic_vector(to_unsigned(12,8) ,
53038	 => std_logic_vector(to_unsigned(12,8) ,
53039	 => std_logic_vector(to_unsigned(14,8) ,
53040	 => std_logic_vector(to_unsigned(12,8) ,
53041	 => std_logic_vector(to_unsigned(17,8) ,
53042	 => std_logic_vector(to_unsigned(35,8) ,
53043	 => std_logic_vector(to_unsigned(23,8) ,
53044	 => std_logic_vector(to_unsigned(18,8) ,
53045	 => std_logic_vector(to_unsigned(18,8) ,
53046	 => std_logic_vector(to_unsigned(17,8) ,
53047	 => std_logic_vector(to_unsigned(20,8) ,
53048	 => std_logic_vector(to_unsigned(49,8) ,
53049	 => std_logic_vector(to_unsigned(64,8) ,
53050	 => std_logic_vector(to_unsigned(51,8) ,
53051	 => std_logic_vector(to_unsigned(28,8) ,
53052	 => std_logic_vector(to_unsigned(25,8) ,
53053	 => std_logic_vector(to_unsigned(33,8) ,
53054	 => std_logic_vector(to_unsigned(27,8) ,
53055	 => std_logic_vector(to_unsigned(21,8) ,
53056	 => std_logic_vector(to_unsigned(28,8) ,
53057	 => std_logic_vector(to_unsigned(8,8) ,
53058	 => std_logic_vector(to_unsigned(0,8) ,
53059	 => std_logic_vector(to_unsigned(1,8) ,
53060	 => std_logic_vector(to_unsigned(13,8) ,
53061	 => std_logic_vector(to_unsigned(25,8) ,
53062	 => std_logic_vector(to_unsigned(18,8) ,
53063	 => std_logic_vector(to_unsigned(24,8) ,
53064	 => std_logic_vector(to_unsigned(27,8) ,
53065	 => std_logic_vector(to_unsigned(22,8) ,
53066	 => std_logic_vector(to_unsigned(19,8) ,
53067	 => std_logic_vector(to_unsigned(15,8) ,
53068	 => std_logic_vector(to_unsigned(12,8) ,
53069	 => std_logic_vector(to_unsigned(14,8) ,
53070	 => std_logic_vector(to_unsigned(12,8) ,
53071	 => std_logic_vector(to_unsigned(11,8) ,
53072	 => std_logic_vector(to_unsigned(11,8) ,
53073	 => std_logic_vector(to_unsigned(11,8) ,
53074	 => std_logic_vector(to_unsigned(9,8) ,
53075	 => std_logic_vector(to_unsigned(12,8) ,
53076	 => std_logic_vector(to_unsigned(10,8) ,
53077	 => std_logic_vector(to_unsigned(8,8) ,
53078	 => std_logic_vector(to_unsigned(5,8) ,
53079	 => std_logic_vector(to_unsigned(1,8) ,
53080	 => std_logic_vector(to_unsigned(0,8) ,
53081	 => std_logic_vector(to_unsigned(0,8) ,
53082	 => std_logic_vector(to_unsigned(0,8) ,
53083	 => std_logic_vector(to_unsigned(2,8) ,
53084	 => std_logic_vector(to_unsigned(9,8) ,
53085	 => std_logic_vector(to_unsigned(10,8) ,
53086	 => std_logic_vector(to_unsigned(11,8) ,
53087	 => std_logic_vector(to_unsigned(13,8) ,
53088	 => std_logic_vector(to_unsigned(17,8) ,
53089	 => std_logic_vector(to_unsigned(10,8) ,
53090	 => std_logic_vector(to_unsigned(19,8) ,
53091	 => std_logic_vector(to_unsigned(17,8) ,
53092	 => std_logic_vector(to_unsigned(23,8) ,
53093	 => std_logic_vector(to_unsigned(22,8) ,
53094	 => std_logic_vector(to_unsigned(17,8) ,
53095	 => std_logic_vector(to_unsigned(14,8) ,
53096	 => std_logic_vector(to_unsigned(11,8) ,
53097	 => std_logic_vector(to_unsigned(6,8) ,
53098	 => std_logic_vector(to_unsigned(5,8) ,
53099	 => std_logic_vector(to_unsigned(13,8) ,
53100	 => std_logic_vector(to_unsigned(17,8) ,
53101	 => std_logic_vector(to_unsigned(14,8) ,
53102	 => std_logic_vector(to_unsigned(11,8) ,
53103	 => std_logic_vector(to_unsigned(2,8) ,
53104	 => std_logic_vector(to_unsigned(6,8) ,
53105	 => std_logic_vector(to_unsigned(15,8) ,
53106	 => std_logic_vector(to_unsigned(9,8) ,
53107	 => std_logic_vector(to_unsigned(39,8) ,
53108	 => std_logic_vector(to_unsigned(21,8) ,
53109	 => std_logic_vector(to_unsigned(12,8) ,
53110	 => std_logic_vector(to_unsigned(6,8) ,
53111	 => std_logic_vector(to_unsigned(3,8) ,
53112	 => std_logic_vector(to_unsigned(15,8) ,
53113	 => std_logic_vector(to_unsigned(20,8) ,
53114	 => std_logic_vector(to_unsigned(32,8) ,
53115	 => std_logic_vector(to_unsigned(49,8) ,
53116	 => std_logic_vector(to_unsigned(41,8) ,
53117	 => std_logic_vector(to_unsigned(35,8) ,
53118	 => std_logic_vector(to_unsigned(54,8) ,
53119	 => std_logic_vector(to_unsigned(72,8) ,
53120	 => std_logic_vector(to_unsigned(61,8) ,
53121	 => std_logic_vector(to_unsigned(118,8) ,
53122	 => std_logic_vector(to_unsigned(118,8) ,
53123	 => std_logic_vector(to_unsigned(121,8) ,
53124	 => std_logic_vector(to_unsigned(124,8) ,
53125	 => std_logic_vector(to_unsigned(130,8) ,
53126	 => std_logic_vector(to_unsigned(116,8) ,
53127	 => std_logic_vector(to_unsigned(112,8) ,
53128	 => std_logic_vector(to_unsigned(127,8) ,
53129	 => std_logic_vector(to_unsigned(133,8) ,
53130	 => std_logic_vector(to_unsigned(124,8) ,
53131	 => std_logic_vector(to_unsigned(118,8) ,
53132	 => std_logic_vector(to_unsigned(107,8) ,
53133	 => std_logic_vector(to_unsigned(101,8) ,
53134	 => std_logic_vector(to_unsigned(101,8) ,
53135	 => std_logic_vector(to_unsigned(109,8) ,
53136	 => std_logic_vector(to_unsigned(115,8) ,
53137	 => std_logic_vector(to_unsigned(114,8) ,
53138	 => std_logic_vector(to_unsigned(119,8) ,
53139	 => std_logic_vector(to_unsigned(92,8) ,
53140	 => std_logic_vector(to_unsigned(82,8) ,
53141	 => std_logic_vector(to_unsigned(96,8) ,
53142	 => std_logic_vector(to_unsigned(63,8) ,
53143	 => std_logic_vector(to_unsigned(48,8) ,
53144	 => std_logic_vector(to_unsigned(48,8) ,
53145	 => std_logic_vector(to_unsigned(37,8) ,
53146	 => std_logic_vector(to_unsigned(37,8) ,
53147	 => std_logic_vector(to_unsigned(48,8) ,
53148	 => std_logic_vector(to_unsigned(76,8) ,
53149	 => std_logic_vector(to_unsigned(78,8) ,
53150	 => std_logic_vector(to_unsigned(81,8) ,
53151	 => std_logic_vector(to_unsigned(86,8) ,
53152	 => std_logic_vector(to_unsigned(64,8) ,
53153	 => std_logic_vector(to_unsigned(44,8) ,
53154	 => std_logic_vector(to_unsigned(41,8) ,
53155	 => std_logic_vector(to_unsigned(28,8) ,
53156	 => std_logic_vector(to_unsigned(28,8) ,
53157	 => std_logic_vector(to_unsigned(29,8) ,
53158	 => std_logic_vector(to_unsigned(35,8) ,
53159	 => std_logic_vector(to_unsigned(35,8) ,
53160	 => std_logic_vector(to_unsigned(43,8) ,
53161	 => std_logic_vector(to_unsigned(40,8) ,
53162	 => std_logic_vector(to_unsigned(35,8) ,
53163	 => std_logic_vector(to_unsigned(42,8) ,
53164	 => std_logic_vector(to_unsigned(45,8) ,
53165	 => std_logic_vector(to_unsigned(45,8) ,
53166	 => std_logic_vector(to_unsigned(45,8) ,
53167	 => std_logic_vector(to_unsigned(50,8) ,
53168	 => std_logic_vector(to_unsigned(52,8) ,
53169	 => std_logic_vector(to_unsigned(69,8) ,
53170	 => std_logic_vector(to_unsigned(91,8) ,
53171	 => std_logic_vector(to_unsigned(93,8) ,
53172	 => std_logic_vector(to_unsigned(108,8) ,
53173	 => std_logic_vector(to_unsigned(112,8) ,
53174	 => std_logic_vector(to_unsigned(90,8) ,
53175	 => std_logic_vector(to_unsigned(82,8) ,
53176	 => std_logic_vector(to_unsigned(64,8) ,
53177	 => std_logic_vector(to_unsigned(61,8) ,
53178	 => std_logic_vector(to_unsigned(71,8) ,
53179	 => std_logic_vector(to_unsigned(80,8) ,
53180	 => std_logic_vector(to_unsigned(81,8) ,
53181	 => std_logic_vector(to_unsigned(77,8) ,
53182	 => std_logic_vector(to_unsigned(91,8) ,
53183	 => std_logic_vector(to_unsigned(73,8) ,
53184	 => std_logic_vector(to_unsigned(58,8) ,
53185	 => std_logic_vector(to_unsigned(71,8) ,
53186	 => std_logic_vector(to_unsigned(82,8) ,
53187	 => std_logic_vector(to_unsigned(88,8) ,
53188	 => std_logic_vector(to_unsigned(87,8) ,
53189	 => std_logic_vector(to_unsigned(84,8) ,
53190	 => std_logic_vector(to_unsigned(115,8) ,
53191	 => std_logic_vector(to_unsigned(131,8) ,
53192	 => std_logic_vector(to_unsigned(95,8) ,
53193	 => std_logic_vector(to_unsigned(74,8) ,
53194	 => std_logic_vector(to_unsigned(93,8) ,
53195	 => std_logic_vector(to_unsigned(91,8) ,
53196	 => std_logic_vector(to_unsigned(88,8) ,
53197	 => std_logic_vector(to_unsigned(85,8) ,
53198	 => std_logic_vector(to_unsigned(90,8) ,
53199	 => std_logic_vector(to_unsigned(95,8) ,
53200	 => std_logic_vector(to_unsigned(65,8) ,
53201	 => std_logic_vector(to_unsigned(17,8) ,
53202	 => std_logic_vector(to_unsigned(23,8) ,
53203	 => std_logic_vector(to_unsigned(24,8) ,
53204	 => std_logic_vector(to_unsigned(23,8) ,
53205	 => std_logic_vector(to_unsigned(34,8) ,
53206	 => std_logic_vector(to_unsigned(45,8) ,
53207	 => std_logic_vector(to_unsigned(41,8) ,
53208	 => std_logic_vector(to_unsigned(93,8) ,
53209	 => std_logic_vector(to_unsigned(97,8) ,
53210	 => std_logic_vector(to_unsigned(45,8) ,
53211	 => std_logic_vector(to_unsigned(51,8) ,
53212	 => std_logic_vector(to_unsigned(58,8) ,
53213	 => std_logic_vector(to_unsigned(61,8) ,
53214	 => std_logic_vector(to_unsigned(80,8) ,
53215	 => std_logic_vector(to_unsigned(107,8) ,
53216	 => std_logic_vector(to_unsigned(119,8) ,
53217	 => std_logic_vector(to_unsigned(118,8) ,
53218	 => std_logic_vector(to_unsigned(119,8) ,
53219	 => std_logic_vector(to_unsigned(124,8) ,
53220	 => std_logic_vector(to_unsigned(128,8) ,
53221	 => std_logic_vector(to_unsigned(139,8) ,
53222	 => std_logic_vector(to_unsigned(99,8) ,
53223	 => std_logic_vector(to_unsigned(58,8) ,
53224	 => std_logic_vector(to_unsigned(54,8) ,
53225	 => std_logic_vector(to_unsigned(51,8) ,
53226	 => std_logic_vector(to_unsigned(40,8) ,
53227	 => std_logic_vector(to_unsigned(41,8) ,
53228	 => std_logic_vector(to_unsigned(37,8) ,
53229	 => std_logic_vector(to_unsigned(37,8) ,
53230	 => std_logic_vector(to_unsigned(37,8) ,
53231	 => std_logic_vector(to_unsigned(38,8) ,
53232	 => std_logic_vector(to_unsigned(35,8) ,
53233	 => std_logic_vector(to_unsigned(37,8) ,
53234	 => std_logic_vector(to_unsigned(37,8) ,
53235	 => std_logic_vector(to_unsigned(39,8) ,
53236	 => std_logic_vector(to_unsigned(43,8) ,
53237	 => std_logic_vector(to_unsigned(39,8) ,
53238	 => std_logic_vector(to_unsigned(33,8) ,
53239	 => std_logic_vector(to_unsigned(19,8) ,
53240	 => std_logic_vector(to_unsigned(16,8) ,
53241	 => std_logic_vector(to_unsigned(20,8) ,
53242	 => std_logic_vector(to_unsigned(18,8) ,
53243	 => std_logic_vector(to_unsigned(20,8) ,
53244	 => std_logic_vector(to_unsigned(53,8) ,
53245	 => std_logic_vector(to_unsigned(67,8) ,
53246	 => std_logic_vector(to_unsigned(45,8) ,
53247	 => std_logic_vector(to_unsigned(38,8) ,
53248	 => std_logic_vector(to_unsigned(39,8) ,
53249	 => std_logic_vector(to_unsigned(57,8) ,
53250	 => std_logic_vector(to_unsigned(46,8) ,
53251	 => std_logic_vector(to_unsigned(36,8) ,
53252	 => std_logic_vector(to_unsigned(44,8) ,
53253	 => std_logic_vector(to_unsigned(29,8) ,
53254	 => std_logic_vector(to_unsigned(14,8) ,
53255	 => std_logic_vector(to_unsigned(17,8) ,
53256	 => std_logic_vector(to_unsigned(27,8) ,
53257	 => std_logic_vector(to_unsigned(29,8) ,
53258	 => std_logic_vector(to_unsigned(17,8) ,
53259	 => std_logic_vector(to_unsigned(12,8) ,
53260	 => std_logic_vector(to_unsigned(7,8) ,
53261	 => std_logic_vector(to_unsigned(17,8) ,
53262	 => std_logic_vector(to_unsigned(60,8) ,
53263	 => std_logic_vector(to_unsigned(32,8) ,
53264	 => std_logic_vector(to_unsigned(41,8) ,
53265	 => std_logic_vector(to_unsigned(71,8) ,
53266	 => std_logic_vector(to_unsigned(55,8) ,
53267	 => std_logic_vector(to_unsigned(32,8) ,
53268	 => std_logic_vector(to_unsigned(16,8) ,
53269	 => std_logic_vector(to_unsigned(27,8) ,
53270	 => std_logic_vector(to_unsigned(47,8) ,
53271	 => std_logic_vector(to_unsigned(13,8) ,
53272	 => std_logic_vector(to_unsigned(38,8) ,
53273	 => std_logic_vector(to_unsigned(49,8) ,
53274	 => std_logic_vector(to_unsigned(47,8) ,
53275	 => std_logic_vector(to_unsigned(37,8) ,
53276	 => std_logic_vector(to_unsigned(71,8) ,
53277	 => std_logic_vector(to_unsigned(48,8) ,
53278	 => std_logic_vector(to_unsigned(10,8) ,
53279	 => std_logic_vector(to_unsigned(9,8) ,
53280	 => std_logic_vector(to_unsigned(7,8) ,
53281	 => std_logic_vector(to_unsigned(38,8) ,
53282	 => std_logic_vector(to_unsigned(45,8) ,
53283	 => std_logic_vector(to_unsigned(37,8) ,
53284	 => std_logic_vector(to_unsigned(39,8) ,
53285	 => std_logic_vector(to_unsigned(33,8) ,
53286	 => std_logic_vector(to_unsigned(24,8) ,
53287	 => std_logic_vector(to_unsigned(19,8) ,
53288	 => std_logic_vector(to_unsigned(43,8) ,
53289	 => std_logic_vector(to_unsigned(16,8) ,
53290	 => std_logic_vector(to_unsigned(8,8) ,
53291	 => std_logic_vector(to_unsigned(4,8) ,
53292	 => std_logic_vector(to_unsigned(11,8) ,
53293	 => std_logic_vector(to_unsigned(61,8) ,
53294	 => std_logic_vector(to_unsigned(20,8) ,
53295	 => std_logic_vector(to_unsigned(12,8) ,
53296	 => std_logic_vector(to_unsigned(22,8) ,
53297	 => std_logic_vector(to_unsigned(19,8) ,
53298	 => std_logic_vector(to_unsigned(15,8) ,
53299	 => std_logic_vector(to_unsigned(15,8) ,
53300	 => std_logic_vector(to_unsigned(16,8) ,
53301	 => std_logic_vector(to_unsigned(17,8) ,
53302	 => std_logic_vector(to_unsigned(17,8) ,
53303	 => std_logic_vector(to_unsigned(23,8) ,
53304	 => std_logic_vector(to_unsigned(23,8) ,
53305	 => std_logic_vector(to_unsigned(31,8) ,
53306	 => std_logic_vector(to_unsigned(32,8) ,
53307	 => std_logic_vector(to_unsigned(40,8) ,
53308	 => std_logic_vector(to_unsigned(31,8) ,
53309	 => std_logic_vector(to_unsigned(15,8) ,
53310	 => std_logic_vector(to_unsigned(13,8) ,
53311	 => std_logic_vector(to_unsigned(20,8) ,
53312	 => std_logic_vector(to_unsigned(29,8) ,
53313	 => std_logic_vector(to_unsigned(31,8) ,
53314	 => std_logic_vector(to_unsigned(40,8) ,
53315	 => std_logic_vector(to_unsigned(29,8) ,
53316	 => std_logic_vector(to_unsigned(12,8) ,
53317	 => std_logic_vector(to_unsigned(10,8) ,
53318	 => std_logic_vector(to_unsigned(9,8) ,
53319	 => std_logic_vector(to_unsigned(13,8) ,
53320	 => std_logic_vector(to_unsigned(18,8) ,
53321	 => std_logic_vector(to_unsigned(17,8) ,
53322	 => std_logic_vector(to_unsigned(14,8) ,
53323	 => std_logic_vector(to_unsigned(20,8) ,
53324	 => std_logic_vector(to_unsigned(22,8) ,
53325	 => std_logic_vector(to_unsigned(15,8) ,
53326	 => std_logic_vector(to_unsigned(13,8) ,
53327	 => std_logic_vector(to_unsigned(24,8) ,
53328	 => std_logic_vector(to_unsigned(25,8) ,
53329	 => std_logic_vector(to_unsigned(7,8) ,
53330	 => std_logic_vector(to_unsigned(12,8) ,
53331	 => std_logic_vector(to_unsigned(19,8) ,
53332	 => std_logic_vector(to_unsigned(20,8) ,
53333	 => std_logic_vector(to_unsigned(19,8) ,
53334	 => std_logic_vector(to_unsigned(12,8) ,
53335	 => std_logic_vector(to_unsigned(23,8) ,
53336	 => std_logic_vector(to_unsigned(28,8) ,
53337	 => std_logic_vector(to_unsigned(18,8) ,
53338	 => std_logic_vector(to_unsigned(16,8) ,
53339	 => std_logic_vector(to_unsigned(17,8) ,
53340	 => std_logic_vector(to_unsigned(11,8) ,
53341	 => std_logic_vector(to_unsigned(13,8) ,
53342	 => std_logic_vector(to_unsigned(33,8) ,
53343	 => std_logic_vector(to_unsigned(37,8) ,
53344	 => std_logic_vector(to_unsigned(15,8) ,
53345	 => std_logic_vector(to_unsigned(10,8) ,
53346	 => std_logic_vector(to_unsigned(10,8) ,
53347	 => std_logic_vector(to_unsigned(10,8) ,
53348	 => std_logic_vector(to_unsigned(11,8) ,
53349	 => std_logic_vector(to_unsigned(10,8) ,
53350	 => std_logic_vector(to_unsigned(17,8) ,
53351	 => std_logic_vector(to_unsigned(30,8) ,
53352	 => std_logic_vector(to_unsigned(28,8) ,
53353	 => std_logic_vector(to_unsigned(32,8) ,
53354	 => std_logic_vector(to_unsigned(20,8) ,
53355	 => std_logic_vector(to_unsigned(11,8) ,
53356	 => std_logic_vector(to_unsigned(12,8) ,
53357	 => std_logic_vector(to_unsigned(13,8) ,
53358	 => std_logic_vector(to_unsigned(19,8) ,
53359	 => std_logic_vector(to_unsigned(16,8) ,
53360	 => std_logic_vector(to_unsigned(18,8) ,
53361	 => std_logic_vector(to_unsigned(31,8) ,
53362	 => std_logic_vector(to_unsigned(22,8) ,
53363	 => std_logic_vector(to_unsigned(22,8) ,
53364	 => std_logic_vector(to_unsigned(27,8) ,
53365	 => std_logic_vector(to_unsigned(25,8) ,
53366	 => std_logic_vector(to_unsigned(26,8) ,
53367	 => std_logic_vector(to_unsigned(29,8) ,
53368	 => std_logic_vector(to_unsigned(45,8) ,
53369	 => std_logic_vector(to_unsigned(32,8) ,
53370	 => std_logic_vector(to_unsigned(33,8) ,
53371	 => std_logic_vector(to_unsigned(30,8) ,
53372	 => std_logic_vector(to_unsigned(17,8) ,
53373	 => std_logic_vector(to_unsigned(24,8) ,
53374	 => std_logic_vector(to_unsigned(35,8) ,
53375	 => std_logic_vector(to_unsigned(26,8) ,
53376	 => std_logic_vector(to_unsigned(27,8) ,
53377	 => std_logic_vector(to_unsigned(16,8) ,
53378	 => std_logic_vector(to_unsigned(1,8) ,
53379	 => std_logic_vector(to_unsigned(0,8) ,
53380	 => std_logic_vector(to_unsigned(3,8) ,
53381	 => std_logic_vector(to_unsigned(18,8) ,
53382	 => std_logic_vector(to_unsigned(14,8) ,
53383	 => std_logic_vector(to_unsigned(22,8) ,
53384	 => std_logic_vector(to_unsigned(18,8) ,
53385	 => std_logic_vector(to_unsigned(17,8) ,
53386	 => std_logic_vector(to_unsigned(15,8) ,
53387	 => std_logic_vector(to_unsigned(13,8) ,
53388	 => std_logic_vector(to_unsigned(15,8) ,
53389	 => std_logic_vector(to_unsigned(20,8) ,
53390	 => std_logic_vector(to_unsigned(16,8) ,
53391	 => std_logic_vector(to_unsigned(9,8) ,
53392	 => std_logic_vector(to_unsigned(10,8) ,
53393	 => std_logic_vector(to_unsigned(15,8) ,
53394	 => std_logic_vector(to_unsigned(11,8) ,
53395	 => std_logic_vector(to_unsigned(8,8) ,
53396	 => std_logic_vector(to_unsigned(10,8) ,
53397	 => std_logic_vector(to_unsigned(7,8) ,
53398	 => std_logic_vector(to_unsigned(7,8) ,
53399	 => std_logic_vector(to_unsigned(2,8) ,
53400	 => std_logic_vector(to_unsigned(0,8) ,
53401	 => std_logic_vector(to_unsigned(0,8) ,
53402	 => std_logic_vector(to_unsigned(0,8) ,
53403	 => std_logic_vector(to_unsigned(1,8) ,
53404	 => std_logic_vector(to_unsigned(9,8) ,
53405	 => std_logic_vector(to_unsigned(14,8) ,
53406	 => std_logic_vector(to_unsigned(12,8) ,
53407	 => std_logic_vector(to_unsigned(12,8) ,
53408	 => std_logic_vector(to_unsigned(7,8) ,
53409	 => std_logic_vector(to_unsigned(3,8) ,
53410	 => std_logic_vector(to_unsigned(13,8) ,
53411	 => std_logic_vector(to_unsigned(15,8) ,
53412	 => std_logic_vector(to_unsigned(22,8) ,
53413	 => std_logic_vector(to_unsigned(22,8) ,
53414	 => std_logic_vector(to_unsigned(17,8) ,
53415	 => std_logic_vector(to_unsigned(15,8) ,
53416	 => std_logic_vector(to_unsigned(20,8) ,
53417	 => std_logic_vector(to_unsigned(12,8) ,
53418	 => std_logic_vector(to_unsigned(10,8) ,
53419	 => std_logic_vector(to_unsigned(20,8) ,
53420	 => std_logic_vector(to_unsigned(41,8) ,
53421	 => std_logic_vector(to_unsigned(45,8) ,
53422	 => std_logic_vector(to_unsigned(35,8) ,
53423	 => std_logic_vector(to_unsigned(25,8) ,
53424	 => std_logic_vector(to_unsigned(29,8) ,
53425	 => std_logic_vector(to_unsigned(31,8) ,
53426	 => std_logic_vector(to_unsigned(24,8) ,
53427	 => std_logic_vector(to_unsigned(45,8) ,
53428	 => std_logic_vector(to_unsigned(34,8) ,
53429	 => std_logic_vector(to_unsigned(25,8) ,
53430	 => std_logic_vector(to_unsigned(13,8) ,
53431	 => std_logic_vector(to_unsigned(10,8) ,
53432	 => std_logic_vector(to_unsigned(19,8) ,
53433	 => std_logic_vector(to_unsigned(18,8) ,
53434	 => std_logic_vector(to_unsigned(13,8) ,
53435	 => std_logic_vector(to_unsigned(27,8) ,
53436	 => std_logic_vector(to_unsigned(56,8) ,
53437	 => std_logic_vector(to_unsigned(45,8) ,
53438	 => std_logic_vector(to_unsigned(46,8) ,
53439	 => std_logic_vector(to_unsigned(37,8) ,
53440	 => std_logic_vector(to_unsigned(59,8) ,
53441	 => std_logic_vector(to_unsigned(130,8) ,
53442	 => std_logic_vector(to_unsigned(134,8) ,
53443	 => std_logic_vector(to_unsigned(133,8) ,
53444	 => std_logic_vector(to_unsigned(115,8) ,
53445	 => std_logic_vector(to_unsigned(96,8) ,
53446	 => std_logic_vector(to_unsigned(103,8) ,
53447	 => std_logic_vector(to_unsigned(111,8) ,
53448	 => std_logic_vector(to_unsigned(119,8) ,
53449	 => std_logic_vector(to_unsigned(115,8) ,
53450	 => std_logic_vector(to_unsigned(105,8) ,
53451	 => std_logic_vector(to_unsigned(115,8) ,
53452	 => std_logic_vector(to_unsigned(125,8) ,
53453	 => std_logic_vector(to_unsigned(124,8) ,
53454	 => std_logic_vector(to_unsigned(114,8) ,
53455	 => std_logic_vector(to_unsigned(111,8) ,
53456	 => std_logic_vector(to_unsigned(124,8) ,
53457	 => std_logic_vector(to_unsigned(127,8) ,
53458	 => std_logic_vector(to_unsigned(111,8) ,
53459	 => std_logic_vector(to_unsigned(84,8) ,
53460	 => std_logic_vector(to_unsigned(78,8) ,
53461	 => std_logic_vector(to_unsigned(99,8) ,
53462	 => std_logic_vector(to_unsigned(59,8) ,
53463	 => std_logic_vector(to_unsigned(35,8) ,
53464	 => std_logic_vector(to_unsigned(49,8) ,
53465	 => std_logic_vector(to_unsigned(51,8) ,
53466	 => std_logic_vector(to_unsigned(60,8) ,
53467	 => std_logic_vector(to_unsigned(88,8) ,
53468	 => std_logic_vector(to_unsigned(92,8) ,
53469	 => std_logic_vector(to_unsigned(74,8) ,
53470	 => std_logic_vector(to_unsigned(64,8) ,
53471	 => std_logic_vector(to_unsigned(65,8) ,
53472	 => std_logic_vector(to_unsigned(68,8) ,
53473	 => std_logic_vector(to_unsigned(49,8) ,
53474	 => std_logic_vector(to_unsigned(45,8) ,
53475	 => std_logic_vector(to_unsigned(30,8) ,
53476	 => std_logic_vector(to_unsigned(23,8) ,
53477	 => std_logic_vector(to_unsigned(25,8) ,
53478	 => std_logic_vector(to_unsigned(29,8) ,
53479	 => std_logic_vector(to_unsigned(37,8) ,
53480	 => std_logic_vector(to_unsigned(53,8) ,
53481	 => std_logic_vector(to_unsigned(63,8) ,
53482	 => std_logic_vector(to_unsigned(67,8) ,
53483	 => std_logic_vector(to_unsigned(67,8) ,
53484	 => std_logic_vector(to_unsigned(66,8) ,
53485	 => std_logic_vector(to_unsigned(66,8) ,
53486	 => std_logic_vector(to_unsigned(62,8) ,
53487	 => std_logic_vector(to_unsigned(53,8) ,
53488	 => std_logic_vector(to_unsigned(49,8) ,
53489	 => std_logic_vector(to_unsigned(73,8) ,
53490	 => std_logic_vector(to_unsigned(87,8) ,
53491	 => std_logic_vector(to_unsigned(76,8) ,
53492	 => std_logic_vector(to_unsigned(101,8) ,
53493	 => std_logic_vector(to_unsigned(91,8) ,
53494	 => std_logic_vector(to_unsigned(81,8) ,
53495	 => std_logic_vector(to_unsigned(88,8) ,
53496	 => std_logic_vector(to_unsigned(92,8) ,
53497	 => std_logic_vector(to_unsigned(91,8) ,
53498	 => std_logic_vector(to_unsigned(78,8) ,
53499	 => std_logic_vector(to_unsigned(74,8) ,
53500	 => std_logic_vector(to_unsigned(79,8) ,
53501	 => std_logic_vector(to_unsigned(76,8) ,
53502	 => std_logic_vector(to_unsigned(85,8) ,
53503	 => std_logic_vector(to_unsigned(85,8) ,
53504	 => std_logic_vector(to_unsigned(65,8) ,
53505	 => std_logic_vector(to_unsigned(54,8) ,
53506	 => std_logic_vector(to_unsigned(65,8) ,
53507	 => std_logic_vector(to_unsigned(82,8) ,
53508	 => std_logic_vector(to_unsigned(96,8) ,
53509	 => std_logic_vector(to_unsigned(60,8) ,
53510	 => std_logic_vector(to_unsigned(104,8) ,
53511	 => std_logic_vector(to_unsigned(146,8) ,
53512	 => std_logic_vector(to_unsigned(136,8) ,
53513	 => std_logic_vector(to_unsigned(105,8) ,
53514	 => std_logic_vector(to_unsigned(74,8) ,
53515	 => std_logic_vector(to_unsigned(64,8) ,
53516	 => std_logic_vector(to_unsigned(64,8) ,
53517	 => std_logic_vector(to_unsigned(84,8) ,
53518	 => std_logic_vector(to_unsigned(96,8) ,
53519	 => std_logic_vector(to_unsigned(85,8) ,
53520	 => std_logic_vector(to_unsigned(74,8) ,
53521	 => std_logic_vector(to_unsigned(35,8) ,
53522	 => std_logic_vector(to_unsigned(28,8) ,
53523	 => std_logic_vector(to_unsigned(35,8) ,
53524	 => std_logic_vector(to_unsigned(27,8) ,
53525	 => std_logic_vector(to_unsigned(29,8) ,
53526	 => std_logic_vector(to_unsigned(27,8) ,
53527	 => std_logic_vector(to_unsigned(32,8) ,
53528	 => std_logic_vector(to_unsigned(43,8) ,
53529	 => std_logic_vector(to_unsigned(42,8) ,
53530	 => std_logic_vector(to_unsigned(50,8) ,
53531	 => std_logic_vector(to_unsigned(63,8) ,
53532	 => std_logic_vector(to_unsigned(65,8) ,
53533	 => std_logic_vector(to_unsigned(71,8) ,
53534	 => std_logic_vector(to_unsigned(97,8) ,
53535	 => std_logic_vector(to_unsigned(124,8) ,
53536	 => std_logic_vector(to_unsigned(111,8) ,
53537	 => std_logic_vector(to_unsigned(96,8) ,
53538	 => std_logic_vector(to_unsigned(112,8) ,
53539	 => std_logic_vector(to_unsigned(114,8) ,
53540	 => std_logic_vector(to_unsigned(105,8) ,
53541	 => std_logic_vector(to_unsigned(93,8) ,
53542	 => std_logic_vector(to_unsigned(71,8) ,
53543	 => std_logic_vector(to_unsigned(65,8) ,
53544	 => std_logic_vector(to_unsigned(67,8) ,
53545	 => std_logic_vector(to_unsigned(66,8) ,
53546	 => std_logic_vector(to_unsigned(51,8) ,
53547	 => std_logic_vector(to_unsigned(35,8) ,
53548	 => std_logic_vector(to_unsigned(35,8) ,
53549	 => std_logic_vector(to_unsigned(38,8) ,
53550	 => std_logic_vector(to_unsigned(39,8) ,
53551	 => std_logic_vector(to_unsigned(35,8) ,
53552	 => std_logic_vector(to_unsigned(34,8) ,
53553	 => std_logic_vector(to_unsigned(37,8) ,
53554	 => std_logic_vector(to_unsigned(45,8) ,
53555	 => std_logic_vector(to_unsigned(43,8) ,
53556	 => std_logic_vector(to_unsigned(43,8) ,
53557	 => std_logic_vector(to_unsigned(37,8) ,
53558	 => std_logic_vector(to_unsigned(32,8) ,
53559	 => std_logic_vector(to_unsigned(22,8) ,
53560	 => std_logic_vector(to_unsigned(19,8) ,
53561	 => std_logic_vector(to_unsigned(17,8) ,
53562	 => std_logic_vector(to_unsigned(15,8) ,
53563	 => std_logic_vector(to_unsigned(27,8) ,
53564	 => std_logic_vector(to_unsigned(62,8) ,
53565	 => std_logic_vector(to_unsigned(70,8) ,
53566	 => std_logic_vector(to_unsigned(44,8) ,
53567	 => std_logic_vector(to_unsigned(38,8) ,
53568	 => std_logic_vector(to_unsigned(41,8) ,
53569	 => std_logic_vector(to_unsigned(54,8) ,
53570	 => std_logic_vector(to_unsigned(30,8) ,
53571	 => std_logic_vector(to_unsigned(13,8) ,
53572	 => std_logic_vector(to_unsigned(20,8) ,
53573	 => std_logic_vector(to_unsigned(18,8) ,
53574	 => std_logic_vector(to_unsigned(15,8) ,
53575	 => std_logic_vector(to_unsigned(16,8) ,
53576	 => std_logic_vector(to_unsigned(17,8) ,
53577	 => std_logic_vector(to_unsigned(19,8) ,
53578	 => std_logic_vector(to_unsigned(12,8) ,
53579	 => std_logic_vector(to_unsigned(9,8) ,
53580	 => std_logic_vector(to_unsigned(6,8) ,
53581	 => std_logic_vector(to_unsigned(22,8) ,
53582	 => std_logic_vector(to_unsigned(63,8) ,
53583	 => std_logic_vector(to_unsigned(22,8) ,
53584	 => std_logic_vector(to_unsigned(29,8) ,
53585	 => std_logic_vector(to_unsigned(67,8) ,
53586	 => std_logic_vector(to_unsigned(29,8) ,
53587	 => std_logic_vector(to_unsigned(19,8) ,
53588	 => std_logic_vector(to_unsigned(24,8) ,
53589	 => std_logic_vector(to_unsigned(33,8) ,
53590	 => std_logic_vector(to_unsigned(64,8) ,
53591	 => std_logic_vector(to_unsigned(31,8) ,
53592	 => std_logic_vector(to_unsigned(42,8) ,
53593	 => std_logic_vector(to_unsigned(42,8) ,
53594	 => std_logic_vector(to_unsigned(41,8) ,
53595	 => std_logic_vector(to_unsigned(22,8) ,
53596	 => std_logic_vector(to_unsigned(45,8) ,
53597	 => std_logic_vector(to_unsigned(48,8) ,
53598	 => std_logic_vector(to_unsigned(12,8) ,
53599	 => std_logic_vector(to_unsigned(8,8) ,
53600	 => std_logic_vector(to_unsigned(6,8) ,
53601	 => std_logic_vector(to_unsigned(38,8) ,
53602	 => std_logic_vector(to_unsigned(38,8) ,
53603	 => std_logic_vector(to_unsigned(35,8) ,
53604	 => std_logic_vector(to_unsigned(45,8) ,
53605	 => std_logic_vector(to_unsigned(41,8) ,
53606	 => std_logic_vector(to_unsigned(39,8) ,
53607	 => std_logic_vector(to_unsigned(34,8) ,
53608	 => std_logic_vector(to_unsigned(39,8) ,
53609	 => std_logic_vector(to_unsigned(17,8) ,
53610	 => std_logic_vector(to_unsigned(8,8) ,
53611	 => std_logic_vector(to_unsigned(4,8) ,
53612	 => std_logic_vector(to_unsigned(10,8) ,
53613	 => std_logic_vector(to_unsigned(61,8) ,
53614	 => std_logic_vector(to_unsigned(31,8) ,
53615	 => std_logic_vector(to_unsigned(20,8) ,
53616	 => std_logic_vector(to_unsigned(18,8) ,
53617	 => std_logic_vector(to_unsigned(19,8) ,
53618	 => std_logic_vector(to_unsigned(17,8) ,
53619	 => std_logic_vector(to_unsigned(14,8) ,
53620	 => std_logic_vector(to_unsigned(17,8) ,
53621	 => std_logic_vector(to_unsigned(20,8) ,
53622	 => std_logic_vector(to_unsigned(19,8) ,
53623	 => std_logic_vector(to_unsigned(22,8) ,
53624	 => std_logic_vector(to_unsigned(22,8) ,
53625	 => std_logic_vector(to_unsigned(27,8) ,
53626	 => std_logic_vector(to_unsigned(32,8) ,
53627	 => std_logic_vector(to_unsigned(41,8) ,
53628	 => std_logic_vector(to_unsigned(26,8) ,
53629	 => std_logic_vector(to_unsigned(9,8) ,
53630	 => std_logic_vector(to_unsigned(12,8) ,
53631	 => std_logic_vector(to_unsigned(30,8) ,
53632	 => std_logic_vector(to_unsigned(17,8) ,
53633	 => std_logic_vector(to_unsigned(10,8) ,
53634	 => std_logic_vector(to_unsigned(22,8) ,
53635	 => std_logic_vector(to_unsigned(26,8) ,
53636	 => std_logic_vector(to_unsigned(18,8) ,
53637	 => std_logic_vector(to_unsigned(9,8) ,
53638	 => std_logic_vector(to_unsigned(6,8) ,
53639	 => std_logic_vector(to_unsigned(10,8) ,
53640	 => std_logic_vector(to_unsigned(18,8) ,
53641	 => std_logic_vector(to_unsigned(8,8) ,
53642	 => std_logic_vector(to_unsigned(9,8) ,
53643	 => std_logic_vector(to_unsigned(16,8) ,
53644	 => std_logic_vector(to_unsigned(17,8) ,
53645	 => std_logic_vector(to_unsigned(16,8) ,
53646	 => std_logic_vector(to_unsigned(30,8) ,
53647	 => std_logic_vector(to_unsigned(24,8) ,
53648	 => std_logic_vector(to_unsigned(18,8) ,
53649	 => std_logic_vector(to_unsigned(18,8) ,
53650	 => std_logic_vector(to_unsigned(15,8) ,
53651	 => std_logic_vector(to_unsigned(9,8) ,
53652	 => std_logic_vector(to_unsigned(6,8) ,
53653	 => std_logic_vector(to_unsigned(9,8) ,
53654	 => std_logic_vector(to_unsigned(15,8) ,
53655	 => std_logic_vector(to_unsigned(10,8) ,
53656	 => std_logic_vector(to_unsigned(12,8) ,
53657	 => std_logic_vector(to_unsigned(12,8) ,
53658	 => std_logic_vector(to_unsigned(20,8) ,
53659	 => std_logic_vector(to_unsigned(28,8) ,
53660	 => std_logic_vector(to_unsigned(12,8) ,
53661	 => std_logic_vector(to_unsigned(11,8) ,
53662	 => std_logic_vector(to_unsigned(34,8) ,
53663	 => std_logic_vector(to_unsigned(33,8) ,
53664	 => std_logic_vector(to_unsigned(22,8) ,
53665	 => std_logic_vector(to_unsigned(20,8) ,
53666	 => std_logic_vector(to_unsigned(20,8) ,
53667	 => std_logic_vector(to_unsigned(23,8) ,
53668	 => std_logic_vector(to_unsigned(19,8) ,
53669	 => std_logic_vector(to_unsigned(17,8) ,
53670	 => std_logic_vector(to_unsigned(31,8) ,
53671	 => std_logic_vector(to_unsigned(32,8) ,
53672	 => std_logic_vector(to_unsigned(25,8) ,
53673	 => std_logic_vector(to_unsigned(32,8) ,
53674	 => std_logic_vector(to_unsigned(22,8) ,
53675	 => std_logic_vector(to_unsigned(11,8) ,
53676	 => std_logic_vector(to_unsigned(22,8) ,
53677	 => std_logic_vector(to_unsigned(20,8) ,
53678	 => std_logic_vector(to_unsigned(16,8) ,
53679	 => std_logic_vector(to_unsigned(15,8) ,
53680	 => std_logic_vector(to_unsigned(18,8) ,
53681	 => std_logic_vector(to_unsigned(22,8) ,
53682	 => std_logic_vector(to_unsigned(24,8) ,
53683	 => std_logic_vector(to_unsigned(28,8) ,
53684	 => std_logic_vector(to_unsigned(29,8) ,
53685	 => std_logic_vector(to_unsigned(33,8) ,
53686	 => std_logic_vector(to_unsigned(39,8) ,
53687	 => std_logic_vector(to_unsigned(43,8) ,
53688	 => std_logic_vector(to_unsigned(42,8) ,
53689	 => std_logic_vector(to_unsigned(35,8) ,
53690	 => std_logic_vector(to_unsigned(39,8) ,
53691	 => std_logic_vector(to_unsigned(28,8) ,
53692	 => std_logic_vector(to_unsigned(22,8) ,
53693	 => std_logic_vector(to_unsigned(29,8) ,
53694	 => std_logic_vector(to_unsigned(29,8) ,
53695	 => std_logic_vector(to_unsigned(27,8) ,
53696	 => std_logic_vector(to_unsigned(25,8) ,
53697	 => std_logic_vector(to_unsigned(15,8) ,
53698	 => std_logic_vector(to_unsigned(2,8) ,
53699	 => std_logic_vector(to_unsigned(0,8) ,
53700	 => std_logic_vector(to_unsigned(2,8) ,
53701	 => std_logic_vector(to_unsigned(15,8) ,
53702	 => std_logic_vector(to_unsigned(15,8) ,
53703	 => std_logic_vector(to_unsigned(19,8) ,
53704	 => std_logic_vector(to_unsigned(12,8) ,
53705	 => std_logic_vector(to_unsigned(16,8) ,
53706	 => std_logic_vector(to_unsigned(13,8) ,
53707	 => std_logic_vector(to_unsigned(7,8) ,
53708	 => std_logic_vector(to_unsigned(8,8) ,
53709	 => std_logic_vector(to_unsigned(9,8) ,
53710	 => std_logic_vector(to_unsigned(9,8) ,
53711	 => std_logic_vector(to_unsigned(8,8) ,
53712	 => std_logic_vector(to_unsigned(9,8) ,
53713	 => std_logic_vector(to_unsigned(10,8) ,
53714	 => std_logic_vector(to_unsigned(7,8) ,
53715	 => std_logic_vector(to_unsigned(7,8) ,
53716	 => std_logic_vector(to_unsigned(7,8) ,
53717	 => std_logic_vector(to_unsigned(7,8) ,
53718	 => std_logic_vector(to_unsigned(10,8) ,
53719	 => std_logic_vector(to_unsigned(2,8) ,
53720	 => std_logic_vector(to_unsigned(0,8) ,
53721	 => std_logic_vector(to_unsigned(0,8) ,
53722	 => std_logic_vector(to_unsigned(0,8) ,
53723	 => std_logic_vector(to_unsigned(0,8) ,
53724	 => std_logic_vector(to_unsigned(10,8) ,
53725	 => std_logic_vector(to_unsigned(18,8) ,
53726	 => std_logic_vector(to_unsigned(12,8) ,
53727	 => std_logic_vector(to_unsigned(13,8) ,
53728	 => std_logic_vector(to_unsigned(18,8) ,
53729	 => std_logic_vector(to_unsigned(17,8) ,
53730	 => std_logic_vector(to_unsigned(17,8) ,
53731	 => std_logic_vector(to_unsigned(14,8) ,
53732	 => std_logic_vector(to_unsigned(23,8) ,
53733	 => std_logic_vector(to_unsigned(22,8) ,
53734	 => std_logic_vector(to_unsigned(14,8) ,
53735	 => std_logic_vector(to_unsigned(5,8) ,
53736	 => std_logic_vector(to_unsigned(4,8) ,
53737	 => std_logic_vector(to_unsigned(5,8) ,
53738	 => std_logic_vector(to_unsigned(6,8) ,
53739	 => std_logic_vector(to_unsigned(18,8) ,
53740	 => std_logic_vector(to_unsigned(36,8) ,
53741	 => std_logic_vector(to_unsigned(30,8) ,
53742	 => std_logic_vector(to_unsigned(30,8) ,
53743	 => std_logic_vector(to_unsigned(37,8) ,
53744	 => std_logic_vector(to_unsigned(40,8) ,
53745	 => std_logic_vector(to_unsigned(39,8) ,
53746	 => std_logic_vector(to_unsigned(32,8) ,
53747	 => std_logic_vector(to_unsigned(41,8) ,
53748	 => std_logic_vector(to_unsigned(21,8) ,
53749	 => std_logic_vector(to_unsigned(23,8) ,
53750	 => std_logic_vector(to_unsigned(23,8) ,
53751	 => std_logic_vector(to_unsigned(25,8) ,
53752	 => std_logic_vector(to_unsigned(36,8) ,
53753	 => std_logic_vector(to_unsigned(43,8) ,
53754	 => std_logic_vector(to_unsigned(44,8) ,
53755	 => std_logic_vector(to_unsigned(58,8) ,
53756	 => std_logic_vector(to_unsigned(82,8) ,
53757	 => std_logic_vector(to_unsigned(82,8) ,
53758	 => std_logic_vector(to_unsigned(70,8) ,
53759	 => std_logic_vector(to_unsigned(22,8) ,
53760	 => std_logic_vector(to_unsigned(44,8) ,
53761	 => std_logic_vector(to_unsigned(128,8) ,
53762	 => std_logic_vector(to_unsigned(114,8) ,
53763	 => std_logic_vector(to_unsigned(101,8) ,
53764	 => std_logic_vector(to_unsigned(108,8) ,
53765	 => std_logic_vector(to_unsigned(104,8) ,
53766	 => std_logic_vector(to_unsigned(104,8) ,
53767	 => std_logic_vector(to_unsigned(112,8) ,
53768	 => std_logic_vector(to_unsigned(118,8) ,
53769	 => std_logic_vector(to_unsigned(122,8) ,
53770	 => std_logic_vector(to_unsigned(121,8) ,
53771	 => std_logic_vector(to_unsigned(124,8) ,
53772	 => std_logic_vector(to_unsigned(130,8) ,
53773	 => std_logic_vector(to_unsigned(128,8) ,
53774	 => std_logic_vector(to_unsigned(114,8) ,
53775	 => std_logic_vector(to_unsigned(70,8) ,
53776	 => std_logic_vector(to_unsigned(88,8) ,
53777	 => std_logic_vector(to_unsigned(103,8) ,
53778	 => std_logic_vector(to_unsigned(82,8) ,
53779	 => std_logic_vector(to_unsigned(99,8) ,
53780	 => std_logic_vector(to_unsigned(108,8) ,
53781	 => std_logic_vector(to_unsigned(77,8) ,
53782	 => std_logic_vector(to_unsigned(64,8) ,
53783	 => std_logic_vector(to_unsigned(54,8) ,
53784	 => std_logic_vector(to_unsigned(71,8) ,
53785	 => std_logic_vector(to_unsigned(111,8) ,
53786	 => std_logic_vector(to_unsigned(80,8) ,
53787	 => std_logic_vector(to_unsigned(68,8) ,
53788	 => std_logic_vector(to_unsigned(56,8) ,
53789	 => std_logic_vector(to_unsigned(73,8) ,
53790	 => std_logic_vector(to_unsigned(108,8) ,
53791	 => std_logic_vector(to_unsigned(103,8) ,
53792	 => std_logic_vector(to_unsigned(82,8) ,
53793	 => std_logic_vector(to_unsigned(47,8) ,
53794	 => std_logic_vector(to_unsigned(38,8) ,
53795	 => std_logic_vector(to_unsigned(27,8) ,
53796	 => std_logic_vector(to_unsigned(22,8) ,
53797	 => std_logic_vector(to_unsigned(22,8) ,
53798	 => std_logic_vector(to_unsigned(29,8) ,
53799	 => std_logic_vector(to_unsigned(33,8) ,
53800	 => std_logic_vector(to_unsigned(36,8) ,
53801	 => std_logic_vector(to_unsigned(38,8) ,
53802	 => std_logic_vector(to_unsigned(45,8) ,
53803	 => std_logic_vector(to_unsigned(63,8) ,
53804	 => std_logic_vector(to_unsigned(72,8) ,
53805	 => std_logic_vector(to_unsigned(79,8) ,
53806	 => std_logic_vector(to_unsigned(77,8) ,
53807	 => std_logic_vector(to_unsigned(82,8) ,
53808	 => std_logic_vector(to_unsigned(80,8) ,
53809	 => std_logic_vector(to_unsigned(86,8) ,
53810	 => std_logic_vector(to_unsigned(97,8) ,
53811	 => std_logic_vector(to_unsigned(82,8) ,
53812	 => std_logic_vector(to_unsigned(101,8) ,
53813	 => std_logic_vector(to_unsigned(77,8) ,
53814	 => std_logic_vector(to_unsigned(63,8) ,
53815	 => std_logic_vector(to_unsigned(103,8) ,
53816	 => std_logic_vector(to_unsigned(88,8) ,
53817	 => std_logic_vector(to_unsigned(85,8) ,
53818	 => std_logic_vector(to_unsigned(90,8) ,
53819	 => std_logic_vector(to_unsigned(95,8) ,
53820	 => std_logic_vector(to_unsigned(101,8) ,
53821	 => std_logic_vector(to_unsigned(96,8) ,
53822	 => std_logic_vector(to_unsigned(92,8) ,
53823	 => std_logic_vector(to_unsigned(104,8) ,
53824	 => std_logic_vector(to_unsigned(99,8) ,
53825	 => std_logic_vector(to_unsigned(95,8) ,
53826	 => std_logic_vector(to_unsigned(84,8) ,
53827	 => std_logic_vector(to_unsigned(86,8) ,
53828	 => std_logic_vector(to_unsigned(90,8) ,
53829	 => std_logic_vector(to_unsigned(78,8) ,
53830	 => std_logic_vector(to_unsigned(119,8) ,
53831	 => std_logic_vector(to_unsigned(134,8) ,
53832	 => std_logic_vector(to_unsigned(96,8) ,
53833	 => std_logic_vector(to_unsigned(65,8) ,
53834	 => std_logic_vector(to_unsigned(61,8) ,
53835	 => std_logic_vector(to_unsigned(69,8) ,
53836	 => std_logic_vector(to_unsigned(69,8) ,
53837	 => std_logic_vector(to_unsigned(66,8) ,
53838	 => std_logic_vector(to_unsigned(84,8) ,
53839	 => std_logic_vector(to_unsigned(87,8) ,
53840	 => std_logic_vector(to_unsigned(93,8) ,
53841	 => std_logic_vector(to_unsigned(56,8) ,
53842	 => std_logic_vector(to_unsigned(18,8) ,
53843	 => std_logic_vector(to_unsigned(42,8) ,
53844	 => std_logic_vector(to_unsigned(37,8) ,
53845	 => std_logic_vector(to_unsigned(24,8) ,
53846	 => std_logic_vector(to_unsigned(24,8) ,
53847	 => std_logic_vector(to_unsigned(19,8) ,
53848	 => std_logic_vector(to_unsigned(18,8) ,
53849	 => std_logic_vector(to_unsigned(19,8) ,
53850	 => std_logic_vector(to_unsigned(39,8) ,
53851	 => std_logic_vector(to_unsigned(79,8) ,
53852	 => std_logic_vector(to_unsigned(66,8) ,
53853	 => std_logic_vector(to_unsigned(57,8) ,
53854	 => std_logic_vector(to_unsigned(68,8) ,
53855	 => std_logic_vector(to_unsigned(82,8) ,
53856	 => std_logic_vector(to_unsigned(88,8) ,
53857	 => std_logic_vector(to_unsigned(90,8) ,
53858	 => std_logic_vector(to_unsigned(88,8) ,
53859	 => std_logic_vector(to_unsigned(81,8) ,
53860	 => std_logic_vector(to_unsigned(71,8) ,
53861	 => std_logic_vector(to_unsigned(68,8) ,
53862	 => std_logic_vector(to_unsigned(67,8) ,
53863	 => std_logic_vector(to_unsigned(67,8) ,
53864	 => std_logic_vector(to_unsigned(65,8) ,
53865	 => std_logic_vector(to_unsigned(73,8) ,
53866	 => std_logic_vector(to_unsigned(65,8) ,
53867	 => std_logic_vector(to_unsigned(50,8) ,
53868	 => std_logic_vector(to_unsigned(35,8) ,
53869	 => std_logic_vector(to_unsigned(32,8) ,
53870	 => std_logic_vector(to_unsigned(32,8) ,
53871	 => std_logic_vector(to_unsigned(32,8) ,
53872	 => std_logic_vector(to_unsigned(36,8) ,
53873	 => std_logic_vector(to_unsigned(39,8) ,
53874	 => std_logic_vector(to_unsigned(39,8) ,
53875	 => std_logic_vector(to_unsigned(42,8) ,
53876	 => std_logic_vector(to_unsigned(36,8) ,
53877	 => std_logic_vector(to_unsigned(35,8) ,
53878	 => std_logic_vector(to_unsigned(31,8) ,
53879	 => std_logic_vector(to_unsigned(19,8) ,
53880	 => std_logic_vector(to_unsigned(14,8) ,
53881	 => std_logic_vector(to_unsigned(16,8) ,
53882	 => std_logic_vector(to_unsigned(17,8) ,
53883	 => std_logic_vector(to_unsigned(29,8) ,
53884	 => std_logic_vector(to_unsigned(62,8) ,
53885	 => std_logic_vector(to_unsigned(77,8) ,
53886	 => std_logic_vector(to_unsigned(48,8) ,
53887	 => std_logic_vector(to_unsigned(39,8) ,
53888	 => std_logic_vector(to_unsigned(39,8) ,
53889	 => std_logic_vector(to_unsigned(46,8) ,
53890	 => std_logic_vector(to_unsigned(27,8) ,
53891	 => std_logic_vector(to_unsigned(12,8) ,
53892	 => std_logic_vector(to_unsigned(16,8) ,
53893	 => std_logic_vector(to_unsigned(13,8) ,
53894	 => std_logic_vector(to_unsigned(13,8) ,
53895	 => std_logic_vector(to_unsigned(12,8) ,
53896	 => std_logic_vector(to_unsigned(12,8) ,
53897	 => std_logic_vector(to_unsigned(13,8) ,
53898	 => std_logic_vector(to_unsigned(11,8) ,
53899	 => std_logic_vector(to_unsigned(8,8) ,
53900	 => std_logic_vector(to_unsigned(7,8) ,
53901	 => std_logic_vector(to_unsigned(17,8) ,
53902	 => std_logic_vector(to_unsigned(65,8) ,
53903	 => std_logic_vector(to_unsigned(32,8) ,
53904	 => std_logic_vector(to_unsigned(34,8) ,
53905	 => std_logic_vector(to_unsigned(70,8) ,
53906	 => std_logic_vector(to_unsigned(26,8) ,
53907	 => std_logic_vector(to_unsigned(7,8) ,
53908	 => std_logic_vector(to_unsigned(5,8) ,
53909	 => std_logic_vector(to_unsigned(13,8) ,
53910	 => std_logic_vector(to_unsigned(48,8) ,
53911	 => std_logic_vector(to_unsigned(32,8) ,
53912	 => std_logic_vector(to_unsigned(51,8) ,
53913	 => std_logic_vector(to_unsigned(45,8) ,
53914	 => std_logic_vector(to_unsigned(42,8) ,
53915	 => std_logic_vector(to_unsigned(37,8) ,
53916	 => std_logic_vector(to_unsigned(47,8) ,
53917	 => std_logic_vector(to_unsigned(45,8) ,
53918	 => std_logic_vector(to_unsigned(29,8) ,
53919	 => std_logic_vector(to_unsigned(20,8) ,
53920	 => std_logic_vector(to_unsigned(17,8) ,
53921	 => std_logic_vector(to_unsigned(46,8) ,
53922	 => std_logic_vector(to_unsigned(30,8) ,
53923	 => std_logic_vector(to_unsigned(27,8) ,
53924	 => std_logic_vector(to_unsigned(28,8) ,
53925	 => std_logic_vector(to_unsigned(23,8) ,
53926	 => std_logic_vector(to_unsigned(23,8) ,
53927	 => std_logic_vector(to_unsigned(18,8) ,
53928	 => std_logic_vector(to_unsigned(34,8) ,
53929	 => std_logic_vector(to_unsigned(15,8) ,
53930	 => std_logic_vector(to_unsigned(7,8) ,
53931	 => std_logic_vector(to_unsigned(2,8) ,
53932	 => std_logic_vector(to_unsigned(7,8) ,
53933	 => std_logic_vector(to_unsigned(52,8) ,
53934	 => std_logic_vector(to_unsigned(23,8) ,
53935	 => std_logic_vector(to_unsigned(16,8) ,
53936	 => std_logic_vector(to_unsigned(15,8) ,
53937	 => std_logic_vector(to_unsigned(16,8) ,
53938	 => std_logic_vector(to_unsigned(17,8) ,
53939	 => std_logic_vector(to_unsigned(16,8) ,
53940	 => std_logic_vector(to_unsigned(15,8) ,
53941	 => std_logic_vector(to_unsigned(17,8) ,
53942	 => std_logic_vector(to_unsigned(18,8) ,
53943	 => std_logic_vector(to_unsigned(20,8) ,
53944	 => std_logic_vector(to_unsigned(19,8) ,
53945	 => std_logic_vector(to_unsigned(27,8) ,
53946	 => std_logic_vector(to_unsigned(41,8) ,
53947	 => std_logic_vector(to_unsigned(26,8) ,
53948	 => std_logic_vector(to_unsigned(13,8) ,
53949	 => std_logic_vector(to_unsigned(14,8) ,
53950	 => std_logic_vector(to_unsigned(13,8) ,
53951	 => std_logic_vector(to_unsigned(23,8) ,
53952	 => std_logic_vector(to_unsigned(15,8) ,
53953	 => std_logic_vector(to_unsigned(9,8) ,
53954	 => std_logic_vector(to_unsigned(23,8) ,
53955	 => std_logic_vector(to_unsigned(32,8) ,
53956	 => std_logic_vector(to_unsigned(22,8) ,
53957	 => std_logic_vector(to_unsigned(27,8) ,
53958	 => std_logic_vector(to_unsigned(29,8) ,
53959	 => std_logic_vector(to_unsigned(22,8) ,
53960	 => std_logic_vector(to_unsigned(24,8) ,
53961	 => std_logic_vector(to_unsigned(17,8) ,
53962	 => std_logic_vector(to_unsigned(19,8) ,
53963	 => std_logic_vector(to_unsigned(18,8) ,
53964	 => std_logic_vector(to_unsigned(16,8) ,
53965	 => std_logic_vector(to_unsigned(14,8) ,
53966	 => std_logic_vector(to_unsigned(44,8) ,
53967	 => std_logic_vector(to_unsigned(58,8) ,
53968	 => std_logic_vector(to_unsigned(41,8) ,
53969	 => std_logic_vector(to_unsigned(14,8) ,
53970	 => std_logic_vector(to_unsigned(8,8) ,
53971	 => std_logic_vector(to_unsigned(17,8) ,
53972	 => std_logic_vector(to_unsigned(24,8) ,
53973	 => std_logic_vector(to_unsigned(19,8) ,
53974	 => std_logic_vector(to_unsigned(10,8) ,
53975	 => std_logic_vector(to_unsigned(10,8) ,
53976	 => std_logic_vector(to_unsigned(8,8) ,
53977	 => std_logic_vector(to_unsigned(11,8) ,
53978	 => std_logic_vector(to_unsigned(25,8) ,
53979	 => std_logic_vector(to_unsigned(18,8) ,
53980	 => std_logic_vector(to_unsigned(12,8) ,
53981	 => std_logic_vector(to_unsigned(17,8) ,
53982	 => std_logic_vector(to_unsigned(33,8) ,
53983	 => std_logic_vector(to_unsigned(37,8) ,
53984	 => std_logic_vector(to_unsigned(28,8) ,
53985	 => std_logic_vector(to_unsigned(21,8) ,
53986	 => std_logic_vector(to_unsigned(25,8) ,
53987	 => std_logic_vector(to_unsigned(23,8) ,
53988	 => std_logic_vector(to_unsigned(21,8) ,
53989	 => std_logic_vector(to_unsigned(29,8) ,
53990	 => std_logic_vector(to_unsigned(34,8) ,
53991	 => std_logic_vector(to_unsigned(27,8) ,
53992	 => std_logic_vector(to_unsigned(26,8) ,
53993	 => std_logic_vector(to_unsigned(16,8) ,
53994	 => std_logic_vector(to_unsigned(9,8) ,
53995	 => std_logic_vector(to_unsigned(17,8) ,
53996	 => std_logic_vector(to_unsigned(24,8) ,
53997	 => std_logic_vector(to_unsigned(20,8) ,
53998	 => std_logic_vector(to_unsigned(10,8) ,
53999	 => std_logic_vector(to_unsigned(20,8) ,
54000	 => std_logic_vector(to_unsigned(19,8) ,
54001	 => std_logic_vector(to_unsigned(14,8) ,
54002	 => std_logic_vector(to_unsigned(16,8) ,
54003	 => std_logic_vector(to_unsigned(16,8) ,
54004	 => std_logic_vector(to_unsigned(16,8) ,
54005	 => std_logic_vector(to_unsigned(16,8) ,
54006	 => std_logic_vector(to_unsigned(22,8) ,
54007	 => std_logic_vector(to_unsigned(23,8) ,
54008	 => std_logic_vector(to_unsigned(21,8) ,
54009	 => std_logic_vector(to_unsigned(72,8) ,
54010	 => std_logic_vector(to_unsigned(81,8) ,
54011	 => std_logic_vector(to_unsigned(36,8) ,
54012	 => std_logic_vector(to_unsigned(35,8) ,
54013	 => std_logic_vector(to_unsigned(28,8) ,
54014	 => std_logic_vector(to_unsigned(22,8) ,
54015	 => std_logic_vector(to_unsigned(24,8) ,
54016	 => std_logic_vector(to_unsigned(18,8) ,
54017	 => std_logic_vector(to_unsigned(13,8) ,
54018	 => std_logic_vector(to_unsigned(5,8) ,
54019	 => std_logic_vector(to_unsigned(0,8) ,
54020	 => std_logic_vector(to_unsigned(0,8) ,
54021	 => std_logic_vector(to_unsigned(7,8) ,
54022	 => std_logic_vector(to_unsigned(12,8) ,
54023	 => std_logic_vector(to_unsigned(22,8) ,
54024	 => std_logic_vector(to_unsigned(14,8) ,
54025	 => std_logic_vector(to_unsigned(17,8) ,
54026	 => std_logic_vector(to_unsigned(12,8) ,
54027	 => std_logic_vector(to_unsigned(9,8) ,
54028	 => std_logic_vector(to_unsigned(12,8) ,
54029	 => std_logic_vector(to_unsigned(15,8) ,
54030	 => std_logic_vector(to_unsigned(10,8) ,
54031	 => std_logic_vector(to_unsigned(7,8) ,
54032	 => std_logic_vector(to_unsigned(9,8) ,
54033	 => std_logic_vector(to_unsigned(9,8) ,
54034	 => std_logic_vector(to_unsigned(6,8) ,
54035	 => std_logic_vector(to_unsigned(8,8) ,
54036	 => std_logic_vector(to_unsigned(7,8) ,
54037	 => std_logic_vector(to_unsigned(6,8) ,
54038	 => std_logic_vector(to_unsigned(8,8) ,
54039	 => std_logic_vector(to_unsigned(2,8) ,
54040	 => std_logic_vector(to_unsigned(0,8) ,
54041	 => std_logic_vector(to_unsigned(0,8) ,
54042	 => std_logic_vector(to_unsigned(0,8) ,
54043	 => std_logic_vector(to_unsigned(0,8) ,
54044	 => std_logic_vector(to_unsigned(3,8) ,
54045	 => std_logic_vector(to_unsigned(11,8) ,
54046	 => std_logic_vector(to_unsigned(8,8) ,
54047	 => std_logic_vector(to_unsigned(7,8) ,
54048	 => std_logic_vector(to_unsigned(8,8) ,
54049	 => std_logic_vector(to_unsigned(12,8) ,
54050	 => std_logic_vector(to_unsigned(17,8) ,
54051	 => std_logic_vector(to_unsigned(15,8) ,
54052	 => std_logic_vector(to_unsigned(29,8) ,
54053	 => std_logic_vector(to_unsigned(19,8) ,
54054	 => std_logic_vector(to_unsigned(19,8) ,
54055	 => std_logic_vector(to_unsigned(19,8) ,
54056	 => std_logic_vector(to_unsigned(14,8) ,
54057	 => std_logic_vector(to_unsigned(10,8) ,
54058	 => std_logic_vector(to_unsigned(7,8) ,
54059	 => std_logic_vector(to_unsigned(19,8) ,
54060	 => std_logic_vector(to_unsigned(37,8) ,
54061	 => std_logic_vector(to_unsigned(25,8) ,
54062	 => std_logic_vector(to_unsigned(27,8) ,
54063	 => std_logic_vector(to_unsigned(23,8) ,
54064	 => std_logic_vector(to_unsigned(18,8) ,
54065	 => std_logic_vector(to_unsigned(20,8) ,
54066	 => std_logic_vector(to_unsigned(19,8) ,
54067	 => std_logic_vector(to_unsigned(38,8) ,
54068	 => std_logic_vector(to_unsigned(17,8) ,
54069	 => std_logic_vector(to_unsigned(14,8) ,
54070	 => std_logic_vector(to_unsigned(5,8) ,
54071	 => std_logic_vector(to_unsigned(3,8) ,
54072	 => std_logic_vector(to_unsigned(13,8) ,
54073	 => std_logic_vector(to_unsigned(17,8) ,
54074	 => std_logic_vector(to_unsigned(29,8) ,
54075	 => std_logic_vector(to_unsigned(41,8) ,
54076	 => std_logic_vector(to_unsigned(27,8) ,
54077	 => std_logic_vector(to_unsigned(27,8) ,
54078	 => std_logic_vector(to_unsigned(54,8) ,
54079	 => std_logic_vector(to_unsigned(64,8) ,
54080	 => std_logic_vector(to_unsigned(82,8) ,
54081	 => std_logic_vector(to_unsigned(104,8) ,
54082	 => std_logic_vector(to_unsigned(88,8) ,
54083	 => std_logic_vector(to_unsigned(87,8) ,
54084	 => std_logic_vector(to_unsigned(87,8) ,
54085	 => std_logic_vector(to_unsigned(73,8) ,
54086	 => std_logic_vector(to_unsigned(61,8) ,
54087	 => std_logic_vector(to_unsigned(79,8) ,
54088	 => std_logic_vector(to_unsigned(95,8) ,
54089	 => std_logic_vector(to_unsigned(87,8) ,
54090	 => std_logic_vector(to_unsigned(101,8) ,
54091	 => std_logic_vector(to_unsigned(88,8) ,
54092	 => std_logic_vector(to_unsigned(96,8) ,
54093	 => std_logic_vector(to_unsigned(112,8) ,
54094	 => std_logic_vector(to_unsigned(87,8) ,
54095	 => std_logic_vector(to_unsigned(52,8) ,
54096	 => std_logic_vector(to_unsigned(74,8) ,
54097	 => std_logic_vector(to_unsigned(99,8) ,
54098	 => std_logic_vector(to_unsigned(96,8) ,
54099	 => std_logic_vector(to_unsigned(108,8) ,
54100	 => std_logic_vector(to_unsigned(104,8) ,
54101	 => std_logic_vector(to_unsigned(62,8) ,
54102	 => std_logic_vector(to_unsigned(50,8) ,
54103	 => std_logic_vector(to_unsigned(64,8) ,
54104	 => std_logic_vector(to_unsigned(66,8) ,
54105	 => std_logic_vector(to_unsigned(77,8) ,
54106	 => std_logic_vector(to_unsigned(62,8) ,
54107	 => std_logic_vector(to_unsigned(64,8) ,
54108	 => std_logic_vector(to_unsigned(85,8) ,
54109	 => std_logic_vector(to_unsigned(115,8) ,
54110	 => std_logic_vector(to_unsigned(128,8) ,
54111	 => std_logic_vector(to_unsigned(74,8) ,
54112	 => std_logic_vector(to_unsigned(43,8) ,
54113	 => std_logic_vector(to_unsigned(35,8) ,
54114	 => std_logic_vector(to_unsigned(37,8) ,
54115	 => std_logic_vector(to_unsigned(25,8) ,
54116	 => std_logic_vector(to_unsigned(17,8) ,
54117	 => std_logic_vector(to_unsigned(19,8) ,
54118	 => std_logic_vector(to_unsigned(25,8) ,
54119	 => std_logic_vector(to_unsigned(26,8) ,
54120	 => std_logic_vector(to_unsigned(32,8) ,
54121	 => std_logic_vector(to_unsigned(37,8) ,
54122	 => std_logic_vector(to_unsigned(32,8) ,
54123	 => std_logic_vector(to_unsigned(34,8) ,
54124	 => std_logic_vector(to_unsigned(36,8) ,
54125	 => std_logic_vector(to_unsigned(37,8) ,
54126	 => std_logic_vector(to_unsigned(45,8) ,
54127	 => std_logic_vector(to_unsigned(49,8) ,
54128	 => std_logic_vector(to_unsigned(58,8) ,
54129	 => std_logic_vector(to_unsigned(77,8) ,
54130	 => std_logic_vector(to_unsigned(97,8) ,
54131	 => std_logic_vector(to_unsigned(92,8) ,
54132	 => std_logic_vector(to_unsigned(104,8) ,
54133	 => std_logic_vector(to_unsigned(105,8) ,
54134	 => std_logic_vector(to_unsigned(101,8) ,
54135	 => std_logic_vector(to_unsigned(116,8) ,
54136	 => std_logic_vector(to_unsigned(95,8) ,
54137	 => std_logic_vector(to_unsigned(88,8) ,
54138	 => std_logic_vector(to_unsigned(104,8) ,
54139	 => std_logic_vector(to_unsigned(100,8) ,
54140	 => std_logic_vector(to_unsigned(111,8) ,
54141	 => std_logic_vector(to_unsigned(80,8) ,
54142	 => std_logic_vector(to_unsigned(92,8) ,
54143	 => std_logic_vector(to_unsigned(105,8) ,
54144	 => std_logic_vector(to_unsigned(78,8) ,
54145	 => std_logic_vector(to_unsigned(105,8) ,
54146	 => std_logic_vector(to_unsigned(108,8) ,
54147	 => std_logic_vector(to_unsigned(97,8) ,
54148	 => std_logic_vector(to_unsigned(93,8) ,
54149	 => std_logic_vector(to_unsigned(108,8) ,
54150	 => std_logic_vector(to_unsigned(104,8) ,
54151	 => std_logic_vector(to_unsigned(93,8) ,
54152	 => std_logic_vector(to_unsigned(85,8) ,
54153	 => std_logic_vector(to_unsigned(78,8) ,
54154	 => std_logic_vector(to_unsigned(95,8) ,
54155	 => std_logic_vector(to_unsigned(111,8) ,
54156	 => std_logic_vector(to_unsigned(82,8) ,
54157	 => std_logic_vector(to_unsigned(59,8) ,
54158	 => std_logic_vector(to_unsigned(96,8) ,
54159	 => std_logic_vector(to_unsigned(116,8) ,
54160	 => std_logic_vector(to_unsigned(92,8) ,
54161	 => std_logic_vector(to_unsigned(76,8) ,
54162	 => std_logic_vector(to_unsigned(30,8) ,
54163	 => std_logic_vector(to_unsigned(28,8) ,
54164	 => std_logic_vector(to_unsigned(33,8) ,
54165	 => std_logic_vector(to_unsigned(30,8) ,
54166	 => std_logic_vector(to_unsigned(23,8) ,
54167	 => std_logic_vector(to_unsigned(22,8) ,
54168	 => std_logic_vector(to_unsigned(27,8) ,
54169	 => std_logic_vector(to_unsigned(37,8) ,
54170	 => std_logic_vector(to_unsigned(53,8) ,
54171	 => std_logic_vector(to_unsigned(63,8) ,
54172	 => std_logic_vector(to_unsigned(62,8) ,
54173	 => std_logic_vector(to_unsigned(61,8) ,
54174	 => std_logic_vector(to_unsigned(67,8) ,
54175	 => std_logic_vector(to_unsigned(66,8) ,
54176	 => std_logic_vector(to_unsigned(65,8) ,
54177	 => std_logic_vector(to_unsigned(72,8) ,
54178	 => std_logic_vector(to_unsigned(69,8) ,
54179	 => std_logic_vector(to_unsigned(63,8) ,
54180	 => std_logic_vector(to_unsigned(72,8) ,
54181	 => std_logic_vector(to_unsigned(77,8) ,
54182	 => std_logic_vector(to_unsigned(76,8) ,
54183	 => std_logic_vector(to_unsigned(76,8) ,
54184	 => std_logic_vector(to_unsigned(77,8) ,
54185	 => std_logic_vector(to_unsigned(66,8) ,
54186	 => std_logic_vector(to_unsigned(66,8) ,
54187	 => std_logic_vector(to_unsigned(72,8) ,
54188	 => std_logic_vector(to_unsigned(49,8) ,
54189	 => std_logic_vector(to_unsigned(32,8) ,
54190	 => std_logic_vector(to_unsigned(33,8) ,
54191	 => std_logic_vector(to_unsigned(34,8) ,
54192	 => std_logic_vector(to_unsigned(29,8) ,
54193	 => std_logic_vector(to_unsigned(37,8) ,
54194	 => std_logic_vector(to_unsigned(40,8) ,
54195	 => std_logic_vector(to_unsigned(37,8) ,
54196	 => std_logic_vector(to_unsigned(35,8) ,
54197	 => std_logic_vector(to_unsigned(35,8) ,
54198	 => std_logic_vector(to_unsigned(30,8) ,
54199	 => std_logic_vector(to_unsigned(22,8) ,
54200	 => std_logic_vector(to_unsigned(14,8) ,
54201	 => std_logic_vector(to_unsigned(14,8) ,
54202	 => std_logic_vector(to_unsigned(17,8) ,
54203	 => std_logic_vector(to_unsigned(18,8) ,
54204	 => std_logic_vector(to_unsigned(49,8) ,
54205	 => std_logic_vector(to_unsigned(78,8) ,
54206	 => std_logic_vector(to_unsigned(48,8) ,
54207	 => std_logic_vector(to_unsigned(38,8) ,
54208	 => std_logic_vector(to_unsigned(38,8) ,
54209	 => std_logic_vector(to_unsigned(46,8) ,
54210	 => std_logic_vector(to_unsigned(23,8) ,
54211	 => std_logic_vector(to_unsigned(9,8) ,
54212	 => std_logic_vector(to_unsigned(13,8) ,
54213	 => std_logic_vector(to_unsigned(13,8) ,
54214	 => std_logic_vector(to_unsigned(13,8) ,
54215	 => std_logic_vector(to_unsigned(15,8) ,
54216	 => std_logic_vector(to_unsigned(13,8) ,
54217	 => std_logic_vector(to_unsigned(21,8) ,
54218	 => std_logic_vector(to_unsigned(20,8) ,
54219	 => std_logic_vector(to_unsigned(12,8) ,
54220	 => std_logic_vector(to_unsigned(8,8) ,
54221	 => std_logic_vector(to_unsigned(13,8) ,
54222	 => std_logic_vector(to_unsigned(60,8) ,
54223	 => std_logic_vector(to_unsigned(20,8) ,
54224	 => std_logic_vector(to_unsigned(20,8) ,
54225	 => std_logic_vector(to_unsigned(67,8) ,
54226	 => std_logic_vector(to_unsigned(43,8) ,
54227	 => std_logic_vector(to_unsigned(12,8) ,
54228	 => std_logic_vector(to_unsigned(9,8) ,
54229	 => std_logic_vector(to_unsigned(13,8) ,
54230	 => std_logic_vector(to_unsigned(42,8) ,
54231	 => std_logic_vector(to_unsigned(30,8) ,
54232	 => std_logic_vector(to_unsigned(41,8) ,
54233	 => std_logic_vector(to_unsigned(27,8) ,
54234	 => std_logic_vector(to_unsigned(29,8) ,
54235	 => std_logic_vector(to_unsigned(16,8) ,
54236	 => std_logic_vector(to_unsigned(34,8) ,
54237	 => std_logic_vector(to_unsigned(28,8) ,
54238	 => std_logic_vector(to_unsigned(8,8) ,
54239	 => std_logic_vector(to_unsigned(10,8) ,
54240	 => std_logic_vector(to_unsigned(9,8) ,
54241	 => std_logic_vector(to_unsigned(36,8) ,
54242	 => std_logic_vector(to_unsigned(40,8) ,
54243	 => std_logic_vector(to_unsigned(32,8) ,
54244	 => std_logic_vector(to_unsigned(32,8) ,
54245	 => std_logic_vector(to_unsigned(26,8) ,
54246	 => std_logic_vector(to_unsigned(24,8) ,
54247	 => std_logic_vector(to_unsigned(22,8) ,
54248	 => std_logic_vector(to_unsigned(36,8) ,
54249	 => std_logic_vector(to_unsigned(19,8) ,
54250	 => std_logic_vector(to_unsigned(9,8) ,
54251	 => std_logic_vector(to_unsigned(5,8) ,
54252	 => std_logic_vector(to_unsigned(9,8) ,
54253	 => std_logic_vector(to_unsigned(44,8) ,
54254	 => std_logic_vector(to_unsigned(18,8) ,
54255	 => std_logic_vector(to_unsigned(11,8) ,
54256	 => std_logic_vector(to_unsigned(14,8) ,
54257	 => std_logic_vector(to_unsigned(13,8) ,
54258	 => std_logic_vector(to_unsigned(17,8) ,
54259	 => std_logic_vector(to_unsigned(17,8) ,
54260	 => std_logic_vector(to_unsigned(16,8) ,
54261	 => std_logic_vector(to_unsigned(17,8) ,
54262	 => std_logic_vector(to_unsigned(15,8) ,
54263	 => std_logic_vector(to_unsigned(22,8) ,
54264	 => std_logic_vector(to_unsigned(22,8) ,
54265	 => std_logic_vector(to_unsigned(29,8) ,
54266	 => std_logic_vector(to_unsigned(27,8) ,
54267	 => std_logic_vector(to_unsigned(12,8) ,
54268	 => std_logic_vector(to_unsigned(13,8) ,
54269	 => std_logic_vector(to_unsigned(18,8) ,
54270	 => std_logic_vector(to_unsigned(19,8) ,
54271	 => std_logic_vector(to_unsigned(22,8) ,
54272	 => std_logic_vector(to_unsigned(13,8) ,
54273	 => std_logic_vector(to_unsigned(11,8) ,
54274	 => std_logic_vector(to_unsigned(34,8) ,
54275	 => std_logic_vector(to_unsigned(43,8) ,
54276	 => std_logic_vector(to_unsigned(20,8) ,
54277	 => std_logic_vector(to_unsigned(32,8) ,
54278	 => std_logic_vector(to_unsigned(33,8) ,
54279	 => std_logic_vector(to_unsigned(30,8) ,
54280	 => std_logic_vector(to_unsigned(25,8) ,
54281	 => std_logic_vector(to_unsigned(29,8) ,
54282	 => std_logic_vector(to_unsigned(29,8) ,
54283	 => std_logic_vector(to_unsigned(22,8) ,
54284	 => std_logic_vector(to_unsigned(20,8) ,
54285	 => std_logic_vector(to_unsigned(27,8) ,
54286	 => std_logic_vector(to_unsigned(41,8) ,
54287	 => std_logic_vector(to_unsigned(48,8) ,
54288	 => std_logic_vector(to_unsigned(42,8) ,
54289	 => std_logic_vector(to_unsigned(17,8) ,
54290	 => std_logic_vector(to_unsigned(10,8) ,
54291	 => std_logic_vector(to_unsigned(31,8) ,
54292	 => std_logic_vector(to_unsigned(71,8) ,
54293	 => std_logic_vector(to_unsigned(54,8) ,
54294	 => std_logic_vector(to_unsigned(10,8) ,
54295	 => std_logic_vector(to_unsigned(30,8) ,
54296	 => std_logic_vector(to_unsigned(50,8) ,
54297	 => std_logic_vector(to_unsigned(30,8) ,
54298	 => std_logic_vector(to_unsigned(12,8) ,
54299	 => std_logic_vector(to_unsigned(16,8) ,
54300	 => std_logic_vector(to_unsigned(15,8) ,
54301	 => std_logic_vector(to_unsigned(17,8) ,
54302	 => std_logic_vector(to_unsigned(29,8) ,
54303	 => std_logic_vector(to_unsigned(32,8) ,
54304	 => std_logic_vector(to_unsigned(23,8) ,
54305	 => std_logic_vector(to_unsigned(23,8) ,
54306	 => std_logic_vector(to_unsigned(25,8) ,
54307	 => std_logic_vector(to_unsigned(24,8) ,
54308	 => std_logic_vector(to_unsigned(29,8) ,
54309	 => std_logic_vector(to_unsigned(36,8) ,
54310	 => std_logic_vector(to_unsigned(32,8) ,
54311	 => std_logic_vector(to_unsigned(31,8) ,
54312	 => std_logic_vector(to_unsigned(17,8) ,
54313	 => std_logic_vector(to_unsigned(7,8) ,
54314	 => std_logic_vector(to_unsigned(16,8) ,
54315	 => std_logic_vector(to_unsigned(23,8) ,
54316	 => std_logic_vector(to_unsigned(15,8) ,
54317	 => std_logic_vector(to_unsigned(8,8) ,
54318	 => std_logic_vector(to_unsigned(8,8) ,
54319	 => std_logic_vector(to_unsigned(38,8) ,
54320	 => std_logic_vector(to_unsigned(69,8) ,
54321	 => std_logic_vector(to_unsigned(55,8) ,
54322	 => std_logic_vector(to_unsigned(39,8) ,
54323	 => std_logic_vector(to_unsigned(17,8) ,
54324	 => std_logic_vector(to_unsigned(19,8) ,
54325	 => std_logic_vector(to_unsigned(16,8) ,
54326	 => std_logic_vector(to_unsigned(13,8) ,
54327	 => std_logic_vector(to_unsigned(14,8) ,
54328	 => std_logic_vector(to_unsigned(19,8) ,
54329	 => std_logic_vector(to_unsigned(51,8) ,
54330	 => std_logic_vector(to_unsigned(24,8) ,
54331	 => std_logic_vector(to_unsigned(15,8) ,
54332	 => std_logic_vector(to_unsigned(22,8) ,
54333	 => std_logic_vector(to_unsigned(23,8) ,
54334	 => std_logic_vector(to_unsigned(23,8) ,
54335	 => std_logic_vector(to_unsigned(20,8) ,
54336	 => std_logic_vector(to_unsigned(21,8) ,
54337	 => std_logic_vector(to_unsigned(24,8) ,
54338	 => std_logic_vector(to_unsigned(16,8) ,
54339	 => std_logic_vector(to_unsigned(1,8) ,
54340	 => std_logic_vector(to_unsigned(0,8) ,
54341	 => std_logic_vector(to_unsigned(4,8) ,
54342	 => std_logic_vector(to_unsigned(12,8) ,
54343	 => std_logic_vector(to_unsigned(19,8) ,
54344	 => std_logic_vector(to_unsigned(15,8) ,
54345	 => std_logic_vector(to_unsigned(18,8) ,
54346	 => std_logic_vector(to_unsigned(10,8) ,
54347	 => std_logic_vector(to_unsigned(7,8) ,
54348	 => std_logic_vector(to_unsigned(9,8) ,
54349	 => std_logic_vector(to_unsigned(9,8) ,
54350	 => std_logic_vector(to_unsigned(9,8) ,
54351	 => std_logic_vector(to_unsigned(8,8) ,
54352	 => std_logic_vector(to_unsigned(9,8) ,
54353	 => std_logic_vector(to_unsigned(9,8) ,
54354	 => std_logic_vector(to_unsigned(8,8) ,
54355	 => std_logic_vector(to_unsigned(8,8) ,
54356	 => std_logic_vector(to_unsigned(9,8) ,
54357	 => std_logic_vector(to_unsigned(7,8) ,
54358	 => std_logic_vector(to_unsigned(10,8) ,
54359	 => std_logic_vector(to_unsigned(5,8) ,
54360	 => std_logic_vector(to_unsigned(0,8) ,
54361	 => std_logic_vector(to_unsigned(0,8) ,
54362	 => std_logic_vector(to_unsigned(0,8) ,
54363	 => std_logic_vector(to_unsigned(0,8) ,
54364	 => std_logic_vector(to_unsigned(1,8) ,
54365	 => std_logic_vector(to_unsigned(12,8) ,
54366	 => std_logic_vector(to_unsigned(11,8) ,
54367	 => std_logic_vector(to_unsigned(7,8) ,
54368	 => std_logic_vector(to_unsigned(4,8) ,
54369	 => std_logic_vector(to_unsigned(3,8) ,
54370	 => std_logic_vector(to_unsigned(10,8) ,
54371	 => std_logic_vector(to_unsigned(14,8) ,
54372	 => std_logic_vector(to_unsigned(22,8) ,
54373	 => std_logic_vector(to_unsigned(20,8) ,
54374	 => std_logic_vector(to_unsigned(15,8) ,
54375	 => std_logic_vector(to_unsigned(6,8) ,
54376	 => std_logic_vector(to_unsigned(8,8) ,
54377	 => std_logic_vector(to_unsigned(12,8) ,
54378	 => std_logic_vector(to_unsigned(9,8) ,
54379	 => std_logic_vector(to_unsigned(16,8) ,
54380	 => std_logic_vector(to_unsigned(29,8) ,
54381	 => std_logic_vector(to_unsigned(24,8) ,
54382	 => std_logic_vector(to_unsigned(24,8) ,
54383	 => std_logic_vector(to_unsigned(24,8) ,
54384	 => std_logic_vector(to_unsigned(30,8) ,
54385	 => std_logic_vector(to_unsigned(33,8) ,
54386	 => std_logic_vector(to_unsigned(30,8) ,
54387	 => std_logic_vector(to_unsigned(41,8) ,
54388	 => std_logic_vector(to_unsigned(33,8) ,
54389	 => std_logic_vector(to_unsigned(32,8) ,
54390	 => std_logic_vector(to_unsigned(25,8) ,
54391	 => std_logic_vector(to_unsigned(19,8) ,
54392	 => std_logic_vector(to_unsigned(27,8) ,
54393	 => std_logic_vector(to_unsigned(29,8) ,
54394	 => std_logic_vector(to_unsigned(23,8) ,
54395	 => std_logic_vector(to_unsigned(27,8) ,
54396	 => std_logic_vector(to_unsigned(14,8) ,
54397	 => std_logic_vector(to_unsigned(8,8) ,
54398	 => std_logic_vector(to_unsigned(20,8) ,
54399	 => std_logic_vector(to_unsigned(36,8) ,
54400	 => std_logic_vector(to_unsigned(70,8) ,
54401	 => std_logic_vector(to_unsigned(100,8) ,
54402	 => std_logic_vector(to_unsigned(101,8) ,
54403	 => std_logic_vector(to_unsigned(96,8) ,
54404	 => std_logic_vector(to_unsigned(72,8) ,
54405	 => std_logic_vector(to_unsigned(55,8) ,
54406	 => std_logic_vector(to_unsigned(40,8) ,
54407	 => std_logic_vector(to_unsigned(59,8) ,
54408	 => std_logic_vector(to_unsigned(72,8) ,
54409	 => std_logic_vector(to_unsigned(61,8) ,
54410	 => std_logic_vector(to_unsigned(69,8) ,
54411	 => std_logic_vector(to_unsigned(67,8) ,
54412	 => std_logic_vector(to_unsigned(72,8) ,
54413	 => std_logic_vector(to_unsigned(86,8) ,
54414	 => std_logic_vector(to_unsigned(79,8) ,
54415	 => std_logic_vector(to_unsigned(86,8) ,
54416	 => std_logic_vector(to_unsigned(92,8) ,
54417	 => std_logic_vector(to_unsigned(115,8) ,
54418	 => std_logic_vector(to_unsigned(107,8) ,
54419	 => std_logic_vector(to_unsigned(97,8) ,
54420	 => std_logic_vector(to_unsigned(72,8) ,
54421	 => std_logic_vector(to_unsigned(69,8) ,
54422	 => std_logic_vector(to_unsigned(41,8) ,
54423	 => std_logic_vector(to_unsigned(34,8) ,
54424	 => std_logic_vector(to_unsigned(47,8) ,
54425	 => std_logic_vector(to_unsigned(57,8) ,
54426	 => std_logic_vector(to_unsigned(91,8) ,
54427	 => std_logic_vector(to_unsigned(95,8) ,
54428	 => std_logic_vector(to_unsigned(92,8) ,
54429	 => std_logic_vector(to_unsigned(71,8) ,
54430	 => std_logic_vector(to_unsigned(51,8) ,
54431	 => std_logic_vector(to_unsigned(40,8) ,
54432	 => std_logic_vector(to_unsigned(48,8) ,
54433	 => std_logic_vector(to_unsigned(41,8) ,
54434	 => std_logic_vector(to_unsigned(31,8) ,
54435	 => std_logic_vector(to_unsigned(29,8) ,
54436	 => std_logic_vector(to_unsigned(17,8) ,
54437	 => std_logic_vector(to_unsigned(23,8) ,
54438	 => std_logic_vector(to_unsigned(24,8) ,
54439	 => std_logic_vector(to_unsigned(27,8) ,
54440	 => std_logic_vector(to_unsigned(32,8) ,
54441	 => std_logic_vector(to_unsigned(46,8) ,
54442	 => std_logic_vector(to_unsigned(41,8) ,
54443	 => std_logic_vector(to_unsigned(39,8) ,
54444	 => std_logic_vector(to_unsigned(49,8) ,
54445	 => std_logic_vector(to_unsigned(47,8) ,
54446	 => std_logic_vector(to_unsigned(52,8) ,
54447	 => std_logic_vector(to_unsigned(57,8) ,
54448	 => std_logic_vector(to_unsigned(50,8) ,
54449	 => std_logic_vector(to_unsigned(53,8) ,
54450	 => std_logic_vector(to_unsigned(88,8) ,
54451	 => std_logic_vector(to_unsigned(70,8) ,
54452	 => std_logic_vector(to_unsigned(84,8) ,
54453	 => std_logic_vector(to_unsigned(93,8) ,
54454	 => std_logic_vector(to_unsigned(76,8) ,
54455	 => std_logic_vector(to_unsigned(109,8) ,
54456	 => std_logic_vector(to_unsigned(88,8) ,
54457	 => std_logic_vector(to_unsigned(82,8) ,
54458	 => std_logic_vector(to_unsigned(104,8) ,
54459	 => std_logic_vector(to_unsigned(86,8) ,
54460	 => std_logic_vector(to_unsigned(114,8) ,
54461	 => std_logic_vector(to_unsigned(97,8) ,
54462	 => std_logic_vector(to_unsigned(108,8) ,
54463	 => std_logic_vector(to_unsigned(119,8) ,
54464	 => std_logic_vector(to_unsigned(93,8) ,
54465	 => std_logic_vector(to_unsigned(114,8) ,
54466	 => std_logic_vector(to_unsigned(108,8) ,
54467	 => std_logic_vector(to_unsigned(86,8) ,
54468	 => std_logic_vector(to_unsigned(93,8) ,
54469	 => std_logic_vector(to_unsigned(91,8) ,
54470	 => std_logic_vector(to_unsigned(74,8) ,
54471	 => std_logic_vector(to_unsigned(45,8) ,
54472	 => std_logic_vector(to_unsigned(92,8) ,
54473	 => std_logic_vector(to_unsigned(112,8) ,
54474	 => std_logic_vector(to_unsigned(108,8) ,
54475	 => std_logic_vector(to_unsigned(90,8) ,
54476	 => std_logic_vector(to_unsigned(57,8) ,
54477	 => std_logic_vector(to_unsigned(69,8) ,
54478	 => std_logic_vector(to_unsigned(116,8) ,
54479	 => std_logic_vector(to_unsigned(93,8) ,
54480	 => std_logic_vector(to_unsigned(66,8) ,
54481	 => std_logic_vector(to_unsigned(71,8) ,
54482	 => std_logic_vector(to_unsigned(55,8) ,
54483	 => std_logic_vector(to_unsigned(34,8) ,
54484	 => std_logic_vector(to_unsigned(29,8) ,
54485	 => std_logic_vector(to_unsigned(29,8) ,
54486	 => std_logic_vector(to_unsigned(34,8) ,
54487	 => std_logic_vector(to_unsigned(31,8) ,
54488	 => std_logic_vector(to_unsigned(30,8) ,
54489	 => std_logic_vector(to_unsigned(55,8) ,
54490	 => std_logic_vector(to_unsigned(59,8) ,
54491	 => std_logic_vector(to_unsigned(56,8) ,
54492	 => std_logic_vector(to_unsigned(63,8) ,
54493	 => std_logic_vector(to_unsigned(72,8) ,
54494	 => std_logic_vector(to_unsigned(73,8) ,
54495	 => std_logic_vector(to_unsigned(66,8) ,
54496	 => std_logic_vector(to_unsigned(66,8) ,
54497	 => std_logic_vector(to_unsigned(61,8) ,
54498	 => std_logic_vector(to_unsigned(62,8) ,
54499	 => std_logic_vector(to_unsigned(71,8) ,
54500	 => std_logic_vector(to_unsigned(77,8) ,
54501	 => std_logic_vector(to_unsigned(72,8) ,
54502	 => std_logic_vector(to_unsigned(76,8) ,
54503	 => std_logic_vector(to_unsigned(71,8) ,
54504	 => std_logic_vector(to_unsigned(69,8) ,
54505	 => std_logic_vector(to_unsigned(70,8) ,
54506	 => std_logic_vector(to_unsigned(68,8) ,
54507	 => std_logic_vector(to_unsigned(63,8) ,
54508	 => std_logic_vector(to_unsigned(62,8) ,
54509	 => std_logic_vector(to_unsigned(46,8) ,
54510	 => std_logic_vector(to_unsigned(37,8) ,
54511	 => std_logic_vector(to_unsigned(42,8) ,
54512	 => std_logic_vector(to_unsigned(38,8) ,
54513	 => std_logic_vector(to_unsigned(32,8) ,
54514	 => std_logic_vector(to_unsigned(31,8) ,
54515	 => std_logic_vector(to_unsigned(32,8) ,
54516	 => std_logic_vector(to_unsigned(31,8) ,
54517	 => std_logic_vector(to_unsigned(30,8) ,
54518	 => std_logic_vector(to_unsigned(29,8) ,
54519	 => std_logic_vector(to_unsigned(25,8) ,
54520	 => std_logic_vector(to_unsigned(17,8) ,
54521	 => std_logic_vector(to_unsigned(17,8) ,
54522	 => std_logic_vector(to_unsigned(17,8) ,
54523	 => std_logic_vector(to_unsigned(13,8) ,
54524	 => std_logic_vector(to_unsigned(40,8) ,
54525	 => std_logic_vector(to_unsigned(73,8) ,
54526	 => std_logic_vector(to_unsigned(43,8) ,
54527	 => std_logic_vector(to_unsigned(35,8) ,
54528	 => std_logic_vector(to_unsigned(35,8) ,
54529	 => std_logic_vector(to_unsigned(46,8) ,
54530	 => std_logic_vector(to_unsigned(23,8) ,
54531	 => std_logic_vector(to_unsigned(9,8) ,
54532	 => std_logic_vector(to_unsigned(12,8) ,
54533	 => std_logic_vector(to_unsigned(10,8) ,
54534	 => std_logic_vector(to_unsigned(10,8) ,
54535	 => std_logic_vector(to_unsigned(13,8) ,
54536	 => std_logic_vector(to_unsigned(17,8) ,
54537	 => std_logic_vector(to_unsigned(30,8) ,
54538	 => std_logic_vector(to_unsigned(31,8) ,
54539	 => std_logic_vector(to_unsigned(20,8) ,
54540	 => std_logic_vector(to_unsigned(10,8) ,
54541	 => std_logic_vector(to_unsigned(11,8) ,
54542	 => std_logic_vector(to_unsigned(48,8) ,
54543	 => std_logic_vector(to_unsigned(27,8) ,
54544	 => std_logic_vector(to_unsigned(24,8) ,
54545	 => std_logic_vector(to_unsigned(62,8) ,
54546	 => std_logic_vector(to_unsigned(46,8) ,
54547	 => std_logic_vector(to_unsigned(14,8) ,
54548	 => std_logic_vector(to_unsigned(8,8) ,
54549	 => std_logic_vector(to_unsigned(10,8) ,
54550	 => std_logic_vector(to_unsigned(47,8) ,
54551	 => std_logic_vector(to_unsigned(41,8) ,
54552	 => std_logic_vector(to_unsigned(40,8) ,
54553	 => std_logic_vector(to_unsigned(40,8) ,
54554	 => std_logic_vector(to_unsigned(43,8) ,
54555	 => std_logic_vector(to_unsigned(25,8) ,
54556	 => std_logic_vector(to_unsigned(41,8) ,
54557	 => std_logic_vector(to_unsigned(32,8) ,
54558	 => std_logic_vector(to_unsigned(7,8) ,
54559	 => std_logic_vector(to_unsigned(5,8) ,
54560	 => std_logic_vector(to_unsigned(3,8) ,
54561	 => std_logic_vector(to_unsigned(29,8) ,
54562	 => std_logic_vector(to_unsigned(30,8) ,
54563	 => std_logic_vector(to_unsigned(25,8) ,
54564	 => std_logic_vector(to_unsigned(35,8) ,
54565	 => std_logic_vector(to_unsigned(32,8) ,
54566	 => std_logic_vector(to_unsigned(28,8) ,
54567	 => std_logic_vector(to_unsigned(31,8) ,
54568	 => std_logic_vector(to_unsigned(32,8) ,
54569	 => std_logic_vector(to_unsigned(17,8) ,
54570	 => std_logic_vector(to_unsigned(22,8) ,
54571	 => std_logic_vector(to_unsigned(15,8) ,
54572	 => std_logic_vector(to_unsigned(18,8) ,
54573	 => std_logic_vector(to_unsigned(45,8) ,
54574	 => std_logic_vector(to_unsigned(20,8) ,
54575	 => std_logic_vector(to_unsigned(12,8) ,
54576	 => std_logic_vector(to_unsigned(16,8) ,
54577	 => std_logic_vector(to_unsigned(13,8) ,
54578	 => std_logic_vector(to_unsigned(15,8) ,
54579	 => std_logic_vector(to_unsigned(17,8) ,
54580	 => std_logic_vector(to_unsigned(19,8) ,
54581	 => std_logic_vector(to_unsigned(12,8) ,
54582	 => std_logic_vector(to_unsigned(12,8) ,
54583	 => std_logic_vector(to_unsigned(25,8) ,
54584	 => std_logic_vector(to_unsigned(25,8) ,
54585	 => std_logic_vector(to_unsigned(17,8) ,
54586	 => std_logic_vector(to_unsigned(14,8) ,
54587	 => std_logic_vector(to_unsigned(19,8) ,
54588	 => std_logic_vector(to_unsigned(19,8) ,
54589	 => std_logic_vector(to_unsigned(15,8) ,
54590	 => std_logic_vector(to_unsigned(16,8) ,
54591	 => std_logic_vector(to_unsigned(22,8) ,
54592	 => std_logic_vector(to_unsigned(20,8) ,
54593	 => std_logic_vector(to_unsigned(30,8) ,
54594	 => std_logic_vector(to_unsigned(44,8) ,
54595	 => std_logic_vector(to_unsigned(23,8) ,
54596	 => std_logic_vector(to_unsigned(15,8) ,
54597	 => std_logic_vector(to_unsigned(51,8) ,
54598	 => std_logic_vector(to_unsigned(55,8) ,
54599	 => std_logic_vector(to_unsigned(35,8) ,
54600	 => std_logic_vector(to_unsigned(19,8) ,
54601	 => std_logic_vector(to_unsigned(32,8) ,
54602	 => std_logic_vector(to_unsigned(35,8) ,
54603	 => std_logic_vector(to_unsigned(23,8) ,
54604	 => std_logic_vector(to_unsigned(17,8) ,
54605	 => std_logic_vector(to_unsigned(27,8) ,
54606	 => std_logic_vector(to_unsigned(22,8) ,
54607	 => std_logic_vector(to_unsigned(22,8) ,
54608	 => std_logic_vector(to_unsigned(27,8) ,
54609	 => std_logic_vector(to_unsigned(21,8) ,
54610	 => std_logic_vector(to_unsigned(13,8) ,
54611	 => std_logic_vector(to_unsigned(21,8) ,
54612	 => std_logic_vector(to_unsigned(45,8) ,
54613	 => std_logic_vector(to_unsigned(44,8) ,
54614	 => std_logic_vector(to_unsigned(14,8) ,
54615	 => std_logic_vector(to_unsigned(42,8) ,
54616	 => std_logic_vector(to_unsigned(77,8) ,
54617	 => std_logic_vector(to_unsigned(39,8) ,
54618	 => std_logic_vector(to_unsigned(8,8) ,
54619	 => std_logic_vector(to_unsigned(28,8) ,
54620	 => std_logic_vector(to_unsigned(18,8) ,
54621	 => std_logic_vector(to_unsigned(18,8) ,
54622	 => std_logic_vector(to_unsigned(26,8) ,
54623	 => std_logic_vector(to_unsigned(20,8) ,
54624	 => std_logic_vector(to_unsigned(13,8) ,
54625	 => std_logic_vector(to_unsigned(12,8) ,
54626	 => std_logic_vector(to_unsigned(15,8) ,
54627	 => std_logic_vector(to_unsigned(26,8) ,
54628	 => std_logic_vector(to_unsigned(34,8) ,
54629	 => std_logic_vector(to_unsigned(30,8) ,
54630	 => std_logic_vector(to_unsigned(36,8) ,
54631	 => std_logic_vector(to_unsigned(19,8) ,
54632	 => std_logic_vector(to_unsigned(8,8) ,
54633	 => std_logic_vector(to_unsigned(16,8) ,
54634	 => std_logic_vector(to_unsigned(25,8) ,
54635	 => std_logic_vector(to_unsigned(15,8) ,
54636	 => std_logic_vector(to_unsigned(10,8) ,
54637	 => std_logic_vector(to_unsigned(8,8) ,
54638	 => std_logic_vector(to_unsigned(7,8) ,
54639	 => std_logic_vector(to_unsigned(47,8) ,
54640	 => std_logic_vector(to_unsigned(95,8) ,
54641	 => std_logic_vector(to_unsigned(88,8) ,
54642	 => std_logic_vector(to_unsigned(43,8) ,
54643	 => std_logic_vector(to_unsigned(10,8) ,
54644	 => std_logic_vector(to_unsigned(17,8) ,
54645	 => std_logic_vector(to_unsigned(18,8) ,
54646	 => std_logic_vector(to_unsigned(20,8) ,
54647	 => std_logic_vector(to_unsigned(16,8) ,
54648	 => std_logic_vector(to_unsigned(19,8) ,
54649	 => std_logic_vector(to_unsigned(25,8) ,
54650	 => std_logic_vector(to_unsigned(12,8) ,
54651	 => std_logic_vector(to_unsigned(16,8) ,
54652	 => std_logic_vector(to_unsigned(12,8) ,
54653	 => std_logic_vector(to_unsigned(12,8) ,
54654	 => std_logic_vector(to_unsigned(17,8) ,
54655	 => std_logic_vector(to_unsigned(18,8) ,
54656	 => std_logic_vector(to_unsigned(17,8) ,
54657	 => std_logic_vector(to_unsigned(15,8) ,
54658	 => std_logic_vector(to_unsigned(17,8) ,
54659	 => std_logic_vector(to_unsigned(1,8) ,
54660	 => std_logic_vector(to_unsigned(0,8) ,
54661	 => std_logic_vector(to_unsigned(2,8) ,
54662	 => std_logic_vector(to_unsigned(9,8) ,
54663	 => std_logic_vector(to_unsigned(18,8) ,
54664	 => std_logic_vector(to_unsigned(15,8) ,
54665	 => std_logic_vector(to_unsigned(18,8) ,
54666	 => std_logic_vector(to_unsigned(11,8) ,
54667	 => std_logic_vector(to_unsigned(6,8) ,
54668	 => std_logic_vector(to_unsigned(8,8) ,
54669	 => std_logic_vector(to_unsigned(9,8) ,
54670	 => std_logic_vector(to_unsigned(8,8) ,
54671	 => std_logic_vector(to_unsigned(8,8) ,
54672	 => std_logic_vector(to_unsigned(7,8) ,
54673	 => std_logic_vector(to_unsigned(11,8) ,
54674	 => std_logic_vector(to_unsigned(8,8) ,
54675	 => std_logic_vector(to_unsigned(8,8) ,
54676	 => std_logic_vector(to_unsigned(7,8) ,
54677	 => std_logic_vector(to_unsigned(5,8) ,
54678	 => std_logic_vector(to_unsigned(8,8) ,
54679	 => std_logic_vector(to_unsigned(7,8) ,
54680	 => std_logic_vector(to_unsigned(1,8) ,
54681	 => std_logic_vector(to_unsigned(0,8) ,
54682	 => std_logic_vector(to_unsigned(0,8) ,
54683	 => std_logic_vector(to_unsigned(0,8) ,
54684	 => std_logic_vector(to_unsigned(1,8) ,
54685	 => std_logic_vector(to_unsigned(12,8) ,
54686	 => std_logic_vector(to_unsigned(15,8) ,
54687	 => std_logic_vector(to_unsigned(16,8) ,
54688	 => std_logic_vector(to_unsigned(19,8) ,
54689	 => std_logic_vector(to_unsigned(15,8) ,
54690	 => std_logic_vector(to_unsigned(17,8) ,
54691	 => std_logic_vector(to_unsigned(18,8) ,
54692	 => std_logic_vector(to_unsigned(17,8) ,
54693	 => std_logic_vector(to_unsigned(16,8) ,
54694	 => std_logic_vector(to_unsigned(13,8) ,
54695	 => std_logic_vector(to_unsigned(8,8) ,
54696	 => std_logic_vector(to_unsigned(4,8) ,
54697	 => std_logic_vector(to_unsigned(4,8) ,
54698	 => std_logic_vector(to_unsigned(5,8) ,
54699	 => std_logic_vector(to_unsigned(17,8) ,
54700	 => std_logic_vector(to_unsigned(13,8) ,
54701	 => std_logic_vector(to_unsigned(10,8) ,
54702	 => std_logic_vector(to_unsigned(8,8) ,
54703	 => std_logic_vector(to_unsigned(5,8) ,
54704	 => std_logic_vector(to_unsigned(13,8) ,
54705	 => std_logic_vector(to_unsigned(21,8) ,
54706	 => std_logic_vector(to_unsigned(23,8) ,
54707	 => std_logic_vector(to_unsigned(40,8) ,
54708	 => std_logic_vector(to_unsigned(17,8) ,
54709	 => std_logic_vector(to_unsigned(30,8) ,
54710	 => std_logic_vector(to_unsigned(40,8) ,
54711	 => std_logic_vector(to_unsigned(43,8) ,
54712	 => std_logic_vector(to_unsigned(46,8) ,
54713	 => std_logic_vector(to_unsigned(35,8) ,
54714	 => std_logic_vector(to_unsigned(52,8) ,
54715	 => std_logic_vector(to_unsigned(58,8) ,
54716	 => std_logic_vector(to_unsigned(40,8) ,
54717	 => std_logic_vector(to_unsigned(47,8) ,
54718	 => std_logic_vector(to_unsigned(51,8) ,
54719	 => std_logic_vector(to_unsigned(41,8) ,
54720	 => std_logic_vector(to_unsigned(87,8) ,
54721	 => std_logic_vector(to_unsigned(80,8) ,
54722	 => std_logic_vector(to_unsigned(77,8) ,
54723	 => std_logic_vector(to_unsigned(92,8) ,
54724	 => std_logic_vector(to_unsigned(71,8) ,
54725	 => std_logic_vector(to_unsigned(47,8) ,
54726	 => std_logic_vector(to_unsigned(42,8) ,
54727	 => std_logic_vector(to_unsigned(72,8) ,
54728	 => std_logic_vector(to_unsigned(87,8) ,
54729	 => std_logic_vector(to_unsigned(72,8) ,
54730	 => std_logic_vector(to_unsigned(68,8) ,
54731	 => std_logic_vector(to_unsigned(80,8) ,
54732	 => std_logic_vector(to_unsigned(73,8) ,
54733	 => std_logic_vector(to_unsigned(81,8) ,
54734	 => std_logic_vector(to_unsigned(95,8) ,
54735	 => std_logic_vector(to_unsigned(103,8) ,
54736	 => std_logic_vector(to_unsigned(96,8) ,
54737	 => std_logic_vector(to_unsigned(91,8) ,
54738	 => std_logic_vector(to_unsigned(85,8) ,
54739	 => std_logic_vector(to_unsigned(80,8) ,
54740	 => std_logic_vector(to_unsigned(78,8) ,
54741	 => std_logic_vector(to_unsigned(55,8) ,
54742	 => std_logic_vector(to_unsigned(41,8) ,
54743	 => std_logic_vector(to_unsigned(67,8) ,
54744	 => std_logic_vector(to_unsigned(87,8) ,
54745	 => std_logic_vector(to_unsigned(85,8) ,
54746	 => std_logic_vector(to_unsigned(103,8) ,
54747	 => std_logic_vector(to_unsigned(65,8) ,
54748	 => std_logic_vector(to_unsigned(37,8) ,
54749	 => std_logic_vector(to_unsigned(37,8) ,
54750	 => std_logic_vector(to_unsigned(64,8) ,
54751	 => std_logic_vector(to_unsigned(80,8) ,
54752	 => std_logic_vector(to_unsigned(65,8) ,
54753	 => std_logic_vector(to_unsigned(44,8) ,
54754	 => std_logic_vector(to_unsigned(35,8) ,
54755	 => std_logic_vector(to_unsigned(24,8) ,
54756	 => std_logic_vector(to_unsigned(23,8) ,
54757	 => std_logic_vector(to_unsigned(32,8) ,
54758	 => std_logic_vector(to_unsigned(29,8) ,
54759	 => std_logic_vector(to_unsigned(32,8) ,
54760	 => std_logic_vector(to_unsigned(27,8) ,
54761	 => std_logic_vector(to_unsigned(41,8) ,
54762	 => std_logic_vector(to_unsigned(47,8) ,
54763	 => std_logic_vector(to_unsigned(38,8) ,
54764	 => std_logic_vector(to_unsigned(41,8) ,
54765	 => std_logic_vector(to_unsigned(41,8) ,
54766	 => std_logic_vector(to_unsigned(43,8) ,
54767	 => std_logic_vector(to_unsigned(56,8) ,
54768	 => std_logic_vector(to_unsigned(59,8) ,
54769	 => std_logic_vector(to_unsigned(55,8) ,
54770	 => std_logic_vector(to_unsigned(79,8) ,
54771	 => std_logic_vector(to_unsigned(81,8) ,
54772	 => std_logic_vector(to_unsigned(88,8) ,
54773	 => std_logic_vector(to_unsigned(91,8) ,
54774	 => std_logic_vector(to_unsigned(77,8) ,
54775	 => std_logic_vector(to_unsigned(95,8) ,
54776	 => std_logic_vector(to_unsigned(86,8) ,
54777	 => std_logic_vector(to_unsigned(76,8) ,
54778	 => std_logic_vector(to_unsigned(84,8) ,
54779	 => std_logic_vector(to_unsigned(71,8) ,
54780	 => std_logic_vector(to_unsigned(95,8) ,
54781	 => std_logic_vector(to_unsigned(67,8) ,
54782	 => std_logic_vector(to_unsigned(91,8) ,
54783	 => std_logic_vector(to_unsigned(115,8) ,
54784	 => std_logic_vector(to_unsigned(111,8) ,
54785	 => std_logic_vector(to_unsigned(121,8) ,
54786	 => std_logic_vector(to_unsigned(136,8) ,
54787	 => std_logic_vector(to_unsigned(109,8) ,
54788	 => std_logic_vector(to_unsigned(79,8) ,
54789	 => std_logic_vector(to_unsigned(82,8) ,
54790	 => std_logic_vector(to_unsigned(74,8) ,
54791	 => std_logic_vector(to_unsigned(50,8) ,
54792	 => std_logic_vector(to_unsigned(82,8) ,
54793	 => std_logic_vector(to_unsigned(100,8) ,
54794	 => std_logic_vector(to_unsigned(84,8) ,
54795	 => std_logic_vector(to_unsigned(74,8) ,
54796	 => std_logic_vector(to_unsigned(72,8) ,
54797	 => std_logic_vector(to_unsigned(72,8) ,
54798	 => std_logic_vector(to_unsigned(85,8) ,
54799	 => std_logic_vector(to_unsigned(67,8) ,
54800	 => std_logic_vector(to_unsigned(53,8) ,
54801	 => std_logic_vector(to_unsigned(54,8) ,
54802	 => std_logic_vector(to_unsigned(46,8) ,
54803	 => std_logic_vector(to_unsigned(60,8) ,
54804	 => std_logic_vector(to_unsigned(58,8) ,
54805	 => std_logic_vector(to_unsigned(37,8) ,
54806	 => std_logic_vector(to_unsigned(32,8) ,
54807	 => std_logic_vector(to_unsigned(41,8) ,
54808	 => std_logic_vector(to_unsigned(44,8) ,
54809	 => std_logic_vector(to_unsigned(52,8) ,
54810	 => std_logic_vector(to_unsigned(51,8) ,
54811	 => std_logic_vector(to_unsigned(53,8) ,
54812	 => std_logic_vector(to_unsigned(57,8) ,
54813	 => std_logic_vector(to_unsigned(61,8) ,
54814	 => std_logic_vector(to_unsigned(54,8) ,
54815	 => std_logic_vector(to_unsigned(56,8) ,
54816	 => std_logic_vector(to_unsigned(65,8) ,
54817	 => std_logic_vector(to_unsigned(62,8) ,
54818	 => std_logic_vector(to_unsigned(64,8) ,
54819	 => std_logic_vector(to_unsigned(71,8) ,
54820	 => std_logic_vector(to_unsigned(71,8) ,
54821	 => std_logic_vector(to_unsigned(66,8) ,
54822	 => std_logic_vector(to_unsigned(62,8) ,
54823	 => std_logic_vector(to_unsigned(64,8) ,
54824	 => std_logic_vector(to_unsigned(65,8) ,
54825	 => std_logic_vector(to_unsigned(73,8) ,
54826	 => std_logic_vector(to_unsigned(69,8) ,
54827	 => std_logic_vector(to_unsigned(62,8) ,
54828	 => std_logic_vector(to_unsigned(63,8) ,
54829	 => std_logic_vector(to_unsigned(57,8) ,
54830	 => std_logic_vector(to_unsigned(45,8) ,
54831	 => std_logic_vector(to_unsigned(49,8) ,
54832	 => std_logic_vector(to_unsigned(51,8) ,
54833	 => std_logic_vector(to_unsigned(45,8) ,
54834	 => std_logic_vector(to_unsigned(39,8) ,
54835	 => std_logic_vector(to_unsigned(38,8) ,
54836	 => std_logic_vector(to_unsigned(33,8) ,
54837	 => std_logic_vector(to_unsigned(30,8) ,
54838	 => std_logic_vector(to_unsigned(32,8) ,
54839	 => std_logic_vector(to_unsigned(23,8) ,
54840	 => std_logic_vector(to_unsigned(14,8) ,
54841	 => std_logic_vector(to_unsigned(14,8) ,
54842	 => std_logic_vector(to_unsigned(17,8) ,
54843	 => std_logic_vector(to_unsigned(17,8) ,
54844	 => std_logic_vector(to_unsigned(44,8) ,
54845	 => std_logic_vector(to_unsigned(74,8) ,
54846	 => std_logic_vector(to_unsigned(41,8) ,
54847	 => std_logic_vector(to_unsigned(35,8) ,
54848	 => std_logic_vector(to_unsigned(35,8) ,
54849	 => std_logic_vector(to_unsigned(41,8) ,
54850	 => std_logic_vector(to_unsigned(39,8) ,
54851	 => std_logic_vector(to_unsigned(31,8) ,
54852	 => std_logic_vector(to_unsigned(30,8) ,
54853	 => std_logic_vector(to_unsigned(24,8) ,
54854	 => std_logic_vector(to_unsigned(19,8) ,
54855	 => std_logic_vector(to_unsigned(19,8) ,
54856	 => std_logic_vector(to_unsigned(27,8) ,
54857	 => std_logic_vector(to_unsigned(22,8) ,
54858	 => std_logic_vector(to_unsigned(21,8) ,
54859	 => std_logic_vector(to_unsigned(24,8) ,
54860	 => std_logic_vector(to_unsigned(10,8) ,
54861	 => std_logic_vector(to_unsigned(9,8) ,
54862	 => std_logic_vector(to_unsigned(46,8) ,
54863	 => std_logic_vector(to_unsigned(24,8) ,
54864	 => std_logic_vector(to_unsigned(25,8) ,
54865	 => std_logic_vector(to_unsigned(64,8) ,
54866	 => std_logic_vector(to_unsigned(49,8) ,
54867	 => std_logic_vector(to_unsigned(14,8) ,
54868	 => std_logic_vector(to_unsigned(7,8) ,
54869	 => std_logic_vector(to_unsigned(12,8) ,
54870	 => std_logic_vector(to_unsigned(35,8) ,
54871	 => std_logic_vector(to_unsigned(17,8) ,
54872	 => std_logic_vector(to_unsigned(30,8) ,
54873	 => std_logic_vector(to_unsigned(37,8) ,
54874	 => std_logic_vector(to_unsigned(39,8) ,
54875	 => std_logic_vector(to_unsigned(19,8) ,
54876	 => std_logic_vector(to_unsigned(37,8) ,
54877	 => std_logic_vector(to_unsigned(49,8) ,
54878	 => std_logic_vector(to_unsigned(9,8) ,
54879	 => std_logic_vector(to_unsigned(7,8) ,
54880	 => std_logic_vector(to_unsigned(6,8) ,
54881	 => std_logic_vector(to_unsigned(34,8) ,
54882	 => std_logic_vector(to_unsigned(41,8) ,
54883	 => std_logic_vector(to_unsigned(27,8) ,
54884	 => std_logic_vector(to_unsigned(30,8) ,
54885	 => std_logic_vector(to_unsigned(24,8) ,
54886	 => std_logic_vector(to_unsigned(25,8) ,
54887	 => std_logic_vector(to_unsigned(25,8) ,
54888	 => std_logic_vector(to_unsigned(27,8) ,
54889	 => std_logic_vector(to_unsigned(17,8) ,
54890	 => std_logic_vector(to_unsigned(43,8) ,
54891	 => std_logic_vector(to_unsigned(36,8) ,
54892	 => std_logic_vector(to_unsigned(18,8) ,
54893	 => std_logic_vector(to_unsigned(39,8) ,
54894	 => std_logic_vector(to_unsigned(20,8) ,
54895	 => std_logic_vector(to_unsigned(12,8) ,
54896	 => std_logic_vector(to_unsigned(13,8) ,
54897	 => std_logic_vector(to_unsigned(15,8) ,
54898	 => std_logic_vector(to_unsigned(16,8) ,
54899	 => std_logic_vector(to_unsigned(13,8) ,
54900	 => std_logic_vector(to_unsigned(13,8) ,
54901	 => std_logic_vector(to_unsigned(8,8) ,
54902	 => std_logic_vector(to_unsigned(12,8) ,
54903	 => std_logic_vector(to_unsigned(23,8) ,
54904	 => std_logic_vector(to_unsigned(12,8) ,
54905	 => std_logic_vector(to_unsigned(12,8) ,
54906	 => std_logic_vector(to_unsigned(30,8) ,
54907	 => std_logic_vector(to_unsigned(23,8) ,
54908	 => std_logic_vector(to_unsigned(8,8) ,
54909	 => std_logic_vector(to_unsigned(7,8) ,
54910	 => std_logic_vector(to_unsigned(14,8) ,
54911	 => std_logic_vector(to_unsigned(28,8) ,
54912	 => std_logic_vector(to_unsigned(49,8) ,
54913	 => std_logic_vector(to_unsigned(51,8) ,
54914	 => std_logic_vector(to_unsigned(17,8) ,
54915	 => std_logic_vector(to_unsigned(11,8) ,
54916	 => std_logic_vector(to_unsigned(22,8) ,
54917	 => std_logic_vector(to_unsigned(47,8) ,
54918	 => std_logic_vector(to_unsigned(64,8) ,
54919	 => std_logic_vector(to_unsigned(41,8) ,
54920	 => std_logic_vector(to_unsigned(17,8) ,
54921	 => std_logic_vector(to_unsigned(44,8) ,
54922	 => std_logic_vector(to_unsigned(72,8) ,
54923	 => std_logic_vector(to_unsigned(46,8) ,
54924	 => std_logic_vector(to_unsigned(17,8) ,
54925	 => std_logic_vector(to_unsigned(27,8) ,
54926	 => std_logic_vector(to_unsigned(19,8) ,
54927	 => std_logic_vector(to_unsigned(13,8) ,
54928	 => std_logic_vector(to_unsigned(13,8) ,
54929	 => std_logic_vector(to_unsigned(21,8) ,
54930	 => std_logic_vector(to_unsigned(17,8) ,
54931	 => std_logic_vector(to_unsigned(12,8) ,
54932	 => std_logic_vector(to_unsigned(12,8) ,
54933	 => std_logic_vector(to_unsigned(12,8) ,
54934	 => std_logic_vector(to_unsigned(17,8) ,
54935	 => std_logic_vector(to_unsigned(19,8) ,
54936	 => std_logic_vector(to_unsigned(29,8) ,
54937	 => std_logic_vector(to_unsigned(25,8) ,
54938	 => std_logic_vector(to_unsigned(15,8) ,
54939	 => std_logic_vector(to_unsigned(28,8) ,
54940	 => std_logic_vector(to_unsigned(16,8) ,
54941	 => std_logic_vector(to_unsigned(18,8) ,
54942	 => std_logic_vector(to_unsigned(31,8) ,
54943	 => std_logic_vector(to_unsigned(26,8) ,
54944	 => std_logic_vector(to_unsigned(9,8) ,
54945	 => std_logic_vector(to_unsigned(9,8) ,
54946	 => std_logic_vector(to_unsigned(19,8) ,
54947	 => std_logic_vector(to_unsigned(22,8) ,
54948	 => std_logic_vector(to_unsigned(24,8) ,
54949	 => std_logic_vector(to_unsigned(29,8) ,
54950	 => std_logic_vector(to_unsigned(23,8) ,
54951	 => std_logic_vector(to_unsigned(14,8) ,
54952	 => std_logic_vector(to_unsigned(16,8) ,
54953	 => std_logic_vector(to_unsigned(25,8) ,
54954	 => std_logic_vector(to_unsigned(25,8) ,
54955	 => std_logic_vector(to_unsigned(19,8) ,
54956	 => std_logic_vector(to_unsigned(11,8) ,
54957	 => std_logic_vector(to_unsigned(11,8) ,
54958	 => std_logic_vector(to_unsigned(12,8) ,
54959	 => std_logic_vector(to_unsigned(57,8) ,
54960	 => std_logic_vector(to_unsigned(93,8) ,
54961	 => std_logic_vector(to_unsigned(91,8) ,
54962	 => std_logic_vector(to_unsigned(34,8) ,
54963	 => std_logic_vector(to_unsigned(8,8) ,
54964	 => std_logic_vector(to_unsigned(18,8) ,
54965	 => std_logic_vector(to_unsigned(13,8) ,
54966	 => std_logic_vector(to_unsigned(13,8) ,
54967	 => std_logic_vector(to_unsigned(14,8) ,
54968	 => std_logic_vector(to_unsigned(16,8) ,
54969	 => std_logic_vector(to_unsigned(19,8) ,
54970	 => std_logic_vector(to_unsigned(14,8) ,
54971	 => std_logic_vector(to_unsigned(20,8) ,
54972	 => std_logic_vector(to_unsigned(16,8) ,
54973	 => std_logic_vector(to_unsigned(12,8) ,
54974	 => std_logic_vector(to_unsigned(14,8) ,
54975	 => std_logic_vector(to_unsigned(19,8) ,
54976	 => std_logic_vector(to_unsigned(12,8) ,
54977	 => std_logic_vector(to_unsigned(9,8) ,
54978	 => std_logic_vector(to_unsigned(14,8) ,
54979	 => std_logic_vector(to_unsigned(5,8) ,
54980	 => std_logic_vector(to_unsigned(0,8) ,
54981	 => std_logic_vector(to_unsigned(0,8) ,
54982	 => std_logic_vector(to_unsigned(7,8) ,
54983	 => std_logic_vector(to_unsigned(24,8) ,
54984	 => std_logic_vector(to_unsigned(13,8) ,
54985	 => std_logic_vector(to_unsigned(18,8) ,
54986	 => std_logic_vector(to_unsigned(9,8) ,
54987	 => std_logic_vector(to_unsigned(7,8) ,
54988	 => std_logic_vector(to_unsigned(10,8) ,
54989	 => std_logic_vector(to_unsigned(10,8) ,
54990	 => std_logic_vector(to_unsigned(8,8) ,
54991	 => std_logic_vector(to_unsigned(8,8) ,
54992	 => std_logic_vector(to_unsigned(8,8) ,
54993	 => std_logic_vector(to_unsigned(10,8) ,
54994	 => std_logic_vector(to_unsigned(10,8) ,
54995	 => std_logic_vector(to_unsigned(9,8) ,
54996	 => std_logic_vector(to_unsigned(7,8) ,
54997	 => std_logic_vector(to_unsigned(6,8) ,
54998	 => std_logic_vector(to_unsigned(7,8) ,
54999	 => std_logic_vector(to_unsigned(7,8) ,
55000	 => std_logic_vector(to_unsigned(1,8) ,
55001	 => std_logic_vector(to_unsigned(0,8) ,
55002	 => std_logic_vector(to_unsigned(0,8) ,
55003	 => std_logic_vector(to_unsigned(0,8) ,
55004	 => std_logic_vector(to_unsigned(0,8) ,
55005	 => std_logic_vector(to_unsigned(7,8) ,
55006	 => std_logic_vector(to_unsigned(11,8) ,
55007	 => std_logic_vector(to_unsigned(9,8) ,
55008	 => std_logic_vector(to_unsigned(15,8) ,
55009	 => std_logic_vector(to_unsigned(22,8) ,
55010	 => std_logic_vector(to_unsigned(24,8) ,
55011	 => std_logic_vector(to_unsigned(23,8) ,
55012	 => std_logic_vector(to_unsigned(23,8) ,
55013	 => std_logic_vector(to_unsigned(19,8) ,
55014	 => std_logic_vector(to_unsigned(17,8) ,
55015	 => std_logic_vector(to_unsigned(17,8) ,
55016	 => std_logic_vector(to_unsigned(15,8) ,
55017	 => std_logic_vector(to_unsigned(10,8) ,
55018	 => std_logic_vector(to_unsigned(6,8) ,
55019	 => std_logic_vector(to_unsigned(16,8) ,
55020	 => std_logic_vector(to_unsigned(29,8) ,
55021	 => std_logic_vector(to_unsigned(24,8) ,
55022	 => std_logic_vector(to_unsigned(21,8) ,
55023	 => std_logic_vector(to_unsigned(17,8) ,
55024	 => std_logic_vector(to_unsigned(18,8) ,
55025	 => std_logic_vector(to_unsigned(17,8) ,
55026	 => std_logic_vector(to_unsigned(23,8) ,
55027	 => std_logic_vector(to_unsigned(39,8) ,
55028	 => std_logic_vector(to_unsigned(22,8) ,
55029	 => std_logic_vector(to_unsigned(25,8) ,
55030	 => std_logic_vector(to_unsigned(19,8) ,
55031	 => std_logic_vector(to_unsigned(22,8) ,
55032	 => std_logic_vector(to_unsigned(24,8) ,
55033	 => std_logic_vector(to_unsigned(15,8) ,
55034	 => std_logic_vector(to_unsigned(22,8) ,
55035	 => std_logic_vector(to_unsigned(29,8) ,
55036	 => std_logic_vector(to_unsigned(7,8) ,
55037	 => std_logic_vector(to_unsigned(6,8) ,
55038	 => std_logic_vector(to_unsigned(38,8) ,
55039	 => std_logic_vector(to_unsigned(60,8) ,
55040	 => std_logic_vector(to_unsigned(91,8) ,
55041	 => std_logic_vector(to_unsigned(82,8) ,
55042	 => std_logic_vector(to_unsigned(70,8) ,
55043	 => std_logic_vector(to_unsigned(87,8) ,
55044	 => std_logic_vector(to_unsigned(84,8) ,
55045	 => std_logic_vector(to_unsigned(59,8) ,
55046	 => std_logic_vector(to_unsigned(32,8) ,
55047	 => std_logic_vector(to_unsigned(66,8) ,
55048	 => std_logic_vector(to_unsigned(105,8) ,
55049	 => std_logic_vector(to_unsigned(73,8) ,
55050	 => std_logic_vector(to_unsigned(73,8) ,
55051	 => std_logic_vector(to_unsigned(90,8) ,
55052	 => std_logic_vector(to_unsigned(84,8) ,
55053	 => std_logic_vector(to_unsigned(96,8) ,
55054	 => std_logic_vector(to_unsigned(93,8) ,
55055	 => std_logic_vector(to_unsigned(64,8) ,
55056	 => std_logic_vector(to_unsigned(86,8) ,
55057	 => std_logic_vector(to_unsigned(93,8) ,
55058	 => std_logic_vector(to_unsigned(80,8) ,
55059	 => std_logic_vector(to_unsigned(80,8) ,
55060	 => std_logic_vector(to_unsigned(73,8) ,
55061	 => std_logic_vector(to_unsigned(46,8) ,
55062	 => std_logic_vector(to_unsigned(33,8) ,
55063	 => std_logic_vector(to_unsigned(66,8) ,
55064	 => std_logic_vector(to_unsigned(95,8) ,
55065	 => std_logic_vector(to_unsigned(59,8) ,
55066	 => std_logic_vector(to_unsigned(41,8) ,
55067	 => std_logic_vector(to_unsigned(34,8) ,
55068	 => std_logic_vector(to_unsigned(45,8) ,
55069	 => std_logic_vector(to_unsigned(69,8) ,
55070	 => std_logic_vector(to_unsigned(100,8) ,
55071	 => std_logic_vector(to_unsigned(78,8) ,
55072	 => std_logic_vector(to_unsigned(65,8) ,
55073	 => std_logic_vector(to_unsigned(41,8) ,
55074	 => std_logic_vector(to_unsigned(30,8) ,
55075	 => std_logic_vector(to_unsigned(27,8) ,
55076	 => std_logic_vector(to_unsigned(20,8) ,
55077	 => std_logic_vector(to_unsigned(21,8) ,
55078	 => std_logic_vector(to_unsigned(22,8) ,
55079	 => std_logic_vector(to_unsigned(27,8) ,
55080	 => std_logic_vector(to_unsigned(27,8) ,
55081	 => std_logic_vector(to_unsigned(39,8) ,
55082	 => std_logic_vector(to_unsigned(43,8) ,
55083	 => std_logic_vector(to_unsigned(41,8) ,
55084	 => std_logic_vector(to_unsigned(40,8) ,
55085	 => std_logic_vector(to_unsigned(34,8) ,
55086	 => std_logic_vector(to_unsigned(37,8) ,
55087	 => std_logic_vector(to_unsigned(41,8) ,
55088	 => std_logic_vector(to_unsigned(41,8) ,
55089	 => std_logic_vector(to_unsigned(56,8) ,
55090	 => std_logic_vector(to_unsigned(73,8) ,
55091	 => std_logic_vector(to_unsigned(68,8) ,
55092	 => std_logic_vector(to_unsigned(81,8) ,
55093	 => std_logic_vector(to_unsigned(86,8) ,
55094	 => std_logic_vector(to_unsigned(76,8) ,
55095	 => std_logic_vector(to_unsigned(92,8) ,
55096	 => std_logic_vector(to_unsigned(100,8) ,
55097	 => std_logic_vector(to_unsigned(95,8) ,
55098	 => std_logic_vector(to_unsigned(96,8) ,
55099	 => std_logic_vector(to_unsigned(87,8) ,
55100	 => std_logic_vector(to_unsigned(96,8) ,
55101	 => std_logic_vector(to_unsigned(82,8) ,
55102	 => std_logic_vector(to_unsigned(92,8) ,
55103	 => std_logic_vector(to_unsigned(90,8) ,
55104	 => std_logic_vector(to_unsigned(65,8) ,
55105	 => std_logic_vector(to_unsigned(84,8) ,
55106	 => std_logic_vector(to_unsigned(114,8) ,
55107	 => std_logic_vector(to_unsigned(93,8) ,
55108	 => std_logic_vector(to_unsigned(77,8) ,
55109	 => std_logic_vector(to_unsigned(85,8) ,
55110	 => std_logic_vector(to_unsigned(112,8) ,
55111	 => std_logic_vector(to_unsigned(124,8) ,
55112	 => std_logic_vector(to_unsigned(109,8) ,
55113	 => std_logic_vector(to_unsigned(101,8) ,
55114	 => std_logic_vector(to_unsigned(93,8) ,
55115	 => std_logic_vector(to_unsigned(90,8) ,
55116	 => std_logic_vector(to_unsigned(87,8) ,
55117	 => std_logic_vector(to_unsigned(66,8) ,
55118	 => std_logic_vector(to_unsigned(67,8) ,
55119	 => std_logic_vector(to_unsigned(58,8) ,
55120	 => std_logic_vector(to_unsigned(41,8) ,
55121	 => std_logic_vector(to_unsigned(41,8) ,
55122	 => std_logic_vector(to_unsigned(48,8) ,
55123	 => std_logic_vector(to_unsigned(72,8) ,
55124	 => std_logic_vector(to_unsigned(91,8) ,
55125	 => std_logic_vector(to_unsigned(48,8) ,
55126	 => std_logic_vector(to_unsigned(48,8) ,
55127	 => std_logic_vector(to_unsigned(60,8) ,
55128	 => std_logic_vector(to_unsigned(50,8) ,
55129	 => std_logic_vector(to_unsigned(45,8) ,
55130	 => std_logic_vector(to_unsigned(51,8) ,
55131	 => std_logic_vector(to_unsigned(51,8) ,
55132	 => std_logic_vector(to_unsigned(51,8) ,
55133	 => std_logic_vector(to_unsigned(58,8) ,
55134	 => std_logic_vector(to_unsigned(59,8) ,
55135	 => std_logic_vector(to_unsigned(62,8) ,
55136	 => std_logic_vector(to_unsigned(61,8) ,
55137	 => std_logic_vector(to_unsigned(64,8) ,
55138	 => std_logic_vector(to_unsigned(69,8) ,
55139	 => std_logic_vector(to_unsigned(72,8) ,
55140	 => std_logic_vector(to_unsigned(66,8) ,
55141	 => std_logic_vector(to_unsigned(66,8) ,
55142	 => std_logic_vector(to_unsigned(68,8) ,
55143	 => std_logic_vector(to_unsigned(71,8) ,
55144	 => std_logic_vector(to_unsigned(67,8) ,
55145	 => std_logic_vector(to_unsigned(71,8) ,
55146	 => std_logic_vector(to_unsigned(64,8) ,
55147	 => std_logic_vector(to_unsigned(64,8) ,
55148	 => std_logic_vector(to_unsigned(64,8) ,
55149	 => std_logic_vector(to_unsigned(58,8) ,
55150	 => std_logic_vector(to_unsigned(53,8) ,
55151	 => std_logic_vector(to_unsigned(46,8) ,
55152	 => std_logic_vector(to_unsigned(48,8) ,
55153	 => std_logic_vector(to_unsigned(56,8) ,
55154	 => std_logic_vector(to_unsigned(56,8) ,
55155	 => std_logic_vector(to_unsigned(45,8) ,
55156	 => std_logic_vector(to_unsigned(37,8) ,
55157	 => std_logic_vector(to_unsigned(37,8) ,
55158	 => std_logic_vector(to_unsigned(38,8) ,
55159	 => std_logic_vector(to_unsigned(35,8) ,
55160	 => std_logic_vector(to_unsigned(22,8) ,
55161	 => std_logic_vector(to_unsigned(13,8) ,
55162	 => std_logic_vector(to_unsigned(15,8) ,
55163	 => std_logic_vector(to_unsigned(19,8) ,
55164	 => std_logic_vector(to_unsigned(42,8) ,
55165	 => std_logic_vector(to_unsigned(67,8) ,
55166	 => std_logic_vector(to_unsigned(49,8) ,
55167	 => std_logic_vector(to_unsigned(44,8) ,
55168	 => std_logic_vector(to_unsigned(41,8) ,
55169	 => std_logic_vector(to_unsigned(44,8) ,
55170	 => std_logic_vector(to_unsigned(50,8) ,
55171	 => std_logic_vector(to_unsigned(48,8) ,
55172	 => std_logic_vector(to_unsigned(45,8) ,
55173	 => std_logic_vector(to_unsigned(43,8) ,
55174	 => std_logic_vector(to_unsigned(36,8) ,
55175	 => std_logic_vector(to_unsigned(30,8) ,
55176	 => std_logic_vector(to_unsigned(32,8) ,
55177	 => std_logic_vector(to_unsigned(27,8) ,
55178	 => std_logic_vector(to_unsigned(20,8) ,
55179	 => std_logic_vector(to_unsigned(24,8) ,
55180	 => std_logic_vector(to_unsigned(17,8) ,
55181	 => std_logic_vector(to_unsigned(17,8) ,
55182	 => std_logic_vector(to_unsigned(39,8) ,
55183	 => std_logic_vector(to_unsigned(16,8) ,
55184	 => std_logic_vector(to_unsigned(13,8) ,
55185	 => std_logic_vector(to_unsigned(48,8) ,
55186	 => std_logic_vector(to_unsigned(41,8) ,
55187	 => std_logic_vector(to_unsigned(11,8) ,
55188	 => std_logic_vector(to_unsigned(6,8) ,
55189	 => std_logic_vector(to_unsigned(9,8) ,
55190	 => std_logic_vector(to_unsigned(37,8) ,
55191	 => std_logic_vector(to_unsigned(30,8) ,
55192	 => std_logic_vector(to_unsigned(40,8) ,
55193	 => std_logic_vector(to_unsigned(33,8) ,
55194	 => std_logic_vector(to_unsigned(35,8) ,
55195	 => std_logic_vector(to_unsigned(13,8) ,
55196	 => std_logic_vector(to_unsigned(27,8) ,
55197	 => std_logic_vector(to_unsigned(53,8) ,
55198	 => std_logic_vector(to_unsigned(10,8) ,
55199	 => std_logic_vector(to_unsigned(6,8) ,
55200	 => std_logic_vector(to_unsigned(4,8) ,
55201	 => std_logic_vector(to_unsigned(35,8) ,
55202	 => std_logic_vector(to_unsigned(37,8) ,
55203	 => std_logic_vector(to_unsigned(22,8) ,
55204	 => std_logic_vector(to_unsigned(27,8) ,
55205	 => std_logic_vector(to_unsigned(27,8) ,
55206	 => std_logic_vector(to_unsigned(29,8) ,
55207	 => std_logic_vector(to_unsigned(29,8) ,
55208	 => std_logic_vector(to_unsigned(30,8) ,
55209	 => std_logic_vector(to_unsigned(24,8) ,
55210	 => std_logic_vector(to_unsigned(46,8) ,
55211	 => std_logic_vector(to_unsigned(48,8) ,
55212	 => std_logic_vector(to_unsigned(44,8) ,
55213	 => std_logic_vector(to_unsigned(55,8) ,
55214	 => std_logic_vector(to_unsigned(24,8) ,
55215	 => std_logic_vector(to_unsigned(6,8) ,
55216	 => std_logic_vector(to_unsigned(12,8) ,
55217	 => std_logic_vector(to_unsigned(11,8) ,
55218	 => std_logic_vector(to_unsigned(7,8) ,
55219	 => std_logic_vector(to_unsigned(10,8) ,
55220	 => std_logic_vector(to_unsigned(11,8) ,
55221	 => std_logic_vector(to_unsigned(12,8) ,
55222	 => std_logic_vector(to_unsigned(13,8) ,
55223	 => std_logic_vector(to_unsigned(22,8) ,
55224	 => std_logic_vector(to_unsigned(34,8) ,
55225	 => std_logic_vector(to_unsigned(45,8) ,
55226	 => std_logic_vector(to_unsigned(42,8) ,
55227	 => std_logic_vector(to_unsigned(15,8) ,
55228	 => std_logic_vector(to_unsigned(6,8) ,
55229	 => std_logic_vector(to_unsigned(7,8) ,
55230	 => std_logic_vector(to_unsigned(11,8) ,
55231	 => std_logic_vector(to_unsigned(41,8) ,
55232	 => std_logic_vector(to_unsigned(48,8) ,
55233	 => std_logic_vector(to_unsigned(18,8) ,
55234	 => std_logic_vector(to_unsigned(12,8) ,
55235	 => std_logic_vector(to_unsigned(24,8) ,
55236	 => std_logic_vector(to_unsigned(24,8) ,
55237	 => std_logic_vector(to_unsigned(30,8) ,
55238	 => std_logic_vector(to_unsigned(29,8) ,
55239	 => std_logic_vector(to_unsigned(28,8) ,
55240	 => std_logic_vector(to_unsigned(22,8) ,
55241	 => std_logic_vector(to_unsigned(37,8) ,
55242	 => std_logic_vector(to_unsigned(50,8) ,
55243	 => std_logic_vector(to_unsigned(34,8) ,
55244	 => std_logic_vector(to_unsigned(18,8) ,
55245	 => std_logic_vector(to_unsigned(24,8) ,
55246	 => std_logic_vector(to_unsigned(30,8) ,
55247	 => std_logic_vector(to_unsigned(18,8) ,
55248	 => std_logic_vector(to_unsigned(15,8) ,
55249	 => std_logic_vector(to_unsigned(23,8) ,
55250	 => std_logic_vector(to_unsigned(20,8) ,
55251	 => std_logic_vector(to_unsigned(20,8) ,
55252	 => std_logic_vector(to_unsigned(19,8) ,
55253	 => std_logic_vector(to_unsigned(16,8) ,
55254	 => std_logic_vector(to_unsigned(14,8) ,
55255	 => std_logic_vector(to_unsigned(14,8) ,
55256	 => std_logic_vector(to_unsigned(15,8) ,
55257	 => std_logic_vector(to_unsigned(17,8) ,
55258	 => std_logic_vector(to_unsigned(17,8) ,
55259	 => std_logic_vector(to_unsigned(23,8) ,
55260	 => std_logic_vector(to_unsigned(15,8) ,
55261	 => std_logic_vector(to_unsigned(15,8) ,
55262	 => std_logic_vector(to_unsigned(31,8) ,
55263	 => std_logic_vector(to_unsigned(38,8) ,
55264	 => std_logic_vector(to_unsigned(13,8) ,
55265	 => std_logic_vector(to_unsigned(8,8) ,
55266	 => std_logic_vector(to_unsigned(17,8) ,
55267	 => std_logic_vector(to_unsigned(6,8) ,
55268	 => std_logic_vector(to_unsigned(5,8) ,
55269	 => std_logic_vector(to_unsigned(12,8) ,
55270	 => std_logic_vector(to_unsigned(9,8) ,
55271	 => std_logic_vector(to_unsigned(19,8) ,
55272	 => std_logic_vector(to_unsigned(29,8) ,
55273	 => std_logic_vector(to_unsigned(29,8) ,
55274	 => std_logic_vector(to_unsigned(21,8) ,
55275	 => std_logic_vector(to_unsigned(14,8) ,
55276	 => std_logic_vector(to_unsigned(14,8) ,
55277	 => std_logic_vector(to_unsigned(18,8) ,
55278	 => std_logic_vector(to_unsigned(14,8) ,
55279	 => std_logic_vector(to_unsigned(57,8) ,
55280	 => std_logic_vector(to_unsigned(99,8) ,
55281	 => std_logic_vector(to_unsigned(91,8) ,
55282	 => std_logic_vector(to_unsigned(45,8) ,
55283	 => std_logic_vector(to_unsigned(14,8) ,
55284	 => std_logic_vector(to_unsigned(16,8) ,
55285	 => std_logic_vector(to_unsigned(14,8) ,
55286	 => std_logic_vector(to_unsigned(13,8) ,
55287	 => std_logic_vector(to_unsigned(16,8) ,
55288	 => std_logic_vector(to_unsigned(17,8) ,
55289	 => std_logic_vector(to_unsigned(16,8) ,
55290	 => std_logic_vector(to_unsigned(13,8) ,
55291	 => std_logic_vector(to_unsigned(24,8) ,
55292	 => std_logic_vector(to_unsigned(16,8) ,
55293	 => std_logic_vector(to_unsigned(13,8) ,
55294	 => std_logic_vector(to_unsigned(18,8) ,
55295	 => std_logic_vector(to_unsigned(19,8) ,
55296	 => std_logic_vector(to_unsigned(12,8) ,
55297	 => std_logic_vector(to_unsigned(9,8) ,
55298	 => std_logic_vector(to_unsigned(13,8) ,
55299	 => std_logic_vector(to_unsigned(6,8) ,
55300	 => std_logic_vector(to_unsigned(1,8) ,
55301	 => std_logic_vector(to_unsigned(0,8) ,
55302	 => std_logic_vector(to_unsigned(3,8) ,
55303	 => std_logic_vector(to_unsigned(20,8) ,
55304	 => std_logic_vector(to_unsigned(11,8) ,
55305	 => std_logic_vector(to_unsigned(18,8) ,
55306	 => std_logic_vector(to_unsigned(11,8) ,
55307	 => std_logic_vector(to_unsigned(6,8) ,
55308	 => std_logic_vector(to_unsigned(7,8) ,
55309	 => std_logic_vector(to_unsigned(7,8) ,
55310	 => std_logic_vector(to_unsigned(7,8) ,
55311	 => std_logic_vector(to_unsigned(8,8) ,
55312	 => std_logic_vector(to_unsigned(9,8) ,
55313	 => std_logic_vector(to_unsigned(8,8) ,
55314	 => std_logic_vector(to_unsigned(9,8) ,
55315	 => std_logic_vector(to_unsigned(8,8) ,
55316	 => std_logic_vector(to_unsigned(8,8) ,
55317	 => std_logic_vector(to_unsigned(7,8) ,
55318	 => std_logic_vector(to_unsigned(10,8) ,
55319	 => std_logic_vector(to_unsigned(16,8) ,
55320	 => std_logic_vector(to_unsigned(2,8) ,
55321	 => std_logic_vector(to_unsigned(0,8) ,
55322	 => std_logic_vector(to_unsigned(0,8) ,
55323	 => std_logic_vector(to_unsigned(0,8) ,
55324	 => std_logic_vector(to_unsigned(0,8) ,
55325	 => std_logic_vector(to_unsigned(4,8) ,
55326	 => std_logic_vector(to_unsigned(11,8) ,
55327	 => std_logic_vector(to_unsigned(3,8) ,
55328	 => std_logic_vector(to_unsigned(7,8) ,
55329	 => std_logic_vector(to_unsigned(9,8) ,
55330	 => std_logic_vector(to_unsigned(13,8) ,
55331	 => std_logic_vector(to_unsigned(19,8) ,
55332	 => std_logic_vector(to_unsigned(22,8) ,
55333	 => std_logic_vector(to_unsigned(25,8) ,
55334	 => std_logic_vector(to_unsigned(15,8) ,
55335	 => std_logic_vector(to_unsigned(7,8) ,
55336	 => std_logic_vector(to_unsigned(8,8) ,
55337	 => std_logic_vector(to_unsigned(7,8) ,
55338	 => std_logic_vector(to_unsigned(6,8) ,
55339	 => std_logic_vector(to_unsigned(14,8) ,
55340	 => std_logic_vector(to_unsigned(20,8) ,
55341	 => std_logic_vector(to_unsigned(20,8) ,
55342	 => std_logic_vector(to_unsigned(17,8) ,
55343	 => std_logic_vector(to_unsigned(20,8) ,
55344	 => std_logic_vector(to_unsigned(24,8) ,
55345	 => std_logic_vector(to_unsigned(25,8) ,
55346	 => std_logic_vector(to_unsigned(29,8) ,
55347	 => std_logic_vector(to_unsigned(35,8) ,
55348	 => std_logic_vector(to_unsigned(27,8) ,
55349	 => std_logic_vector(to_unsigned(30,8) ,
55350	 => std_logic_vector(to_unsigned(24,8) ,
55351	 => std_logic_vector(to_unsigned(24,8) ,
55352	 => std_logic_vector(to_unsigned(35,8) ,
55353	 => std_logic_vector(to_unsigned(32,8) ,
55354	 => std_logic_vector(to_unsigned(26,8) ,
55355	 => std_logic_vector(to_unsigned(37,8) ,
55356	 => std_logic_vector(to_unsigned(14,8) ,
55357	 => std_logic_vector(to_unsigned(11,8) ,
55358	 => std_logic_vector(to_unsigned(35,8) ,
55359	 => std_logic_vector(to_unsigned(32,8) ,
55360	 => std_logic_vector(to_unsigned(82,8) ,
55361	 => std_logic_vector(to_unsigned(96,8) ,
55362	 => std_logic_vector(to_unsigned(87,8) ,
55363	 => std_logic_vector(to_unsigned(88,8) ,
55364	 => std_logic_vector(to_unsigned(84,8) ,
55365	 => std_logic_vector(to_unsigned(65,8) ,
55366	 => std_logic_vector(to_unsigned(30,8) ,
55367	 => std_logic_vector(to_unsigned(55,8) ,
55368	 => std_logic_vector(to_unsigned(65,8) ,
55369	 => std_logic_vector(to_unsigned(54,8) ,
55370	 => std_logic_vector(to_unsigned(85,8) ,
55371	 => std_logic_vector(to_unsigned(60,8) ,
55372	 => std_logic_vector(to_unsigned(61,8) ,
55373	 => std_logic_vector(to_unsigned(105,8) ,
55374	 => std_logic_vector(to_unsigned(92,8) ,
55375	 => std_logic_vector(to_unsigned(62,8) ,
55376	 => std_logic_vector(to_unsigned(87,8) ,
55377	 => std_logic_vector(to_unsigned(86,8) ,
55378	 => std_logic_vector(to_unsigned(53,8) ,
55379	 => std_logic_vector(to_unsigned(58,8) ,
55380	 => std_logic_vector(to_unsigned(58,8) ,
55381	 => std_logic_vector(to_unsigned(50,8) ,
55382	 => std_logic_vector(to_unsigned(35,8) ,
55383	 => std_logic_vector(to_unsigned(24,8) ,
55384	 => std_logic_vector(to_unsigned(37,8) ,
55385	 => std_logic_vector(to_unsigned(33,8) ,
55386	 => std_logic_vector(to_unsigned(57,8) ,
55387	 => std_logic_vector(to_unsigned(79,8) ,
55388	 => std_logic_vector(to_unsigned(73,8) ,
55389	 => std_logic_vector(to_unsigned(66,8) ,
55390	 => std_logic_vector(to_unsigned(76,8) ,
55391	 => std_logic_vector(to_unsigned(84,8) ,
55392	 => std_logic_vector(to_unsigned(111,8) ,
55393	 => std_logic_vector(to_unsigned(50,8) ,
55394	 => std_logic_vector(to_unsigned(30,8) ,
55395	 => std_logic_vector(to_unsigned(28,8) ,
55396	 => std_logic_vector(to_unsigned(25,8) ,
55397	 => std_logic_vector(to_unsigned(35,8) ,
55398	 => std_logic_vector(to_unsigned(28,8) ,
55399	 => std_logic_vector(to_unsigned(29,8) ,
55400	 => std_logic_vector(to_unsigned(27,8) ,
55401	 => std_logic_vector(to_unsigned(30,8) ,
55402	 => std_logic_vector(to_unsigned(29,8) ,
55403	 => std_logic_vector(to_unsigned(37,8) ,
55404	 => std_logic_vector(to_unsigned(45,8) ,
55405	 => std_logic_vector(to_unsigned(50,8) ,
55406	 => std_logic_vector(to_unsigned(50,8) ,
55407	 => std_logic_vector(to_unsigned(56,8) ,
55408	 => std_logic_vector(to_unsigned(54,8) ,
55409	 => std_logic_vector(to_unsigned(49,8) ,
55410	 => std_logic_vector(to_unsigned(74,8) ,
55411	 => std_logic_vector(to_unsigned(76,8) ,
55412	 => std_logic_vector(to_unsigned(80,8) ,
55413	 => std_logic_vector(to_unsigned(85,8) ,
55414	 => std_logic_vector(to_unsigned(71,8) ,
55415	 => std_logic_vector(to_unsigned(92,8) ,
55416	 => std_logic_vector(to_unsigned(86,8) ,
55417	 => std_logic_vector(to_unsigned(79,8) ,
55418	 => std_logic_vector(to_unsigned(91,8) ,
55419	 => std_logic_vector(to_unsigned(73,8) ,
55420	 => std_logic_vector(to_unsigned(84,8) ,
55421	 => std_logic_vector(to_unsigned(81,8) ,
55422	 => std_logic_vector(to_unsigned(79,8) ,
55423	 => std_logic_vector(to_unsigned(96,8) ,
55424	 => std_logic_vector(to_unsigned(81,8) ,
55425	 => std_logic_vector(to_unsigned(76,8) ,
55426	 => std_logic_vector(to_unsigned(99,8) ,
55427	 => std_logic_vector(to_unsigned(95,8) ,
55428	 => std_logic_vector(to_unsigned(104,8) ,
55429	 => std_logic_vector(to_unsigned(105,8) ,
55430	 => std_logic_vector(to_unsigned(119,8) ,
55431	 => std_logic_vector(to_unsigned(128,8) ,
55432	 => std_logic_vector(to_unsigned(124,8) ,
55433	 => std_logic_vector(to_unsigned(125,8) ,
55434	 => std_logic_vector(to_unsigned(119,8) ,
55435	 => std_logic_vector(to_unsigned(107,8) ,
55436	 => std_logic_vector(to_unsigned(101,8) ,
55437	 => std_logic_vector(to_unsigned(77,8) ,
55438	 => std_logic_vector(to_unsigned(60,8) ,
55439	 => std_logic_vector(to_unsigned(45,8) ,
55440	 => std_logic_vector(to_unsigned(38,8) ,
55441	 => std_logic_vector(to_unsigned(60,8) ,
55442	 => std_logic_vector(to_unsigned(88,8) ,
55443	 => std_logic_vector(to_unsigned(97,8) ,
55444	 => std_logic_vector(to_unsigned(87,8) ,
55445	 => std_logic_vector(to_unsigned(67,8) ,
55446	 => std_logic_vector(to_unsigned(70,8) ,
55447	 => std_logic_vector(to_unsigned(55,8) ,
55448	 => std_logic_vector(to_unsigned(41,8) ,
55449	 => std_logic_vector(to_unsigned(43,8) ,
55450	 => std_logic_vector(to_unsigned(51,8) ,
55451	 => std_logic_vector(to_unsigned(57,8) ,
55452	 => std_logic_vector(to_unsigned(58,8) ,
55453	 => std_logic_vector(to_unsigned(57,8) ,
55454	 => std_logic_vector(to_unsigned(61,8) ,
55455	 => std_logic_vector(to_unsigned(66,8) ,
55456	 => std_logic_vector(to_unsigned(68,8) ,
55457	 => std_logic_vector(to_unsigned(68,8) ,
55458	 => std_logic_vector(to_unsigned(68,8) ,
55459	 => std_logic_vector(to_unsigned(68,8) ,
55460	 => std_logic_vector(to_unsigned(63,8) ,
55461	 => std_logic_vector(to_unsigned(62,8) ,
55462	 => std_logic_vector(to_unsigned(63,8) ,
55463	 => std_logic_vector(to_unsigned(65,8) ,
55464	 => std_logic_vector(to_unsigned(64,8) ,
55465	 => std_logic_vector(to_unsigned(67,8) ,
55466	 => std_logic_vector(to_unsigned(65,8) ,
55467	 => std_logic_vector(to_unsigned(61,8) ,
55468	 => std_logic_vector(to_unsigned(59,8) ,
55469	 => std_logic_vector(to_unsigned(54,8) ,
55470	 => std_logic_vector(to_unsigned(48,8) ,
55471	 => std_logic_vector(to_unsigned(51,8) ,
55472	 => std_logic_vector(to_unsigned(57,8) ,
55473	 => std_logic_vector(to_unsigned(56,8) ,
55474	 => std_logic_vector(to_unsigned(42,8) ,
55475	 => std_logic_vector(to_unsigned(27,8) ,
55476	 => std_logic_vector(to_unsigned(27,8) ,
55477	 => std_logic_vector(to_unsigned(61,8) ,
55478	 => std_logic_vector(to_unsigned(81,8) ,
55479	 => std_logic_vector(to_unsigned(49,8) ,
55480	 => std_logic_vector(to_unsigned(25,8) ,
55481	 => std_logic_vector(to_unsigned(15,8) ,
55482	 => std_logic_vector(to_unsigned(18,8) ,
55483	 => std_logic_vector(to_unsigned(21,8) ,
55484	 => std_logic_vector(to_unsigned(37,8) ,
55485	 => std_logic_vector(to_unsigned(65,8) ,
55486	 => std_logic_vector(to_unsigned(55,8) ,
55487	 => std_logic_vector(to_unsigned(48,8) ,
55488	 => std_logic_vector(to_unsigned(46,8) ,
55489	 => std_logic_vector(to_unsigned(51,8) ,
55490	 => std_logic_vector(to_unsigned(45,8) ,
55491	 => std_logic_vector(to_unsigned(46,8) ,
55492	 => std_logic_vector(to_unsigned(49,8) ,
55493	 => std_logic_vector(to_unsigned(42,8) ,
55494	 => std_logic_vector(to_unsigned(35,8) ,
55495	 => std_logic_vector(to_unsigned(27,8) ,
55496	 => std_logic_vector(to_unsigned(18,8) ,
55497	 => std_logic_vector(to_unsigned(23,8) ,
55498	 => std_logic_vector(to_unsigned(24,8) ,
55499	 => std_logic_vector(to_unsigned(22,8) ,
55500	 => std_logic_vector(to_unsigned(33,8) ,
55501	 => std_logic_vector(to_unsigned(37,8) ,
55502	 => std_logic_vector(to_unsigned(37,8) ,
55503	 => std_logic_vector(to_unsigned(30,8) ,
55504	 => std_logic_vector(to_unsigned(24,8) ,
55505	 => std_logic_vector(to_unsigned(43,8) ,
55506	 => std_logic_vector(to_unsigned(41,8) ,
55507	 => std_logic_vector(to_unsigned(17,8) ,
55508	 => std_logic_vector(to_unsigned(7,8) ,
55509	 => std_logic_vector(to_unsigned(9,8) ,
55510	 => std_logic_vector(to_unsigned(37,8) ,
55511	 => std_logic_vector(to_unsigned(27,8) ,
55512	 => std_logic_vector(to_unsigned(32,8) ,
55513	 => std_logic_vector(to_unsigned(37,8) ,
55514	 => std_logic_vector(to_unsigned(37,8) ,
55515	 => std_logic_vector(to_unsigned(27,8) ,
55516	 => std_logic_vector(to_unsigned(39,8) ,
55517	 => std_logic_vector(to_unsigned(41,8) ,
55518	 => std_logic_vector(to_unsigned(11,8) ,
55519	 => std_logic_vector(to_unsigned(6,8) ,
55520	 => std_logic_vector(to_unsigned(4,8) ,
55521	 => std_logic_vector(to_unsigned(35,8) ,
55522	 => std_logic_vector(to_unsigned(28,8) ,
55523	 => std_logic_vector(to_unsigned(19,8) ,
55524	 => std_logic_vector(to_unsigned(24,8) ,
55525	 => std_logic_vector(to_unsigned(18,8) ,
55526	 => std_logic_vector(to_unsigned(18,8) ,
55527	 => std_logic_vector(to_unsigned(20,8) ,
55528	 => std_logic_vector(to_unsigned(27,8) ,
55529	 => std_logic_vector(to_unsigned(19,8) ,
55530	 => std_logic_vector(to_unsigned(29,8) ,
55531	 => std_logic_vector(to_unsigned(37,8) ,
55532	 => std_logic_vector(to_unsigned(54,8) ,
55533	 => std_logic_vector(to_unsigned(29,8) ,
55534	 => std_logic_vector(to_unsigned(15,8) ,
55535	 => std_logic_vector(to_unsigned(14,8) ,
55536	 => std_logic_vector(to_unsigned(28,8) ,
55537	 => std_logic_vector(to_unsigned(41,8) ,
55538	 => std_logic_vector(to_unsigned(38,8) ,
55539	 => std_logic_vector(to_unsigned(35,8) ,
55540	 => std_logic_vector(to_unsigned(18,8) ,
55541	 => std_logic_vector(to_unsigned(8,8) ,
55542	 => std_logic_vector(to_unsigned(15,8) ,
55543	 => std_logic_vector(to_unsigned(30,8) ,
55544	 => std_logic_vector(to_unsigned(28,8) ,
55545	 => std_logic_vector(to_unsigned(30,8) ,
55546	 => std_logic_vector(to_unsigned(20,8) ,
55547	 => std_logic_vector(to_unsigned(7,8) ,
55548	 => std_logic_vector(to_unsigned(8,8) ,
55549	 => std_logic_vector(to_unsigned(18,8) ,
55550	 => std_logic_vector(to_unsigned(37,8) ,
55551	 => std_logic_vector(to_unsigned(44,8) ,
55552	 => std_logic_vector(to_unsigned(20,8) ,
55553	 => std_logic_vector(to_unsigned(10,8) ,
55554	 => std_logic_vector(to_unsigned(24,8) ,
55555	 => std_logic_vector(to_unsigned(24,8) ,
55556	 => std_logic_vector(to_unsigned(19,8) ,
55557	 => std_logic_vector(to_unsigned(49,8) ,
55558	 => std_logic_vector(to_unsigned(47,8) ,
55559	 => std_logic_vector(to_unsigned(32,8) ,
55560	 => std_logic_vector(to_unsigned(19,8) ,
55561	 => std_logic_vector(to_unsigned(29,8) ,
55562	 => std_logic_vector(to_unsigned(29,8) ,
55563	 => std_logic_vector(to_unsigned(19,8) ,
55564	 => std_logic_vector(to_unsigned(19,8) ,
55565	 => std_logic_vector(to_unsigned(23,8) ,
55566	 => std_logic_vector(to_unsigned(18,8) ,
55567	 => std_logic_vector(to_unsigned(20,8) ,
55568	 => std_logic_vector(to_unsigned(25,8) ,
55569	 => std_logic_vector(to_unsigned(22,8) ,
55570	 => std_logic_vector(to_unsigned(16,8) ,
55571	 => std_logic_vector(to_unsigned(17,8) ,
55572	 => std_logic_vector(to_unsigned(28,8) ,
55573	 => std_logic_vector(to_unsigned(32,8) ,
55574	 => std_logic_vector(to_unsigned(15,8) ,
55575	 => std_logic_vector(to_unsigned(25,8) ,
55576	 => std_logic_vector(to_unsigned(22,8) ,
55577	 => std_logic_vector(to_unsigned(9,8) ,
55578	 => std_logic_vector(to_unsigned(15,8) ,
55579	 => std_logic_vector(to_unsigned(24,8) ,
55580	 => std_logic_vector(to_unsigned(19,8) ,
55581	 => std_logic_vector(to_unsigned(18,8) ,
55582	 => std_logic_vector(to_unsigned(28,8) ,
55583	 => std_logic_vector(to_unsigned(23,8) ,
55584	 => std_logic_vector(to_unsigned(17,8) ,
55585	 => std_logic_vector(to_unsigned(26,8) ,
55586	 => std_logic_vector(to_unsigned(22,8) ,
55587	 => std_logic_vector(to_unsigned(22,8) ,
55588	 => std_logic_vector(to_unsigned(20,8) ,
55589	 => std_logic_vector(to_unsigned(24,8) ,
55590	 => std_logic_vector(to_unsigned(25,8) ,
55591	 => std_logic_vector(to_unsigned(25,8) ,
55592	 => std_logic_vector(to_unsigned(23,8) ,
55593	 => std_logic_vector(to_unsigned(21,8) ,
55594	 => std_logic_vector(to_unsigned(13,8) ,
55595	 => std_logic_vector(to_unsigned(12,8) ,
55596	 => std_logic_vector(to_unsigned(22,8) ,
55597	 => std_logic_vector(to_unsigned(26,8) ,
55598	 => std_logic_vector(to_unsigned(16,8) ,
55599	 => std_logic_vector(to_unsigned(51,8) ,
55600	 => std_logic_vector(to_unsigned(71,8) ,
55601	 => std_logic_vector(to_unsigned(71,8) ,
55602	 => std_logic_vector(to_unsigned(47,8) ,
55603	 => std_logic_vector(to_unsigned(18,8) ,
55604	 => std_logic_vector(to_unsigned(15,8) ,
55605	 => std_logic_vector(to_unsigned(13,8) ,
55606	 => std_logic_vector(to_unsigned(14,8) ,
55607	 => std_logic_vector(to_unsigned(17,8) ,
55608	 => std_logic_vector(to_unsigned(15,8) ,
55609	 => std_logic_vector(to_unsigned(13,8) ,
55610	 => std_logic_vector(to_unsigned(12,8) ,
55611	 => std_logic_vector(to_unsigned(15,8) ,
55612	 => std_logic_vector(to_unsigned(17,8) ,
55613	 => std_logic_vector(to_unsigned(16,8) ,
55614	 => std_logic_vector(to_unsigned(14,8) ,
55615	 => std_logic_vector(to_unsigned(16,8) ,
55616	 => std_logic_vector(to_unsigned(10,8) ,
55617	 => std_logic_vector(to_unsigned(8,8) ,
55618	 => std_logic_vector(to_unsigned(12,8) ,
55619	 => std_logic_vector(to_unsigned(11,8) ,
55620	 => std_logic_vector(to_unsigned(3,8) ,
55621	 => std_logic_vector(to_unsigned(0,8) ,
55622	 => std_logic_vector(to_unsigned(3,8) ,
55623	 => std_logic_vector(to_unsigned(19,8) ,
55624	 => std_logic_vector(to_unsigned(12,8) ,
55625	 => std_logic_vector(to_unsigned(15,8) ,
55626	 => std_logic_vector(to_unsigned(13,8) ,
55627	 => std_logic_vector(to_unsigned(8,8) ,
55628	 => std_logic_vector(to_unsigned(8,8) ,
55629	 => std_logic_vector(to_unsigned(9,8) ,
55630	 => std_logic_vector(to_unsigned(12,8) ,
55631	 => std_logic_vector(to_unsigned(11,8) ,
55632	 => std_logic_vector(to_unsigned(8,8) ,
55633	 => std_logic_vector(to_unsigned(8,8) ,
55634	 => std_logic_vector(to_unsigned(7,8) ,
55635	 => std_logic_vector(to_unsigned(8,8) ,
55636	 => std_logic_vector(to_unsigned(8,8) ,
55637	 => std_logic_vector(to_unsigned(7,8) ,
55638	 => std_logic_vector(to_unsigned(5,8) ,
55639	 => std_logic_vector(to_unsigned(12,8) ,
55640	 => std_logic_vector(to_unsigned(6,8) ,
55641	 => std_logic_vector(to_unsigned(0,8) ,
55642	 => std_logic_vector(to_unsigned(0,8) ,
55643	 => std_logic_vector(to_unsigned(0,8) ,
55644	 => std_logic_vector(to_unsigned(0,8) ,
55645	 => std_logic_vector(to_unsigned(2,8) ,
55646	 => std_logic_vector(to_unsigned(13,8) ,
55647	 => std_logic_vector(to_unsigned(12,8) ,
55648	 => std_logic_vector(to_unsigned(23,8) ,
55649	 => std_logic_vector(to_unsigned(19,8) ,
55650	 => std_logic_vector(to_unsigned(12,8) ,
55651	 => std_logic_vector(to_unsigned(18,8) ,
55652	 => std_logic_vector(to_unsigned(17,8) ,
55653	 => std_logic_vector(to_unsigned(17,8) ,
55654	 => std_logic_vector(to_unsigned(15,8) ,
55655	 => std_logic_vector(to_unsigned(10,8) ,
55656	 => std_logic_vector(to_unsigned(10,8) ,
55657	 => std_logic_vector(to_unsigned(7,8) ,
55658	 => std_logic_vector(to_unsigned(8,8) ,
55659	 => std_logic_vector(to_unsigned(17,8) ,
55660	 => std_logic_vector(to_unsigned(18,8) ,
55661	 => std_logic_vector(to_unsigned(16,8) ,
55662	 => std_logic_vector(to_unsigned(13,8) ,
55663	 => std_logic_vector(to_unsigned(10,8) ,
55664	 => std_logic_vector(to_unsigned(12,8) ,
55665	 => std_logic_vector(to_unsigned(15,8) ,
55666	 => std_logic_vector(to_unsigned(20,8) ,
55667	 => std_logic_vector(to_unsigned(30,8) ,
55668	 => std_logic_vector(to_unsigned(11,8) ,
55669	 => std_logic_vector(to_unsigned(43,8) ,
55670	 => std_logic_vector(to_unsigned(22,8) ,
55671	 => std_logic_vector(to_unsigned(24,8) ,
55672	 => std_logic_vector(to_unsigned(33,8) ,
55673	 => std_logic_vector(to_unsigned(24,8) ,
55674	 => std_logic_vector(to_unsigned(27,8) ,
55675	 => std_logic_vector(to_unsigned(32,8) ,
55676	 => std_logic_vector(to_unsigned(21,8) ,
55677	 => std_logic_vector(to_unsigned(35,8) ,
55678	 => std_logic_vector(to_unsigned(53,8) ,
55679	 => std_logic_vector(to_unsigned(52,8) ,
55680	 => std_logic_vector(to_unsigned(104,8) ,
55681	 => std_logic_vector(to_unsigned(96,8) ,
55682	 => std_logic_vector(to_unsigned(95,8) ,
55683	 => std_logic_vector(to_unsigned(96,8) ,
55684	 => std_logic_vector(to_unsigned(69,8) ,
55685	 => std_logic_vector(to_unsigned(37,8) ,
55686	 => std_logic_vector(to_unsigned(32,8) ,
55687	 => std_logic_vector(to_unsigned(50,8) ,
55688	 => std_logic_vector(to_unsigned(57,8) ,
55689	 => std_logic_vector(to_unsigned(66,8) ,
55690	 => std_logic_vector(to_unsigned(81,8) ,
55691	 => std_logic_vector(to_unsigned(55,8) ,
55692	 => std_logic_vector(to_unsigned(64,8) ,
55693	 => std_logic_vector(to_unsigned(99,8) ,
55694	 => std_logic_vector(to_unsigned(95,8) ,
55695	 => std_logic_vector(to_unsigned(111,8) ,
55696	 => std_logic_vector(to_unsigned(108,8) ,
55697	 => std_logic_vector(to_unsigned(74,8) ,
55698	 => std_logic_vector(to_unsigned(51,8) ,
55699	 => std_logic_vector(to_unsigned(53,8) ,
55700	 => std_logic_vector(to_unsigned(71,8) ,
55701	 => std_logic_vector(to_unsigned(49,8) ,
55702	 => std_logic_vector(to_unsigned(31,8) ,
55703	 => std_logic_vector(to_unsigned(37,8) ,
55704	 => std_logic_vector(to_unsigned(69,8) ,
55705	 => std_logic_vector(to_unsigned(69,8) ,
55706	 => std_logic_vector(to_unsigned(77,8) ,
55707	 => std_logic_vector(to_unsigned(80,8) ,
55708	 => std_logic_vector(to_unsigned(72,8) ,
55709	 => std_logic_vector(to_unsigned(91,8) ,
55710	 => std_logic_vector(to_unsigned(97,8) ,
55711	 => std_logic_vector(to_unsigned(96,8) ,
55712	 => std_logic_vector(to_unsigned(100,8) ,
55713	 => std_logic_vector(to_unsigned(55,8) ,
55714	 => std_logic_vector(to_unsigned(23,8) ,
55715	 => std_logic_vector(to_unsigned(28,8) ,
55716	 => std_logic_vector(to_unsigned(20,8) ,
55717	 => std_logic_vector(to_unsigned(22,8) ,
55718	 => std_logic_vector(to_unsigned(30,8) ,
55719	 => std_logic_vector(to_unsigned(35,8) ,
55720	 => std_logic_vector(to_unsigned(27,8) ,
55721	 => std_logic_vector(to_unsigned(30,8) ,
55722	 => std_logic_vector(to_unsigned(31,8) ,
55723	 => std_logic_vector(to_unsigned(35,8) ,
55724	 => std_logic_vector(to_unsigned(35,8) ,
55725	 => std_logic_vector(to_unsigned(32,8) ,
55726	 => std_logic_vector(to_unsigned(36,8) ,
55727	 => std_logic_vector(to_unsigned(44,8) ,
55728	 => std_logic_vector(to_unsigned(49,8) ,
55729	 => std_logic_vector(to_unsigned(47,8) ,
55730	 => std_logic_vector(to_unsigned(64,8) ,
55731	 => std_logic_vector(to_unsigned(56,8) ,
55732	 => std_logic_vector(to_unsigned(59,8) ,
55733	 => std_logic_vector(to_unsigned(79,8) ,
55734	 => std_logic_vector(to_unsigned(81,8) ,
55735	 => std_logic_vector(to_unsigned(87,8) ,
55736	 => std_logic_vector(to_unsigned(73,8) ,
55737	 => std_logic_vector(to_unsigned(70,8) ,
55738	 => std_logic_vector(to_unsigned(79,8) ,
55739	 => std_logic_vector(to_unsigned(70,8) ,
55740	 => std_logic_vector(to_unsigned(80,8) ,
55741	 => std_logic_vector(to_unsigned(56,8) ,
55742	 => std_logic_vector(to_unsigned(58,8) ,
55743	 => std_logic_vector(to_unsigned(92,8) ,
55744	 => std_logic_vector(to_unsigned(86,8) ,
55745	 => std_logic_vector(to_unsigned(114,8) ,
55746	 => std_logic_vector(to_unsigned(144,8) ,
55747	 => std_logic_vector(to_unsigned(99,8) ,
55748	 => std_logic_vector(to_unsigned(91,8) ,
55749	 => std_logic_vector(to_unsigned(107,8) ,
55750	 => std_logic_vector(to_unsigned(103,8) ,
55751	 => std_logic_vector(to_unsigned(99,8) ,
55752	 => std_logic_vector(to_unsigned(104,8) ,
55753	 => std_logic_vector(to_unsigned(112,8) ,
55754	 => std_logic_vector(to_unsigned(116,8) ,
55755	 => std_logic_vector(to_unsigned(111,8) ,
55756	 => std_logic_vector(to_unsigned(108,8) ,
55757	 => std_logic_vector(to_unsigned(66,8) ,
55758	 => std_logic_vector(to_unsigned(45,8) ,
55759	 => std_logic_vector(to_unsigned(60,8) ,
55760	 => std_logic_vector(to_unsigned(87,8) ,
55761	 => std_logic_vector(to_unsigned(104,8) ,
55762	 => std_logic_vector(to_unsigned(103,8) ,
55763	 => std_logic_vector(to_unsigned(95,8) ,
55764	 => std_logic_vector(to_unsigned(80,8) ,
55765	 => std_logic_vector(to_unsigned(72,8) ,
55766	 => std_logic_vector(to_unsigned(63,8) ,
55767	 => std_logic_vector(to_unsigned(39,8) ,
55768	 => std_logic_vector(to_unsigned(37,8) ,
55769	 => std_logic_vector(to_unsigned(43,8) ,
55770	 => std_logic_vector(to_unsigned(49,8) ,
55771	 => std_logic_vector(to_unsigned(57,8) ,
55772	 => std_logic_vector(to_unsigned(59,8) ,
55773	 => std_logic_vector(to_unsigned(54,8) ,
55774	 => std_logic_vector(to_unsigned(61,8) ,
55775	 => std_logic_vector(to_unsigned(62,8) ,
55776	 => std_logic_vector(to_unsigned(63,8) ,
55777	 => std_logic_vector(to_unsigned(66,8) ,
55778	 => std_logic_vector(to_unsigned(65,8) ,
55779	 => std_logic_vector(to_unsigned(60,8) ,
55780	 => std_logic_vector(to_unsigned(62,8) ,
55781	 => std_logic_vector(to_unsigned(59,8) ,
55782	 => std_logic_vector(to_unsigned(60,8) ,
55783	 => std_logic_vector(to_unsigned(59,8) ,
55784	 => std_logic_vector(to_unsigned(55,8) ,
55785	 => std_logic_vector(to_unsigned(61,8) ,
55786	 => std_logic_vector(to_unsigned(62,8) ,
55787	 => std_logic_vector(to_unsigned(58,8) ,
55788	 => std_logic_vector(to_unsigned(57,8) ,
55789	 => std_logic_vector(to_unsigned(52,8) ,
55790	 => std_logic_vector(to_unsigned(41,8) ,
55791	 => std_logic_vector(to_unsigned(45,8) ,
55792	 => std_logic_vector(to_unsigned(42,8) ,
55793	 => std_logic_vector(to_unsigned(34,8) ,
55794	 => std_logic_vector(to_unsigned(32,8) ,
55795	 => std_logic_vector(to_unsigned(35,8) ,
55796	 => std_logic_vector(to_unsigned(66,8) ,
55797	 => std_logic_vector(to_unsigned(109,8) ,
55798	 => std_logic_vector(to_unsigned(99,8) ,
55799	 => std_logic_vector(to_unsigned(53,8) ,
55800	 => std_logic_vector(to_unsigned(25,8) ,
55801	 => std_logic_vector(to_unsigned(12,8) ,
55802	 => std_logic_vector(to_unsigned(16,8) ,
55803	 => std_logic_vector(to_unsigned(19,8) ,
55804	 => std_logic_vector(to_unsigned(27,8) ,
55805	 => std_logic_vector(to_unsigned(52,8) ,
55806	 => std_logic_vector(to_unsigned(47,8) ,
55807	 => std_logic_vector(to_unsigned(49,8) ,
55808	 => std_logic_vector(to_unsigned(50,8) ,
55809	 => std_logic_vector(to_unsigned(42,8) ,
55810	 => std_logic_vector(to_unsigned(40,8) ,
55811	 => std_logic_vector(to_unsigned(46,8) ,
55812	 => std_logic_vector(to_unsigned(51,8) ,
55813	 => std_logic_vector(to_unsigned(40,8) ,
55814	 => std_logic_vector(to_unsigned(35,8) ,
55815	 => std_logic_vector(to_unsigned(26,8) ,
55816	 => std_logic_vector(to_unsigned(16,8) ,
55817	 => std_logic_vector(to_unsigned(18,8) ,
55818	 => std_logic_vector(to_unsigned(22,8) ,
55819	 => std_logic_vector(to_unsigned(29,8) ,
55820	 => std_logic_vector(to_unsigned(37,8) ,
55821	 => std_logic_vector(to_unsigned(39,8) ,
55822	 => std_logic_vector(to_unsigned(36,8) ,
55823	 => std_logic_vector(to_unsigned(49,8) ,
55824	 => std_logic_vector(to_unsigned(57,8) ,
55825	 => std_logic_vector(to_unsigned(35,8) ,
55826	 => std_logic_vector(to_unsigned(36,8) ,
55827	 => std_logic_vector(to_unsigned(32,8) ,
55828	 => std_logic_vector(to_unsigned(24,8) ,
55829	 => std_logic_vector(to_unsigned(27,8) ,
55830	 => std_logic_vector(to_unsigned(31,8) ,
55831	 => std_logic_vector(to_unsigned(24,8) ,
55832	 => std_logic_vector(to_unsigned(32,8) ,
55833	 => std_logic_vector(to_unsigned(32,8) ,
55834	 => std_logic_vector(to_unsigned(29,8) ,
55835	 => std_logic_vector(to_unsigned(12,8) ,
55836	 => std_logic_vector(to_unsigned(26,8) ,
55837	 => std_logic_vector(to_unsigned(30,8) ,
55838	 => std_logic_vector(to_unsigned(6,8) ,
55839	 => std_logic_vector(to_unsigned(5,8) ,
55840	 => std_logic_vector(to_unsigned(3,8) ,
55841	 => std_logic_vector(to_unsigned(25,8) ,
55842	 => std_logic_vector(to_unsigned(45,8) ,
55843	 => std_logic_vector(to_unsigned(26,8) ,
55844	 => std_logic_vector(to_unsigned(22,8) ,
55845	 => std_logic_vector(to_unsigned(27,8) ,
55846	 => std_logic_vector(to_unsigned(33,8) ,
55847	 => std_logic_vector(to_unsigned(15,8) ,
55848	 => std_logic_vector(to_unsigned(23,8) ,
55849	 => std_logic_vector(to_unsigned(30,8) ,
55850	 => std_logic_vector(to_unsigned(22,8) ,
55851	 => std_logic_vector(to_unsigned(14,8) ,
55852	 => std_logic_vector(to_unsigned(17,8) ,
55853	 => std_logic_vector(to_unsigned(13,8) ,
55854	 => std_logic_vector(to_unsigned(13,8) ,
55855	 => std_logic_vector(to_unsigned(16,8) ,
55856	 => std_logic_vector(to_unsigned(26,8) ,
55857	 => std_logic_vector(to_unsigned(52,8) ,
55858	 => std_logic_vector(to_unsigned(51,8) ,
55859	 => std_logic_vector(to_unsigned(35,8) ,
55860	 => std_logic_vector(to_unsigned(33,8) ,
55861	 => std_logic_vector(to_unsigned(25,8) ,
55862	 => std_logic_vector(to_unsigned(25,8) ,
55863	 => std_logic_vector(to_unsigned(22,8) ,
55864	 => std_logic_vector(to_unsigned(9,8) ,
55865	 => std_logic_vector(to_unsigned(12,8) ,
55866	 => std_logic_vector(to_unsigned(12,8) ,
55867	 => std_logic_vector(to_unsigned(9,8) ,
55868	 => std_logic_vector(to_unsigned(29,8) ,
55869	 => std_logic_vector(to_unsigned(55,8) ,
55870	 => std_logic_vector(to_unsigned(48,8) ,
55871	 => std_logic_vector(to_unsigned(19,8) ,
55872	 => std_logic_vector(to_unsigned(12,8) ,
55873	 => std_logic_vector(to_unsigned(24,8) ,
55874	 => std_logic_vector(to_unsigned(21,8) ,
55875	 => std_logic_vector(to_unsigned(19,8) ,
55876	 => std_logic_vector(to_unsigned(23,8) ,
55877	 => std_logic_vector(to_unsigned(59,8) ,
55878	 => std_logic_vector(to_unsigned(63,8) ,
55879	 => std_logic_vector(to_unsigned(40,8) ,
55880	 => std_logic_vector(to_unsigned(18,8) ,
55881	 => std_logic_vector(to_unsigned(45,8) ,
55882	 => std_logic_vector(to_unsigned(59,8) ,
55883	 => std_logic_vector(to_unsigned(37,8) ,
55884	 => std_logic_vector(to_unsigned(17,8) ,
55885	 => std_logic_vector(to_unsigned(24,8) ,
55886	 => std_logic_vector(to_unsigned(16,8) ,
55887	 => std_logic_vector(to_unsigned(14,8) ,
55888	 => std_logic_vector(to_unsigned(18,8) ,
55889	 => std_logic_vector(to_unsigned(20,8) ,
55890	 => std_logic_vector(to_unsigned(18,8) ,
55891	 => std_logic_vector(to_unsigned(16,8) ,
55892	 => std_logic_vector(to_unsigned(17,8) ,
55893	 => std_logic_vector(to_unsigned(20,8) ,
55894	 => std_logic_vector(to_unsigned(16,8) ,
55895	 => std_logic_vector(to_unsigned(24,8) ,
55896	 => std_logic_vector(to_unsigned(20,8) ,
55897	 => std_logic_vector(to_unsigned(11,8) ,
55898	 => std_logic_vector(to_unsigned(17,8) ,
55899	 => std_logic_vector(to_unsigned(34,8) ,
55900	 => std_logic_vector(to_unsigned(18,8) ,
55901	 => std_logic_vector(to_unsigned(21,8) ,
55902	 => std_logic_vector(to_unsigned(28,8) ,
55903	 => std_logic_vector(to_unsigned(18,8) ,
55904	 => std_logic_vector(to_unsigned(12,8) ,
55905	 => std_logic_vector(to_unsigned(16,8) ,
55906	 => std_logic_vector(to_unsigned(15,8) ,
55907	 => std_logic_vector(to_unsigned(27,8) ,
55908	 => std_logic_vector(to_unsigned(40,8) ,
55909	 => std_logic_vector(to_unsigned(37,8) ,
55910	 => std_logic_vector(to_unsigned(43,8) ,
55911	 => std_logic_vector(to_unsigned(41,8) ,
55912	 => std_logic_vector(to_unsigned(20,8) ,
55913	 => std_logic_vector(to_unsigned(12,8) ,
55914	 => std_logic_vector(to_unsigned(10,8) ,
55915	 => std_logic_vector(to_unsigned(16,8) ,
55916	 => std_logic_vector(to_unsigned(22,8) ,
55917	 => std_logic_vector(to_unsigned(17,8) ,
55918	 => std_logic_vector(to_unsigned(15,8) ,
55919	 => std_logic_vector(to_unsigned(61,8) ,
55920	 => std_logic_vector(to_unsigned(73,8) ,
55921	 => std_logic_vector(to_unsigned(76,8) ,
55922	 => std_logic_vector(to_unsigned(40,8) ,
55923	 => std_logic_vector(to_unsigned(10,8) ,
55924	 => std_logic_vector(to_unsigned(14,8) ,
55925	 => std_logic_vector(to_unsigned(13,8) ,
55926	 => std_logic_vector(to_unsigned(12,8) ,
55927	 => std_logic_vector(to_unsigned(13,8) ,
55928	 => std_logic_vector(to_unsigned(13,8) ,
55929	 => std_logic_vector(to_unsigned(12,8) ,
55930	 => std_logic_vector(to_unsigned(10,8) ,
55931	 => std_logic_vector(to_unsigned(12,8) ,
55932	 => std_logic_vector(to_unsigned(18,8) ,
55933	 => std_logic_vector(to_unsigned(22,8) ,
55934	 => std_logic_vector(to_unsigned(12,8) ,
55935	 => std_logic_vector(to_unsigned(13,8) ,
55936	 => std_logic_vector(to_unsigned(14,8) ,
55937	 => std_logic_vector(to_unsigned(13,8) ,
55938	 => std_logic_vector(to_unsigned(13,8) ,
55939	 => std_logic_vector(to_unsigned(24,8) ,
55940	 => std_logic_vector(to_unsigned(8,8) ,
55941	 => std_logic_vector(to_unsigned(0,8) ,
55942	 => std_logic_vector(to_unsigned(1,8) ,
55943	 => std_logic_vector(to_unsigned(12,8) ,
55944	 => std_logic_vector(to_unsigned(15,8) ,
55945	 => std_logic_vector(to_unsigned(12,8) ,
55946	 => std_logic_vector(to_unsigned(14,8) ,
55947	 => std_logic_vector(to_unsigned(16,8) ,
55948	 => std_logic_vector(to_unsigned(16,8) ,
55949	 => std_logic_vector(to_unsigned(12,8) ,
55950	 => std_logic_vector(to_unsigned(13,8) ,
55951	 => std_logic_vector(to_unsigned(12,8) ,
55952	 => std_logic_vector(to_unsigned(8,8) ,
55953	 => std_logic_vector(to_unsigned(7,8) ,
55954	 => std_logic_vector(to_unsigned(9,8) ,
55955	 => std_logic_vector(to_unsigned(7,8) ,
55956	 => std_logic_vector(to_unsigned(8,8) ,
55957	 => std_logic_vector(to_unsigned(10,8) ,
55958	 => std_logic_vector(to_unsigned(7,8) ,
55959	 => std_logic_vector(to_unsigned(11,8) ,
55960	 => std_logic_vector(to_unsigned(7,8) ,
55961	 => std_logic_vector(to_unsigned(0,8) ,
55962	 => std_logic_vector(to_unsigned(0,8) ,
55963	 => std_logic_vector(to_unsigned(0,8) ,
55964	 => std_logic_vector(to_unsigned(0,8) ,
55965	 => std_logic_vector(to_unsigned(1,8) ,
55966	 => std_logic_vector(to_unsigned(7,8) ,
55967	 => std_logic_vector(to_unsigned(10,8) ,
55968	 => std_logic_vector(to_unsigned(10,8) ,
55969	 => std_logic_vector(to_unsigned(18,8) ,
55970	 => std_logic_vector(to_unsigned(14,8) ,
55971	 => std_logic_vector(to_unsigned(17,8) ,
55972	 => std_logic_vector(to_unsigned(17,8) ,
55973	 => std_logic_vector(to_unsigned(17,8) ,
55974	 => std_logic_vector(to_unsigned(16,8) ,
55975	 => std_logic_vector(to_unsigned(17,8) ,
55976	 => std_logic_vector(to_unsigned(16,8) ,
55977	 => std_logic_vector(to_unsigned(8,8) ,
55978	 => std_logic_vector(to_unsigned(9,8) ,
55979	 => std_logic_vector(to_unsigned(17,8) ,
55980	 => std_logic_vector(to_unsigned(25,8) ,
55981	 => std_logic_vector(to_unsigned(25,8) ,
55982	 => std_logic_vector(to_unsigned(25,8) ,
55983	 => std_logic_vector(to_unsigned(19,8) ,
55984	 => std_logic_vector(to_unsigned(25,8) ,
55985	 => std_logic_vector(to_unsigned(25,8) ,
55986	 => std_logic_vector(to_unsigned(24,8) ,
55987	 => std_logic_vector(to_unsigned(23,8) ,
55988	 => std_logic_vector(to_unsigned(15,8) ,
55989	 => std_logic_vector(to_unsigned(40,8) ,
55990	 => std_logic_vector(to_unsigned(32,8) ,
55991	 => std_logic_vector(to_unsigned(51,8) ,
55992	 => std_logic_vector(to_unsigned(35,8) ,
55993	 => std_logic_vector(to_unsigned(20,8) ,
55994	 => std_logic_vector(to_unsigned(19,8) ,
55995	 => std_logic_vector(to_unsigned(14,8) ,
55996	 => std_logic_vector(to_unsigned(2,8) ,
55997	 => std_logic_vector(to_unsigned(4,8) ,
55998	 => std_logic_vector(to_unsigned(17,8) ,
55999	 => std_logic_vector(to_unsigned(26,8) ,
56000	 => std_logic_vector(to_unsigned(105,8) ,
56001	 => std_logic_vector(to_unsigned(95,8) ,
56002	 => std_logic_vector(to_unsigned(69,8) ,
56003	 => std_logic_vector(to_unsigned(81,8) ,
56004	 => std_logic_vector(to_unsigned(80,8) ,
56005	 => std_logic_vector(to_unsigned(45,8) ,
56006	 => std_logic_vector(to_unsigned(29,8) ,
56007	 => std_logic_vector(to_unsigned(37,8) ,
56008	 => std_logic_vector(to_unsigned(56,8) ,
56009	 => std_logic_vector(to_unsigned(51,8) ,
56010	 => std_logic_vector(to_unsigned(76,8) ,
56011	 => std_logic_vector(to_unsigned(77,8) ,
56012	 => std_logic_vector(to_unsigned(73,8) ,
56013	 => std_logic_vector(to_unsigned(95,8) ,
56014	 => std_logic_vector(to_unsigned(97,8) ,
56015	 => std_logic_vector(to_unsigned(70,8) ,
56016	 => std_logic_vector(to_unsigned(73,8) ,
56017	 => std_logic_vector(to_unsigned(96,8) ,
56018	 => std_logic_vector(to_unsigned(82,8) ,
56019	 => std_logic_vector(to_unsigned(73,8) ,
56020	 => std_logic_vector(to_unsigned(71,8) ,
56021	 => std_logic_vector(to_unsigned(42,8) ,
56022	 => std_logic_vector(to_unsigned(30,8) ,
56023	 => std_logic_vector(to_unsigned(35,8) ,
56024	 => std_logic_vector(to_unsigned(67,8) ,
56025	 => std_logic_vector(to_unsigned(69,8) ,
56026	 => std_logic_vector(to_unsigned(57,8) ,
56027	 => std_logic_vector(to_unsigned(96,8) ,
56028	 => std_logic_vector(to_unsigned(115,8) ,
56029	 => std_logic_vector(to_unsigned(124,8) ,
56030	 => std_logic_vector(to_unsigned(115,8) ,
56031	 => std_logic_vector(to_unsigned(91,8) ,
56032	 => std_logic_vector(to_unsigned(81,8) ,
56033	 => std_logic_vector(to_unsigned(59,8) ,
56034	 => std_logic_vector(to_unsigned(24,8) ,
56035	 => std_logic_vector(to_unsigned(26,8) ,
56036	 => std_logic_vector(to_unsigned(23,8) ,
56037	 => std_logic_vector(to_unsigned(27,8) ,
56038	 => std_logic_vector(to_unsigned(22,8) ,
56039	 => std_logic_vector(to_unsigned(21,8) ,
56040	 => std_logic_vector(to_unsigned(20,8) ,
56041	 => std_logic_vector(to_unsigned(36,8) ,
56042	 => std_logic_vector(to_unsigned(45,8) ,
56043	 => std_logic_vector(to_unsigned(41,8) ,
56044	 => std_logic_vector(to_unsigned(50,8) ,
56045	 => std_logic_vector(to_unsigned(45,8) ,
56046	 => std_logic_vector(to_unsigned(37,8) ,
56047	 => std_logic_vector(to_unsigned(39,8) ,
56048	 => std_logic_vector(to_unsigned(41,8) ,
56049	 => std_logic_vector(to_unsigned(42,8) ,
56050	 => std_logic_vector(to_unsigned(61,8) ,
56051	 => std_logic_vector(to_unsigned(59,8) ,
56052	 => std_logic_vector(to_unsigned(61,8) ,
56053	 => std_logic_vector(to_unsigned(70,8) ,
56054	 => std_logic_vector(to_unsigned(53,8) ,
56055	 => std_logic_vector(to_unsigned(72,8) ,
56056	 => std_logic_vector(to_unsigned(67,8) ,
56057	 => std_logic_vector(to_unsigned(44,8) ,
56058	 => std_logic_vector(to_unsigned(55,8) ,
56059	 => std_logic_vector(to_unsigned(54,8) ,
56060	 => std_logic_vector(to_unsigned(59,8) ,
56061	 => std_logic_vector(to_unsigned(59,8) ,
56062	 => std_logic_vector(to_unsigned(60,8) ,
56063	 => std_logic_vector(to_unsigned(81,8) ,
56064	 => std_logic_vector(to_unsigned(76,8) ,
56065	 => std_logic_vector(to_unsigned(114,8) ,
56066	 => std_logic_vector(to_unsigned(138,8) ,
56067	 => std_logic_vector(to_unsigned(85,8) ,
56068	 => std_logic_vector(to_unsigned(77,8) ,
56069	 => std_logic_vector(to_unsigned(112,8) ,
56070	 => std_logic_vector(to_unsigned(107,8) ,
56071	 => std_logic_vector(to_unsigned(96,8) ,
56072	 => std_logic_vector(to_unsigned(109,8) ,
56073	 => std_logic_vector(to_unsigned(115,8) ,
56074	 => std_logic_vector(to_unsigned(104,8) ,
56075	 => std_logic_vector(to_unsigned(100,8) ,
56076	 => std_logic_vector(to_unsigned(104,8) ,
56077	 => std_logic_vector(to_unsigned(78,8) ,
56078	 => std_logic_vector(to_unsigned(72,8) ,
56079	 => std_logic_vector(to_unsigned(112,8) ,
56080	 => std_logic_vector(to_unsigned(128,8) ,
56081	 => std_logic_vector(to_unsigned(111,8) ,
56082	 => std_logic_vector(to_unsigned(84,8) ,
56083	 => std_logic_vector(to_unsigned(96,8) ,
56084	 => std_logic_vector(to_unsigned(92,8) ,
56085	 => std_logic_vector(to_unsigned(50,8) ,
56086	 => std_logic_vector(to_unsigned(41,8) ,
56087	 => std_logic_vector(to_unsigned(39,8) ,
56088	 => std_logic_vector(to_unsigned(39,8) ,
56089	 => std_logic_vector(to_unsigned(41,8) ,
56090	 => std_logic_vector(to_unsigned(42,8) ,
56091	 => std_logic_vector(to_unsigned(45,8) ,
56092	 => std_logic_vector(to_unsigned(50,8) ,
56093	 => std_logic_vector(to_unsigned(54,8) ,
56094	 => std_logic_vector(to_unsigned(63,8) ,
56095	 => std_logic_vector(to_unsigned(61,8) ,
56096	 => std_logic_vector(to_unsigned(55,8) ,
56097	 => std_logic_vector(to_unsigned(61,8) ,
56098	 => std_logic_vector(to_unsigned(61,8) ,
56099	 => std_logic_vector(to_unsigned(63,8) ,
56100	 => std_logic_vector(to_unsigned(64,8) ,
56101	 => std_logic_vector(to_unsigned(59,8) ,
56102	 => std_logic_vector(to_unsigned(61,8) ,
56103	 => std_logic_vector(to_unsigned(62,8) ,
56104	 => std_logic_vector(to_unsigned(56,8) ,
56105	 => std_logic_vector(to_unsigned(59,8) ,
56106	 => std_logic_vector(to_unsigned(65,8) ,
56107	 => std_logic_vector(to_unsigned(59,8) ,
56108	 => std_logic_vector(to_unsigned(55,8) ,
56109	 => std_logic_vector(to_unsigned(45,8) ,
56110	 => std_logic_vector(to_unsigned(46,8) ,
56111	 => std_logic_vector(to_unsigned(54,8) ,
56112	 => std_logic_vector(to_unsigned(45,8) ,
56113	 => std_logic_vector(to_unsigned(32,8) ,
56114	 => std_logic_vector(to_unsigned(51,8) ,
56115	 => std_logic_vector(to_unsigned(104,8) ,
56116	 => std_logic_vector(to_unsigned(115,8) ,
56117	 => std_logic_vector(to_unsigned(72,8) ,
56118	 => std_logic_vector(to_unsigned(67,8) ,
56119	 => std_logic_vector(to_unsigned(57,8) ,
56120	 => std_logic_vector(to_unsigned(27,8) ,
56121	 => std_logic_vector(to_unsigned(12,8) ,
56122	 => std_logic_vector(to_unsigned(12,8) ,
56123	 => std_logic_vector(to_unsigned(14,8) ,
56124	 => std_logic_vector(to_unsigned(25,8) ,
56125	 => std_logic_vector(to_unsigned(41,8) ,
56126	 => std_logic_vector(to_unsigned(42,8) ,
56127	 => std_logic_vector(to_unsigned(45,8) ,
56128	 => std_logic_vector(to_unsigned(41,8) ,
56129	 => std_logic_vector(to_unsigned(41,8) ,
56130	 => std_logic_vector(to_unsigned(47,8) ,
56131	 => std_logic_vector(to_unsigned(50,8) ,
56132	 => std_logic_vector(to_unsigned(48,8) ,
56133	 => std_logic_vector(to_unsigned(37,8) ,
56134	 => std_logic_vector(to_unsigned(35,8) ,
56135	 => std_logic_vector(to_unsigned(35,8) ,
56136	 => std_logic_vector(to_unsigned(30,8) ,
56137	 => std_logic_vector(to_unsigned(27,8) ,
56138	 => std_logic_vector(to_unsigned(33,8) ,
56139	 => std_logic_vector(to_unsigned(40,8) ,
56140	 => std_logic_vector(to_unsigned(36,8) ,
56141	 => std_logic_vector(to_unsigned(35,8) ,
56142	 => std_logic_vector(to_unsigned(47,8) ,
56143	 => std_logic_vector(to_unsigned(71,8) ,
56144	 => std_logic_vector(to_unsigned(32,8) ,
56145	 => std_logic_vector(to_unsigned(24,8) ,
56146	 => std_logic_vector(to_unsigned(23,8) ,
56147	 => std_logic_vector(to_unsigned(8,8) ,
56148	 => std_logic_vector(to_unsigned(8,8) ,
56149	 => std_logic_vector(to_unsigned(13,8) ,
56150	 => std_logic_vector(to_unsigned(24,8) ,
56151	 => std_logic_vector(to_unsigned(23,8) ,
56152	 => std_logic_vector(to_unsigned(27,8) ,
56153	 => std_logic_vector(to_unsigned(27,8) ,
56154	 => std_logic_vector(to_unsigned(29,8) ,
56155	 => std_logic_vector(to_unsigned(32,8) ,
56156	 => std_logic_vector(to_unsigned(34,8) ,
56157	 => std_logic_vector(to_unsigned(29,8) ,
56158	 => std_logic_vector(to_unsigned(17,8) ,
56159	 => std_logic_vector(to_unsigned(10,8) ,
56160	 => std_logic_vector(to_unsigned(6,8) ,
56161	 => std_logic_vector(to_unsigned(29,8) ,
56162	 => std_logic_vector(to_unsigned(25,8) ,
56163	 => std_logic_vector(to_unsigned(9,8) ,
56164	 => std_logic_vector(to_unsigned(23,8) ,
56165	 => std_logic_vector(to_unsigned(28,8) ,
56166	 => std_logic_vector(to_unsigned(34,8) ,
56167	 => std_logic_vector(to_unsigned(30,8) ,
56168	 => std_logic_vector(to_unsigned(32,8) ,
56169	 => std_logic_vector(to_unsigned(32,8) ,
56170	 => std_logic_vector(to_unsigned(30,8) ,
56171	 => std_logic_vector(to_unsigned(21,8) ,
56172	 => std_logic_vector(to_unsigned(22,8) ,
56173	 => std_logic_vector(to_unsigned(24,8) ,
56174	 => std_logic_vector(to_unsigned(22,8) ,
56175	 => std_logic_vector(to_unsigned(18,8) ,
56176	 => std_logic_vector(to_unsigned(15,8) ,
56177	 => std_logic_vector(to_unsigned(13,8) ,
56178	 => std_logic_vector(to_unsigned(21,8) ,
56179	 => std_logic_vector(to_unsigned(21,8) ,
56180	 => std_logic_vector(to_unsigned(37,8) ,
56181	 => std_logic_vector(to_unsigned(38,8) ,
56182	 => std_logic_vector(to_unsigned(35,8) ,
56183	 => std_logic_vector(to_unsigned(29,8) ,
56184	 => std_logic_vector(to_unsigned(26,8) ,
56185	 => std_logic_vector(to_unsigned(30,8) ,
56186	 => std_logic_vector(to_unsigned(21,8) ,
56187	 => std_logic_vector(to_unsigned(28,8) ,
56188	 => std_logic_vector(to_unsigned(51,8) ,
56189	 => std_logic_vector(to_unsigned(43,8) ,
56190	 => std_logic_vector(to_unsigned(16,8) ,
56191	 => std_logic_vector(to_unsigned(11,8) ,
56192	 => std_logic_vector(to_unsigned(30,8) ,
56193	 => std_logic_vector(to_unsigned(21,8) ,
56194	 => std_logic_vector(to_unsigned(22,8) ,
56195	 => std_logic_vector(to_unsigned(23,8) ,
56196	 => std_logic_vector(to_unsigned(27,8) ,
56197	 => std_logic_vector(to_unsigned(33,8) ,
56198	 => std_logic_vector(to_unsigned(35,8) ,
56199	 => std_logic_vector(to_unsigned(30,8) ,
56200	 => std_logic_vector(to_unsigned(21,8) ,
56201	 => std_logic_vector(to_unsigned(39,8) ,
56202	 => std_logic_vector(to_unsigned(63,8) ,
56203	 => std_logic_vector(to_unsigned(49,8) ,
56204	 => std_logic_vector(to_unsigned(17,8) ,
56205	 => std_logic_vector(to_unsigned(26,8) ,
56206	 => std_logic_vector(to_unsigned(24,8) ,
56207	 => std_logic_vector(to_unsigned(22,8) ,
56208	 => std_logic_vector(to_unsigned(23,8) ,
56209	 => std_logic_vector(to_unsigned(17,8) ,
56210	 => std_logic_vector(to_unsigned(19,8) ,
56211	 => std_logic_vector(to_unsigned(17,8) ,
56212	 => std_logic_vector(to_unsigned(15,8) ,
56213	 => std_logic_vector(to_unsigned(13,8) ,
56214	 => std_logic_vector(to_unsigned(15,8) ,
56215	 => std_logic_vector(to_unsigned(12,8) ,
56216	 => std_logic_vector(to_unsigned(12,8) ,
56217	 => std_logic_vector(to_unsigned(12,8) ,
56218	 => std_logic_vector(to_unsigned(16,8) ,
56219	 => std_logic_vector(to_unsigned(42,8) ,
56220	 => std_logic_vector(to_unsigned(25,8) ,
56221	 => std_logic_vector(to_unsigned(14,8) ,
56222	 => std_logic_vector(to_unsigned(22,8) ,
56223	 => std_logic_vector(to_unsigned(25,8) ,
56224	 => std_logic_vector(to_unsigned(15,8) ,
56225	 => std_logic_vector(to_unsigned(7,8) ,
56226	 => std_logic_vector(to_unsigned(10,8) ,
56227	 => std_logic_vector(to_unsigned(11,8) ,
56228	 => std_logic_vector(to_unsigned(16,8) ,
56229	 => std_logic_vector(to_unsigned(18,8) ,
56230	 => std_logic_vector(to_unsigned(22,8) ,
56231	 => std_logic_vector(to_unsigned(23,8) ,
56232	 => std_logic_vector(to_unsigned(16,8) ,
56233	 => std_logic_vector(to_unsigned(15,8) ,
56234	 => std_logic_vector(to_unsigned(18,8) ,
56235	 => std_logic_vector(to_unsigned(21,8) ,
56236	 => std_logic_vector(to_unsigned(20,8) ,
56237	 => std_logic_vector(to_unsigned(17,8) ,
56238	 => std_logic_vector(to_unsigned(18,8) ,
56239	 => std_logic_vector(to_unsigned(66,8) ,
56240	 => std_logic_vector(to_unsigned(88,8) ,
56241	 => std_logic_vector(to_unsigned(87,8) ,
56242	 => std_logic_vector(to_unsigned(37,8) ,
56243	 => std_logic_vector(to_unsigned(9,8) ,
56244	 => std_logic_vector(to_unsigned(13,8) ,
56245	 => std_logic_vector(to_unsigned(13,8) ,
56246	 => std_logic_vector(to_unsigned(12,8) ,
56247	 => std_logic_vector(to_unsigned(13,8) ,
56248	 => std_logic_vector(to_unsigned(15,8) ,
56249	 => std_logic_vector(to_unsigned(12,8) ,
56250	 => std_logic_vector(to_unsigned(9,8) ,
56251	 => std_logic_vector(to_unsigned(13,8) ,
56252	 => std_logic_vector(to_unsigned(17,8) ,
56253	 => std_logic_vector(to_unsigned(19,8) ,
56254	 => std_logic_vector(to_unsigned(17,8) ,
56255	 => std_logic_vector(to_unsigned(16,8) ,
56256	 => std_logic_vector(to_unsigned(31,8) ,
56257	 => std_logic_vector(to_unsigned(33,8) ,
56258	 => std_logic_vector(to_unsigned(11,8) ,
56259	 => std_logic_vector(to_unsigned(19,8) ,
56260	 => std_logic_vector(to_unsigned(15,8) ,
56261	 => std_logic_vector(to_unsigned(1,8) ,
56262	 => std_logic_vector(to_unsigned(0,8) ,
56263	 => std_logic_vector(to_unsigned(5,8) ,
56264	 => std_logic_vector(to_unsigned(13,8) ,
56265	 => std_logic_vector(to_unsigned(18,8) ,
56266	 => std_logic_vector(to_unsigned(20,8) ,
56267	 => std_logic_vector(to_unsigned(20,8) ,
56268	 => std_logic_vector(to_unsigned(24,8) ,
56269	 => std_logic_vector(to_unsigned(22,8) ,
56270	 => std_logic_vector(to_unsigned(13,8) ,
56271	 => std_logic_vector(to_unsigned(13,8) ,
56272	 => std_logic_vector(to_unsigned(19,8) ,
56273	 => std_logic_vector(to_unsigned(14,8) ,
56274	 => std_logic_vector(to_unsigned(12,8) ,
56275	 => std_logic_vector(to_unsigned(8,8) ,
56276	 => std_logic_vector(to_unsigned(6,8) ,
56277	 => std_logic_vector(to_unsigned(8,8) ,
56278	 => std_logic_vector(to_unsigned(6,8) ,
56279	 => std_logic_vector(to_unsigned(11,8) ,
56280	 => std_logic_vector(to_unsigned(12,8) ,
56281	 => std_logic_vector(to_unsigned(1,8) ,
56282	 => std_logic_vector(to_unsigned(0,8) ,
56283	 => std_logic_vector(to_unsigned(0,8) ,
56284	 => std_logic_vector(to_unsigned(0,8) ,
56285	 => std_logic_vector(to_unsigned(0,8) ,
56286	 => std_logic_vector(to_unsigned(9,8) ,
56287	 => std_logic_vector(to_unsigned(14,8) ,
56288	 => std_logic_vector(to_unsigned(1,8) ,
56289	 => std_logic_vector(to_unsigned(10,8) ,
56290	 => std_logic_vector(to_unsigned(29,8) ,
56291	 => std_logic_vector(to_unsigned(17,8) ,
56292	 => std_logic_vector(to_unsigned(13,8) ,
56293	 => std_logic_vector(to_unsigned(20,8) ,
56294	 => std_logic_vector(to_unsigned(25,8) ,
56295	 => std_logic_vector(to_unsigned(25,8) ,
56296	 => std_logic_vector(to_unsigned(17,8) ,
56297	 => std_logic_vector(to_unsigned(13,8) ,
56298	 => std_logic_vector(to_unsigned(13,8) ,
56299	 => std_logic_vector(to_unsigned(14,8) ,
56300	 => std_logic_vector(to_unsigned(9,8) ,
56301	 => std_logic_vector(to_unsigned(13,8) ,
56302	 => std_logic_vector(to_unsigned(9,8) ,
56303	 => std_logic_vector(to_unsigned(8,8) ,
56304	 => std_logic_vector(to_unsigned(18,8) ,
56305	 => std_logic_vector(to_unsigned(14,8) ,
56306	 => std_logic_vector(to_unsigned(27,8) ,
56307	 => std_logic_vector(to_unsigned(26,8) ,
56308	 => std_logic_vector(to_unsigned(5,8) ,
56309	 => std_logic_vector(to_unsigned(7,8) ,
56310	 => std_logic_vector(to_unsigned(12,8) ,
56311	 => std_logic_vector(to_unsigned(32,8) ,
56312	 => std_logic_vector(to_unsigned(43,8) ,
56313	 => std_logic_vector(to_unsigned(29,8) ,
56314	 => std_logic_vector(to_unsigned(32,8) ,
56315	 => std_logic_vector(to_unsigned(26,8) ,
56316	 => std_logic_vector(to_unsigned(17,8) ,
56317	 => std_logic_vector(to_unsigned(27,8) ,
56318	 => std_logic_vector(to_unsigned(35,8) ,
56319	 => std_logic_vector(to_unsigned(31,8) ,
56320	 => std_logic_vector(to_unsigned(103,8) ,
56321	 => std_logic_vector(to_unsigned(99,8) ,
56322	 => std_logic_vector(to_unsigned(81,8) ,
56323	 => std_logic_vector(to_unsigned(80,8) ,
56324	 => std_logic_vector(to_unsigned(79,8) ,
56325	 => std_logic_vector(to_unsigned(48,8) ,
56326	 => std_logic_vector(to_unsigned(25,8) ,
56327	 => std_logic_vector(to_unsigned(35,8) ,
56328	 => std_logic_vector(to_unsigned(51,8) ,
56329	 => std_logic_vector(to_unsigned(43,8) ,
56330	 => std_logic_vector(to_unsigned(71,8) ,
56331	 => std_logic_vector(to_unsigned(58,8) ,
56332	 => std_logic_vector(to_unsigned(50,8) ,
56333	 => std_logic_vector(to_unsigned(91,8) ,
56334	 => std_logic_vector(to_unsigned(99,8) ,
56335	 => std_logic_vector(to_unsigned(76,8) ,
56336	 => std_logic_vector(to_unsigned(84,8) ,
56337	 => std_logic_vector(to_unsigned(87,8) ,
56338	 => std_logic_vector(to_unsigned(67,8) ,
56339	 => std_logic_vector(to_unsigned(70,8) ,
56340	 => std_logic_vector(to_unsigned(67,8) ,
56341	 => std_logic_vector(to_unsigned(35,8) ,
56342	 => std_logic_vector(to_unsigned(35,8) ,
56343	 => std_logic_vector(to_unsigned(43,8) ,
56344	 => std_logic_vector(to_unsigned(66,8) ,
56345	 => std_logic_vector(to_unsigned(93,8) ,
56346	 => std_logic_vector(to_unsigned(105,8) ,
56347	 => std_logic_vector(to_unsigned(103,8) ,
56348	 => std_logic_vector(to_unsigned(107,8) ,
56349	 => std_logic_vector(to_unsigned(82,8) ,
56350	 => std_logic_vector(to_unsigned(101,8) ,
56351	 => std_logic_vector(to_unsigned(96,8) ,
56352	 => std_logic_vector(to_unsigned(62,8) ,
56353	 => std_logic_vector(to_unsigned(55,8) ,
56354	 => std_logic_vector(to_unsigned(26,8) ,
56355	 => std_logic_vector(to_unsigned(19,8) ,
56356	 => std_logic_vector(to_unsigned(35,8) ,
56357	 => std_logic_vector(to_unsigned(70,8) ,
56358	 => std_logic_vector(to_unsigned(28,8) ,
56359	 => std_logic_vector(to_unsigned(30,8) ,
56360	 => std_logic_vector(to_unsigned(32,8) ,
56361	 => std_logic_vector(to_unsigned(28,8) ,
56362	 => std_logic_vector(to_unsigned(30,8) ,
56363	 => std_logic_vector(to_unsigned(35,8) ,
56364	 => std_logic_vector(to_unsigned(43,8) ,
56365	 => std_logic_vector(to_unsigned(50,8) ,
56366	 => std_logic_vector(to_unsigned(45,8) ,
56367	 => std_logic_vector(to_unsigned(48,8) ,
56368	 => std_logic_vector(to_unsigned(54,8) ,
56369	 => std_logic_vector(to_unsigned(45,8) ,
56370	 => std_logic_vector(to_unsigned(58,8) ,
56371	 => std_logic_vector(to_unsigned(66,8) ,
56372	 => std_logic_vector(to_unsigned(66,8) ,
56373	 => std_logic_vector(to_unsigned(76,8) ,
56374	 => std_logic_vector(to_unsigned(60,8) ,
56375	 => std_logic_vector(to_unsigned(70,8) ,
56376	 => std_logic_vector(to_unsigned(69,8) ,
56377	 => std_logic_vector(to_unsigned(45,8) ,
56378	 => std_logic_vector(to_unsigned(52,8) ,
56379	 => std_logic_vector(to_unsigned(53,8) ,
56380	 => std_logic_vector(to_unsigned(66,8) ,
56381	 => std_logic_vector(to_unsigned(49,8) ,
56382	 => std_logic_vector(to_unsigned(41,8) ,
56383	 => std_logic_vector(to_unsigned(81,8) ,
56384	 => std_logic_vector(to_unsigned(92,8) ,
56385	 => std_logic_vector(to_unsigned(79,8) ,
56386	 => std_logic_vector(to_unsigned(80,8) ,
56387	 => std_logic_vector(to_unsigned(84,8) ,
56388	 => std_logic_vector(to_unsigned(93,8) ,
56389	 => std_logic_vector(to_unsigned(96,8) ,
56390	 => std_logic_vector(to_unsigned(95,8) ,
56391	 => std_logic_vector(to_unsigned(88,8) ,
56392	 => std_logic_vector(to_unsigned(95,8) ,
56393	 => std_logic_vector(to_unsigned(93,8) ,
56394	 => std_logic_vector(to_unsigned(97,8) ,
56395	 => std_logic_vector(to_unsigned(104,8) ,
56396	 => std_logic_vector(to_unsigned(97,8) ,
56397	 => std_logic_vector(to_unsigned(115,8) ,
56398	 => std_logic_vector(to_unsigned(116,8) ,
56399	 => std_logic_vector(to_unsigned(130,8) ,
56400	 => std_logic_vector(to_unsigned(130,8) ,
56401	 => std_logic_vector(to_unsigned(115,8) ,
56402	 => std_logic_vector(to_unsigned(91,8) ,
56403	 => std_logic_vector(to_unsigned(101,8) ,
56404	 => std_logic_vector(to_unsigned(87,8) ,
56405	 => std_logic_vector(to_unsigned(51,8) ,
56406	 => std_logic_vector(to_unsigned(32,8) ,
56407	 => std_logic_vector(to_unsigned(36,8) ,
56408	 => std_logic_vector(to_unsigned(39,8) ,
56409	 => std_logic_vector(to_unsigned(39,8) ,
56410	 => std_logic_vector(to_unsigned(41,8) ,
56411	 => std_logic_vector(to_unsigned(42,8) ,
56412	 => std_logic_vector(to_unsigned(45,8) ,
56413	 => std_logic_vector(to_unsigned(47,8) ,
56414	 => std_logic_vector(to_unsigned(51,8) ,
56415	 => std_logic_vector(to_unsigned(54,8) ,
56416	 => std_logic_vector(to_unsigned(54,8) ,
56417	 => std_logic_vector(to_unsigned(55,8) ,
56418	 => std_logic_vector(to_unsigned(53,8) ,
56419	 => std_logic_vector(to_unsigned(60,8) ,
56420	 => std_logic_vector(to_unsigned(61,8) ,
56421	 => std_logic_vector(to_unsigned(60,8) ,
56422	 => std_logic_vector(to_unsigned(62,8) ,
56423	 => std_logic_vector(to_unsigned(59,8) ,
56424	 => std_logic_vector(to_unsigned(59,8) ,
56425	 => std_logic_vector(to_unsigned(60,8) ,
56426	 => std_logic_vector(to_unsigned(55,8) ,
56427	 => std_logic_vector(to_unsigned(49,8) ,
56428	 => std_logic_vector(to_unsigned(48,8) ,
56429	 => std_logic_vector(to_unsigned(46,8) ,
56430	 => std_logic_vector(to_unsigned(60,8) ,
56431	 => std_logic_vector(to_unsigned(69,8) ,
56432	 => std_logic_vector(to_unsigned(68,8) ,
56433	 => std_logic_vector(to_unsigned(79,8) ,
56434	 => std_logic_vector(to_unsigned(112,8) ,
56435	 => std_logic_vector(to_unsigned(104,8) ,
56436	 => std_logic_vector(to_unsigned(81,8) ,
56437	 => std_logic_vector(to_unsigned(55,8) ,
56438	 => std_logic_vector(to_unsigned(57,8) ,
56439	 => std_logic_vector(to_unsigned(57,8) ,
56440	 => std_logic_vector(to_unsigned(25,8) ,
56441	 => std_logic_vector(to_unsigned(11,8) ,
56442	 => std_logic_vector(to_unsigned(18,8) ,
56443	 => std_logic_vector(to_unsigned(30,8) ,
56444	 => std_logic_vector(to_unsigned(44,8) ,
56445	 => std_logic_vector(to_unsigned(50,8) ,
56446	 => std_logic_vector(to_unsigned(51,8) ,
56447	 => std_logic_vector(to_unsigned(51,8) ,
56448	 => std_logic_vector(to_unsigned(58,8) ,
56449	 => std_logic_vector(to_unsigned(71,8) ,
56450	 => std_logic_vector(to_unsigned(57,8) ,
56451	 => std_logic_vector(to_unsigned(48,8) ,
56452	 => std_logic_vector(to_unsigned(47,8) ,
56453	 => std_logic_vector(to_unsigned(44,8) ,
56454	 => std_logic_vector(to_unsigned(43,8) ,
56455	 => std_logic_vector(to_unsigned(37,8) ,
56456	 => std_logic_vector(to_unsigned(36,8) ,
56457	 => std_logic_vector(to_unsigned(38,8) ,
56458	 => std_logic_vector(to_unsigned(41,8) ,
56459	 => std_logic_vector(to_unsigned(38,8) ,
56460	 => std_logic_vector(to_unsigned(35,8) ,
56461	 => std_logic_vector(to_unsigned(50,8) ,
56462	 => std_logic_vector(to_unsigned(68,8) ,
56463	 => std_logic_vector(to_unsigned(28,8) ,
56464	 => std_logic_vector(to_unsigned(6,8) ,
56465	 => std_logic_vector(to_unsigned(29,8) ,
56466	 => std_logic_vector(to_unsigned(32,8) ,
56467	 => std_logic_vector(to_unsigned(9,8) ,
56468	 => std_logic_vector(to_unsigned(5,8) ,
56469	 => std_logic_vector(to_unsigned(6,8) ,
56470	 => std_logic_vector(to_unsigned(54,8) ,
56471	 => std_logic_vector(to_unsigned(14,8) ,
56472	 => std_logic_vector(to_unsigned(24,8) ,
56473	 => std_logic_vector(to_unsigned(41,8) ,
56474	 => std_logic_vector(to_unsigned(34,8) ,
56475	 => std_logic_vector(to_unsigned(29,8) ,
56476	 => std_logic_vector(to_unsigned(23,8) ,
56477	 => std_logic_vector(to_unsigned(24,8) ,
56478	 => std_logic_vector(to_unsigned(17,8) ,
56479	 => std_logic_vector(to_unsigned(19,8) ,
56480	 => std_logic_vector(to_unsigned(23,8) ,
56481	 => std_logic_vector(to_unsigned(38,8) ,
56482	 => std_logic_vector(to_unsigned(29,8) ,
56483	 => std_logic_vector(to_unsigned(19,8) ,
56484	 => std_logic_vector(to_unsigned(27,8) ,
56485	 => std_logic_vector(to_unsigned(23,8) ,
56486	 => std_logic_vector(to_unsigned(38,8) ,
56487	 => std_logic_vector(to_unsigned(22,8) ,
56488	 => std_logic_vector(to_unsigned(11,8) ,
56489	 => std_logic_vector(to_unsigned(15,8) ,
56490	 => std_logic_vector(to_unsigned(13,8) ,
56491	 => std_logic_vector(to_unsigned(25,8) ,
56492	 => std_logic_vector(to_unsigned(24,8) ,
56493	 => std_logic_vector(to_unsigned(27,8) ,
56494	 => std_logic_vector(to_unsigned(32,8) ,
56495	 => std_logic_vector(to_unsigned(43,8) ,
56496	 => std_logic_vector(to_unsigned(37,8) ,
56497	 => std_logic_vector(to_unsigned(27,8) ,
56498	 => std_logic_vector(to_unsigned(35,8) ,
56499	 => std_logic_vector(to_unsigned(31,8) ,
56500	 => std_logic_vector(to_unsigned(37,8) ,
56501	 => std_logic_vector(to_unsigned(41,8) ,
56502	 => std_logic_vector(to_unsigned(37,8) ,
56503	 => std_logic_vector(to_unsigned(37,8) ,
56504	 => std_logic_vector(to_unsigned(50,8) ,
56505	 => std_logic_vector(to_unsigned(29,8) ,
56506	 => std_logic_vector(to_unsigned(26,8) ,
56507	 => std_logic_vector(to_unsigned(52,8) ,
56508	 => std_logic_vector(to_unsigned(41,8) ,
56509	 => std_logic_vector(to_unsigned(17,8) ,
56510	 => std_logic_vector(to_unsigned(12,8) ,
56511	 => std_logic_vector(to_unsigned(41,8) ,
56512	 => std_logic_vector(to_unsigned(40,8) ,
56513	 => std_logic_vector(to_unsigned(17,8) ,
56514	 => std_logic_vector(to_unsigned(19,8) ,
56515	 => std_logic_vector(to_unsigned(8,8) ,
56516	 => std_logic_vector(to_unsigned(23,8) ,
56517	 => std_logic_vector(to_unsigned(16,8) ,
56518	 => std_logic_vector(to_unsigned(10,8) ,
56519	 => std_logic_vector(to_unsigned(17,8) ,
56520	 => std_logic_vector(to_unsigned(25,8) ,
56521	 => std_logic_vector(to_unsigned(19,8) ,
56522	 => std_logic_vector(to_unsigned(26,8) ,
56523	 => std_logic_vector(to_unsigned(27,8) ,
56524	 => std_logic_vector(to_unsigned(22,8) ,
56525	 => std_logic_vector(to_unsigned(24,8) ,
56526	 => std_logic_vector(to_unsigned(32,8) ,
56527	 => std_logic_vector(to_unsigned(41,8) ,
56528	 => std_logic_vector(to_unsigned(35,8) ,
56529	 => std_logic_vector(to_unsigned(17,8) ,
56530	 => std_logic_vector(to_unsigned(14,8) ,
56531	 => std_logic_vector(to_unsigned(20,8) ,
56532	 => std_logic_vector(to_unsigned(23,8) ,
56533	 => std_logic_vector(to_unsigned(28,8) ,
56534	 => std_logic_vector(to_unsigned(13,8) ,
56535	 => std_logic_vector(to_unsigned(10,8) ,
56536	 => std_logic_vector(to_unsigned(17,8) ,
56537	 => std_logic_vector(to_unsigned(19,8) ,
56538	 => std_logic_vector(to_unsigned(15,8) ,
56539	 => std_logic_vector(to_unsigned(29,8) ,
56540	 => std_logic_vector(to_unsigned(42,8) ,
56541	 => std_logic_vector(to_unsigned(35,8) ,
56542	 => std_logic_vector(to_unsigned(22,8) ,
56543	 => std_logic_vector(to_unsigned(19,8) ,
56544	 => std_logic_vector(to_unsigned(10,8) ,
56545	 => std_logic_vector(to_unsigned(5,8) ,
56546	 => std_logic_vector(to_unsigned(9,8) ,
56547	 => std_logic_vector(to_unsigned(13,8) ,
56548	 => std_logic_vector(to_unsigned(13,8) ,
56549	 => std_logic_vector(to_unsigned(11,8) ,
56550	 => std_logic_vector(to_unsigned(13,8) ,
56551	 => std_logic_vector(to_unsigned(17,8) ,
56552	 => std_logic_vector(to_unsigned(17,8) ,
56553	 => std_logic_vector(to_unsigned(16,8) ,
56554	 => std_logic_vector(to_unsigned(22,8) ,
56555	 => std_logic_vector(to_unsigned(23,8) ,
56556	 => std_logic_vector(to_unsigned(27,8) ,
56557	 => std_logic_vector(to_unsigned(23,8) ,
56558	 => std_logic_vector(to_unsigned(26,8) ,
56559	 => std_logic_vector(to_unsigned(65,8) ,
56560	 => std_logic_vector(to_unsigned(86,8) ,
56561	 => std_logic_vector(to_unsigned(90,8) ,
56562	 => std_logic_vector(to_unsigned(35,8) ,
56563	 => std_logic_vector(to_unsigned(10,8) ,
56564	 => std_logic_vector(to_unsigned(16,8) ,
56565	 => std_logic_vector(to_unsigned(12,8) ,
56566	 => std_logic_vector(to_unsigned(10,8) ,
56567	 => std_logic_vector(to_unsigned(13,8) ,
56568	 => std_logic_vector(to_unsigned(16,8) ,
56569	 => std_logic_vector(to_unsigned(10,8) ,
56570	 => std_logic_vector(to_unsigned(9,8) ,
56571	 => std_logic_vector(to_unsigned(14,8) ,
56572	 => std_logic_vector(to_unsigned(15,8) ,
56573	 => std_logic_vector(to_unsigned(16,8) ,
56574	 => std_logic_vector(to_unsigned(13,8) ,
56575	 => std_logic_vector(to_unsigned(11,8) ,
56576	 => std_logic_vector(to_unsigned(17,8) ,
56577	 => std_logic_vector(to_unsigned(19,8) ,
56578	 => std_logic_vector(to_unsigned(11,8) ,
56579	 => std_logic_vector(to_unsigned(12,8) ,
56580	 => std_logic_vector(to_unsigned(17,8) ,
56581	 => std_logic_vector(to_unsigned(3,8) ,
56582	 => std_logic_vector(to_unsigned(0,8) ,
56583	 => std_logic_vector(to_unsigned(2,8) ,
56584	 => std_logic_vector(to_unsigned(18,8) ,
56585	 => std_logic_vector(to_unsigned(28,8) ,
56586	 => std_logic_vector(to_unsigned(22,8) ,
56587	 => std_logic_vector(to_unsigned(22,8) ,
56588	 => std_logic_vector(to_unsigned(17,8) ,
56589	 => std_logic_vector(to_unsigned(16,8) ,
56590	 => std_logic_vector(to_unsigned(16,8) ,
56591	 => std_logic_vector(to_unsigned(16,8) ,
56592	 => std_logic_vector(to_unsigned(18,8) ,
56593	 => std_logic_vector(to_unsigned(11,8) ,
56594	 => std_logic_vector(to_unsigned(9,8) ,
56595	 => std_logic_vector(to_unsigned(8,8) ,
56596	 => std_logic_vector(to_unsigned(8,8) ,
56597	 => std_logic_vector(to_unsigned(9,8) ,
56598	 => std_logic_vector(to_unsigned(6,8) ,
56599	 => std_logic_vector(to_unsigned(10,8) ,
56600	 => std_logic_vector(to_unsigned(7,8) ,
56601	 => std_logic_vector(to_unsigned(1,8) ,
56602	 => std_logic_vector(to_unsigned(0,8) ,
56603	 => std_logic_vector(to_unsigned(0,8) ,
56604	 => std_logic_vector(to_unsigned(0,8) ,
56605	 => std_logic_vector(to_unsigned(0,8) ,
56606	 => std_logic_vector(to_unsigned(8,8) ,
56607	 => std_logic_vector(to_unsigned(30,8) ,
56608	 => std_logic_vector(to_unsigned(17,8) ,
56609	 => std_logic_vector(to_unsigned(27,8) ,
56610	 => std_logic_vector(to_unsigned(33,8) ,
56611	 => std_logic_vector(to_unsigned(20,8) ,
56612	 => std_logic_vector(to_unsigned(19,8) ,
56613	 => std_logic_vector(to_unsigned(20,8) ,
56614	 => std_logic_vector(to_unsigned(16,8) ,
56615	 => std_logic_vector(to_unsigned(14,8) ,
56616	 => std_logic_vector(to_unsigned(19,8) ,
56617	 => std_logic_vector(to_unsigned(19,8) ,
56618	 => std_logic_vector(to_unsigned(25,8) ,
56619	 => std_logic_vector(to_unsigned(19,8) ,
56620	 => std_logic_vector(to_unsigned(8,8) ,
56621	 => std_logic_vector(to_unsigned(12,8) ,
56622	 => std_logic_vector(to_unsigned(8,8) ,
56623	 => std_logic_vector(to_unsigned(7,8) ,
56624	 => std_logic_vector(to_unsigned(11,8) ,
56625	 => std_logic_vector(to_unsigned(5,8) ,
56626	 => std_logic_vector(to_unsigned(25,8) ,
56627	 => std_logic_vector(to_unsigned(30,8) ,
56628	 => std_logic_vector(to_unsigned(3,8) ,
56629	 => std_logic_vector(to_unsigned(5,8) ,
56630	 => std_logic_vector(to_unsigned(5,8) ,
56631	 => std_logic_vector(to_unsigned(16,8) ,
56632	 => std_logic_vector(to_unsigned(30,8) ,
56633	 => std_logic_vector(to_unsigned(30,8) ,
56634	 => std_logic_vector(to_unsigned(32,8) ,
56635	 => std_logic_vector(to_unsigned(29,8) ,
56636	 => std_logic_vector(to_unsigned(18,8) ,
56637	 => std_logic_vector(to_unsigned(39,8) ,
56638	 => std_logic_vector(to_unsigned(32,8) ,
56639	 => std_logic_vector(to_unsigned(27,8) ,
56640	 => std_logic_vector(to_unsigned(62,8) ,
56641	 => std_logic_vector(to_unsigned(96,8) ,
56642	 => std_logic_vector(to_unsigned(82,8) ,
56643	 => std_logic_vector(to_unsigned(76,8) ,
56644	 => std_logic_vector(to_unsigned(74,8) ,
56645	 => std_logic_vector(to_unsigned(44,8) ,
56646	 => std_logic_vector(to_unsigned(30,8) ,
56647	 => std_logic_vector(to_unsigned(35,8) ,
56648	 => std_logic_vector(to_unsigned(57,8) ,
56649	 => std_logic_vector(to_unsigned(59,8) ,
56650	 => std_logic_vector(to_unsigned(76,8) ,
56651	 => std_logic_vector(to_unsigned(63,8) ,
56652	 => std_logic_vector(to_unsigned(52,8) ,
56653	 => std_logic_vector(to_unsigned(85,8) ,
56654	 => std_logic_vector(to_unsigned(101,8) ,
56655	 => std_logic_vector(to_unsigned(73,8) ,
56656	 => std_logic_vector(to_unsigned(72,8) ,
56657	 => std_logic_vector(to_unsigned(86,8) ,
56658	 => std_logic_vector(to_unsigned(62,8) ,
56659	 => std_logic_vector(to_unsigned(62,8) ,
56660	 => std_logic_vector(to_unsigned(80,8) ,
56661	 => std_logic_vector(to_unsigned(44,8) ,
56662	 => std_logic_vector(to_unsigned(37,8) ,
56663	 => std_logic_vector(to_unsigned(88,8) ,
56664	 => std_logic_vector(to_unsigned(92,8) ,
56665	 => std_logic_vector(to_unsigned(96,8) ,
56666	 => std_logic_vector(to_unsigned(116,8) ,
56667	 => std_logic_vector(to_unsigned(85,8) ,
56668	 => std_logic_vector(to_unsigned(76,8) ,
56669	 => std_logic_vector(to_unsigned(59,8) ,
56670	 => std_logic_vector(to_unsigned(82,8) ,
56671	 => std_logic_vector(to_unsigned(105,8) ,
56672	 => std_logic_vector(to_unsigned(80,8) ,
56673	 => std_logic_vector(to_unsigned(61,8) ,
56674	 => std_logic_vector(to_unsigned(29,8) ,
56675	 => std_logic_vector(to_unsigned(23,8) ,
56676	 => std_logic_vector(to_unsigned(37,8) ,
56677	 => std_logic_vector(to_unsigned(81,8) ,
56678	 => std_logic_vector(to_unsigned(37,8) ,
56679	 => std_logic_vector(to_unsigned(58,8) ,
56680	 => std_logic_vector(to_unsigned(65,8) ,
56681	 => std_logic_vector(to_unsigned(52,8) ,
56682	 => std_logic_vector(to_unsigned(42,8) ,
56683	 => std_logic_vector(to_unsigned(41,8) ,
56684	 => std_logic_vector(to_unsigned(41,8) ,
56685	 => std_logic_vector(to_unsigned(41,8) ,
56686	 => std_logic_vector(to_unsigned(41,8) ,
56687	 => std_logic_vector(to_unsigned(41,8) ,
56688	 => std_logic_vector(to_unsigned(39,8) ,
56689	 => std_logic_vector(to_unsigned(46,8) ,
56690	 => std_logic_vector(to_unsigned(62,8) ,
56691	 => std_logic_vector(to_unsigned(60,8) ,
56692	 => std_logic_vector(to_unsigned(52,8) ,
56693	 => std_logic_vector(to_unsigned(65,8) ,
56694	 => std_logic_vector(to_unsigned(47,8) ,
56695	 => std_logic_vector(to_unsigned(48,8) ,
56696	 => std_logic_vector(to_unsigned(69,8) ,
56697	 => std_logic_vector(to_unsigned(63,8) ,
56698	 => std_logic_vector(to_unsigned(60,8) ,
56699	 => std_logic_vector(to_unsigned(58,8) ,
56700	 => std_logic_vector(to_unsigned(68,8) ,
56701	 => std_logic_vector(to_unsigned(51,8) ,
56702	 => std_logic_vector(to_unsigned(37,8) ,
56703	 => std_logic_vector(to_unsigned(85,8) ,
56704	 => std_logic_vector(to_unsigned(109,8) ,
56705	 => std_logic_vector(to_unsigned(95,8) ,
56706	 => std_logic_vector(to_unsigned(100,8) ,
56707	 => std_logic_vector(to_unsigned(85,8) ,
56708	 => std_logic_vector(to_unsigned(82,8) ,
56709	 => std_logic_vector(to_unsigned(87,8) ,
56710	 => std_logic_vector(to_unsigned(92,8) ,
56711	 => std_logic_vector(to_unsigned(92,8) ,
56712	 => std_logic_vector(to_unsigned(90,8) ,
56713	 => std_logic_vector(to_unsigned(85,8) ,
56714	 => std_logic_vector(to_unsigned(93,8) ,
56715	 => std_logic_vector(to_unsigned(109,8) ,
56716	 => std_logic_vector(to_unsigned(115,8) ,
56717	 => std_logic_vector(to_unsigned(133,8) ,
56718	 => std_logic_vector(to_unsigned(133,8) ,
56719	 => std_logic_vector(to_unsigned(131,8) ,
56720	 => std_logic_vector(to_unsigned(128,8) ,
56721	 => std_logic_vector(to_unsigned(104,8) ,
56722	 => std_logic_vector(to_unsigned(84,8) ,
56723	 => std_logic_vector(to_unsigned(84,8) ,
56724	 => std_logic_vector(to_unsigned(74,8) ,
56725	 => std_logic_vector(to_unsigned(71,8) ,
56726	 => std_logic_vector(to_unsigned(32,8) ,
56727	 => std_logic_vector(to_unsigned(32,8) ,
56728	 => std_logic_vector(to_unsigned(37,8) ,
56729	 => std_logic_vector(to_unsigned(39,8) ,
56730	 => std_logic_vector(to_unsigned(40,8) ,
56731	 => std_logic_vector(to_unsigned(39,8) ,
56732	 => std_logic_vector(to_unsigned(39,8) ,
56733	 => std_logic_vector(to_unsigned(42,8) ,
56734	 => std_logic_vector(to_unsigned(50,8) ,
56735	 => std_logic_vector(to_unsigned(54,8) ,
56736	 => std_logic_vector(to_unsigned(55,8) ,
56737	 => std_logic_vector(to_unsigned(57,8) ,
56738	 => std_logic_vector(to_unsigned(54,8) ,
56739	 => std_logic_vector(to_unsigned(60,8) ,
56740	 => std_logic_vector(to_unsigned(59,8) ,
56741	 => std_logic_vector(to_unsigned(55,8) ,
56742	 => std_logic_vector(to_unsigned(58,8) ,
56743	 => std_logic_vector(to_unsigned(60,8) ,
56744	 => std_logic_vector(to_unsigned(59,8) ,
56745	 => std_logic_vector(to_unsigned(54,8) ,
56746	 => std_logic_vector(to_unsigned(55,8) ,
56747	 => std_logic_vector(to_unsigned(52,8) ,
56748	 => std_logic_vector(to_unsigned(61,8) ,
56749	 => std_logic_vector(to_unsigned(66,8) ,
56750	 => std_logic_vector(to_unsigned(62,8) ,
56751	 => std_logic_vector(to_unsigned(68,8) ,
56752	 => std_logic_vector(to_unsigned(96,8) ,
56753	 => std_logic_vector(to_unsigned(111,8) ,
56754	 => std_logic_vector(to_unsigned(80,8) ,
56755	 => std_logic_vector(to_unsigned(61,8) ,
56756	 => std_logic_vector(to_unsigned(76,8) ,
56757	 => std_logic_vector(to_unsigned(54,8) ,
56758	 => std_logic_vector(to_unsigned(63,8) ,
56759	 => std_logic_vector(to_unsigned(60,8) ,
56760	 => std_logic_vector(to_unsigned(24,8) ,
56761	 => std_logic_vector(to_unsigned(17,8) ,
56762	 => std_logic_vector(to_unsigned(34,8) ,
56763	 => std_logic_vector(to_unsigned(51,8) ,
56764	 => std_logic_vector(to_unsigned(58,8) ,
56765	 => std_logic_vector(to_unsigned(61,8) ,
56766	 => std_logic_vector(to_unsigned(65,8) ,
56767	 => std_logic_vector(to_unsigned(62,8) ,
56768	 => std_logic_vector(to_unsigned(67,8) ,
56769	 => std_logic_vector(to_unsigned(64,8) ,
56770	 => std_logic_vector(to_unsigned(35,8) ,
56771	 => std_logic_vector(to_unsigned(29,8) ,
56772	 => std_logic_vector(to_unsigned(37,8) ,
56773	 => std_logic_vector(to_unsigned(36,8) ,
56774	 => std_logic_vector(to_unsigned(41,8) ,
56775	 => std_logic_vector(to_unsigned(37,8) ,
56776	 => std_logic_vector(to_unsigned(35,8) ,
56777	 => std_logic_vector(to_unsigned(40,8) ,
56778	 => std_logic_vector(to_unsigned(36,8) ,
56779	 => std_logic_vector(to_unsigned(40,8) ,
56780	 => std_logic_vector(to_unsigned(57,8) ,
56781	 => std_logic_vector(to_unsigned(51,8) ,
56782	 => std_logic_vector(to_unsigned(23,8) ,
56783	 => std_logic_vector(to_unsigned(11,8) ,
56784	 => std_logic_vector(to_unsigned(11,8) ,
56785	 => std_logic_vector(to_unsigned(30,8) ,
56786	 => std_logic_vector(to_unsigned(40,8) ,
56787	 => std_logic_vector(to_unsigned(11,8) ,
56788	 => std_logic_vector(to_unsigned(7,8) ,
56789	 => std_logic_vector(to_unsigned(8,8) ,
56790	 => std_logic_vector(to_unsigned(65,8) ,
56791	 => std_logic_vector(to_unsigned(33,8) ,
56792	 => std_logic_vector(to_unsigned(40,8) ,
56793	 => std_logic_vector(to_unsigned(54,8) ,
56794	 => std_logic_vector(to_unsigned(59,8) ,
56795	 => std_logic_vector(to_unsigned(17,8) ,
56796	 => std_logic_vector(to_unsigned(22,8) ,
56797	 => std_logic_vector(to_unsigned(39,8) ,
56798	 => std_logic_vector(to_unsigned(4,8) ,
56799	 => std_logic_vector(to_unsigned(5,8) ,
56800	 => std_logic_vector(to_unsigned(6,8) ,
56801	 => std_logic_vector(to_unsigned(18,8) ,
56802	 => std_logic_vector(to_unsigned(32,8) ,
56803	 => std_logic_vector(to_unsigned(32,8) ,
56804	 => std_logic_vector(to_unsigned(29,8) ,
56805	 => std_logic_vector(to_unsigned(54,8) ,
56806	 => std_logic_vector(to_unsigned(44,8) ,
56807	 => std_logic_vector(to_unsigned(15,8) ,
56808	 => std_logic_vector(to_unsigned(19,8) ,
56809	 => std_logic_vector(to_unsigned(16,8) ,
56810	 => std_logic_vector(to_unsigned(8,8) ,
56811	 => std_logic_vector(to_unsigned(16,8) ,
56812	 => std_logic_vector(to_unsigned(20,8) ,
56813	 => std_logic_vector(to_unsigned(18,8) ,
56814	 => std_logic_vector(to_unsigned(27,8) ,
56815	 => std_logic_vector(to_unsigned(45,8) ,
56816	 => std_logic_vector(to_unsigned(47,8) ,
56817	 => std_logic_vector(to_unsigned(45,8) ,
56818	 => std_logic_vector(to_unsigned(49,8) ,
56819	 => std_logic_vector(to_unsigned(49,8) ,
56820	 => std_logic_vector(to_unsigned(50,8) ,
56821	 => std_logic_vector(to_unsigned(54,8) ,
56822	 => std_logic_vector(to_unsigned(43,8) ,
56823	 => std_logic_vector(to_unsigned(41,8) ,
56824	 => std_logic_vector(to_unsigned(24,8) ,
56825	 => std_logic_vector(to_unsigned(14,8) ,
56826	 => std_logic_vector(to_unsigned(21,8) ,
56827	 => std_logic_vector(to_unsigned(37,8) ,
56828	 => std_logic_vector(to_unsigned(32,8) ,
56829	 => std_logic_vector(to_unsigned(24,8) ,
56830	 => std_logic_vector(to_unsigned(45,8) ,
56831	 => std_logic_vector(to_unsigned(62,8) ,
56832	 => std_logic_vector(to_unsigned(19,8) ,
56833	 => std_logic_vector(to_unsigned(8,8) ,
56834	 => std_logic_vector(to_unsigned(7,8) ,
56835	 => std_logic_vector(to_unsigned(8,8) ,
56836	 => std_logic_vector(to_unsigned(23,8) ,
56837	 => std_logic_vector(to_unsigned(20,8) ,
56838	 => std_logic_vector(to_unsigned(10,8) ,
56839	 => std_logic_vector(to_unsigned(16,8) ,
56840	 => std_logic_vector(to_unsigned(27,8) ,
56841	 => std_logic_vector(to_unsigned(8,8) ,
56842	 => std_logic_vector(to_unsigned(3,8) ,
56843	 => std_logic_vector(to_unsigned(10,8) ,
56844	 => std_logic_vector(to_unsigned(27,8) ,
56845	 => std_logic_vector(to_unsigned(23,8) ,
56846	 => std_logic_vector(to_unsigned(17,8) ,
56847	 => std_logic_vector(to_unsigned(17,8) ,
56848	 => std_logic_vector(to_unsigned(23,8) ,
56849	 => std_logic_vector(to_unsigned(24,8) ,
56850	 => std_logic_vector(to_unsigned(17,8) ,
56851	 => std_logic_vector(to_unsigned(22,8) ,
56852	 => std_logic_vector(to_unsigned(30,8) ,
56853	 => std_logic_vector(to_unsigned(29,8) ,
56854	 => std_logic_vector(to_unsigned(17,8) ,
56855	 => std_logic_vector(to_unsigned(18,8) ,
56856	 => std_logic_vector(to_unsigned(31,8) ,
56857	 => std_logic_vector(to_unsigned(26,8) ,
56858	 => std_logic_vector(to_unsigned(15,8) ,
56859	 => std_logic_vector(to_unsigned(30,8) ,
56860	 => std_logic_vector(to_unsigned(77,8) ,
56861	 => std_logic_vector(to_unsigned(119,8) ,
56862	 => std_logic_vector(to_unsigned(72,8) ,
56863	 => std_logic_vector(to_unsigned(37,8) ,
56864	 => std_logic_vector(to_unsigned(10,8) ,
56865	 => std_logic_vector(to_unsigned(6,8) ,
56866	 => std_logic_vector(to_unsigned(7,8) ,
56867	 => std_logic_vector(to_unsigned(12,8) ,
56868	 => std_logic_vector(to_unsigned(13,8) ,
56869	 => std_logic_vector(to_unsigned(12,8) ,
56870	 => std_logic_vector(to_unsigned(10,8) ,
56871	 => std_logic_vector(to_unsigned(13,8) ,
56872	 => std_logic_vector(to_unsigned(17,8) ,
56873	 => std_logic_vector(to_unsigned(17,8) ,
56874	 => std_logic_vector(to_unsigned(14,8) ,
56875	 => std_logic_vector(to_unsigned(16,8) ,
56876	 => std_logic_vector(to_unsigned(22,8) ,
56877	 => std_logic_vector(to_unsigned(22,8) ,
56878	 => std_logic_vector(to_unsigned(25,8) ,
56879	 => std_logic_vector(to_unsigned(58,8) ,
56880	 => std_logic_vector(to_unsigned(71,8) ,
56881	 => std_logic_vector(to_unsigned(74,8) ,
56882	 => std_logic_vector(to_unsigned(27,8) ,
56883	 => std_logic_vector(to_unsigned(9,8) ,
56884	 => std_logic_vector(to_unsigned(14,8) ,
56885	 => std_logic_vector(to_unsigned(10,8) ,
56886	 => std_logic_vector(to_unsigned(11,8) ,
56887	 => std_logic_vector(to_unsigned(14,8) ,
56888	 => std_logic_vector(to_unsigned(12,8) ,
56889	 => std_logic_vector(to_unsigned(9,8) ,
56890	 => std_logic_vector(to_unsigned(10,8) ,
56891	 => std_logic_vector(to_unsigned(12,8) ,
56892	 => std_logic_vector(to_unsigned(11,8) ,
56893	 => std_logic_vector(to_unsigned(12,8) ,
56894	 => std_logic_vector(to_unsigned(11,8) ,
56895	 => std_logic_vector(to_unsigned(9,8) ,
56896	 => std_logic_vector(to_unsigned(9,8) ,
56897	 => std_logic_vector(to_unsigned(10,8) ,
56898	 => std_logic_vector(to_unsigned(14,8) ,
56899	 => std_logic_vector(to_unsigned(15,8) ,
56900	 => std_logic_vector(to_unsigned(16,8) ,
56901	 => std_logic_vector(to_unsigned(6,8) ,
56902	 => std_logic_vector(to_unsigned(0,8) ,
56903	 => std_logic_vector(to_unsigned(1,8) ,
56904	 => std_logic_vector(to_unsigned(18,8) ,
56905	 => std_logic_vector(to_unsigned(26,8) ,
56906	 => std_logic_vector(to_unsigned(24,8) ,
56907	 => std_logic_vector(to_unsigned(22,8) ,
56908	 => std_logic_vector(to_unsigned(12,8) ,
56909	 => std_logic_vector(to_unsigned(16,8) ,
56910	 => std_logic_vector(to_unsigned(25,8) ,
56911	 => std_logic_vector(to_unsigned(22,8) ,
56912	 => std_logic_vector(to_unsigned(16,8) ,
56913	 => std_logic_vector(to_unsigned(6,8) ,
56914	 => std_logic_vector(to_unsigned(4,8) ,
56915	 => std_logic_vector(to_unsigned(5,8) ,
56916	 => std_logic_vector(to_unsigned(7,8) ,
56917	 => std_logic_vector(to_unsigned(9,8) ,
56918	 => std_logic_vector(to_unsigned(8,8) ,
56919	 => std_logic_vector(to_unsigned(10,8) ,
56920	 => std_logic_vector(to_unsigned(8,8) ,
56921	 => std_logic_vector(to_unsigned(3,8) ,
56922	 => std_logic_vector(to_unsigned(0,8) ,
56923	 => std_logic_vector(to_unsigned(0,8) ,
56924	 => std_logic_vector(to_unsigned(0,8) ,
56925	 => std_logic_vector(to_unsigned(0,8) ,
56926	 => std_logic_vector(to_unsigned(4,8) ,
56927	 => std_logic_vector(to_unsigned(14,8) ,
56928	 => std_logic_vector(to_unsigned(8,8) ,
56929	 => std_logic_vector(to_unsigned(15,8) ,
56930	 => std_logic_vector(to_unsigned(17,8) ,
56931	 => std_logic_vector(to_unsigned(17,8) ,
56932	 => std_logic_vector(to_unsigned(17,8) ,
56933	 => std_logic_vector(to_unsigned(22,8) ,
56934	 => std_logic_vector(to_unsigned(10,8) ,
56935	 => std_logic_vector(to_unsigned(7,8) ,
56936	 => std_logic_vector(to_unsigned(8,8) ,
56937	 => std_logic_vector(to_unsigned(6,8) ,
56938	 => std_logic_vector(to_unsigned(8,8) ,
56939	 => std_logic_vector(to_unsigned(10,8) ,
56940	 => std_logic_vector(to_unsigned(6,8) ,
56941	 => std_logic_vector(to_unsigned(7,8) ,
56942	 => std_logic_vector(to_unsigned(8,8) ,
56943	 => std_logic_vector(to_unsigned(9,8) ,
56944	 => std_logic_vector(to_unsigned(8,8) ,
56945	 => std_logic_vector(to_unsigned(6,8) ,
56946	 => std_logic_vector(to_unsigned(10,8) ,
56947	 => std_logic_vector(to_unsigned(11,8) ,
56948	 => std_logic_vector(to_unsigned(8,8) ,
56949	 => std_logic_vector(to_unsigned(11,8) ,
56950	 => std_logic_vector(to_unsigned(9,8) ,
56951	 => std_logic_vector(to_unsigned(7,8) ,
56952	 => std_logic_vector(to_unsigned(8,8) ,
56953	 => std_logic_vector(to_unsigned(11,8) ,
56954	 => std_logic_vector(to_unsigned(13,8) ,
56955	 => std_logic_vector(to_unsigned(11,8) ,
56956	 => std_logic_vector(to_unsigned(3,8) ,
56957	 => std_logic_vector(to_unsigned(10,8) ,
56958	 => std_logic_vector(to_unsigned(13,8) ,
56959	 => std_logic_vector(to_unsigned(12,8) ,
56960	 => std_logic_vector(to_unsigned(24,8) ,
56961	 => std_logic_vector(to_unsigned(92,8) ,
56962	 => std_logic_vector(to_unsigned(63,8) ,
56963	 => std_logic_vector(to_unsigned(65,8) ,
56964	 => std_logic_vector(to_unsigned(81,8) ,
56965	 => std_logic_vector(to_unsigned(51,8) ,
56966	 => std_logic_vector(to_unsigned(32,8) ,
56967	 => std_logic_vector(to_unsigned(35,8) ,
56968	 => std_logic_vector(to_unsigned(57,8) ,
56969	 => std_logic_vector(to_unsigned(49,8) ,
56970	 => std_logic_vector(to_unsigned(85,8) ,
56971	 => std_logic_vector(to_unsigned(68,8) ,
56972	 => std_logic_vector(to_unsigned(50,8) ,
56973	 => std_logic_vector(to_unsigned(82,8) ,
56974	 => std_logic_vector(to_unsigned(105,8) ,
56975	 => std_logic_vector(to_unsigned(56,8) ,
56976	 => std_logic_vector(to_unsigned(49,8) ,
56977	 => std_logic_vector(to_unsigned(92,8) ,
56978	 => std_logic_vector(to_unsigned(77,8) ,
56979	 => std_logic_vector(to_unsigned(84,8) ,
56980	 => std_logic_vector(to_unsigned(95,8) ,
56981	 => std_logic_vector(to_unsigned(82,8) ,
56982	 => std_logic_vector(to_unsigned(41,8) ,
56983	 => std_logic_vector(to_unsigned(50,8) ,
56984	 => std_logic_vector(to_unsigned(81,8) ,
56985	 => std_logic_vector(to_unsigned(80,8) ,
56986	 => std_logic_vector(to_unsigned(78,8) ,
56987	 => std_logic_vector(to_unsigned(87,8) ,
56988	 => std_logic_vector(to_unsigned(56,8) ,
56989	 => std_logic_vector(to_unsigned(47,8) ,
56990	 => std_logic_vector(to_unsigned(78,8) ,
56991	 => std_logic_vector(to_unsigned(100,8) ,
56992	 => std_logic_vector(to_unsigned(90,8) ,
56993	 => std_logic_vector(to_unsigned(68,8) ,
56994	 => std_logic_vector(to_unsigned(28,8) ,
56995	 => std_logic_vector(to_unsigned(20,8) ,
56996	 => std_logic_vector(to_unsigned(32,8) ,
56997	 => std_logic_vector(to_unsigned(74,8) ,
56998	 => std_logic_vector(to_unsigned(41,8) ,
56999	 => std_logic_vector(to_unsigned(43,8) ,
57000	 => std_logic_vector(to_unsigned(69,8) ,
57001	 => std_logic_vector(to_unsigned(59,8) ,
57002	 => std_logic_vector(to_unsigned(35,8) ,
57003	 => std_logic_vector(to_unsigned(39,8) ,
57004	 => std_logic_vector(to_unsigned(49,8) ,
57005	 => std_logic_vector(to_unsigned(43,8) ,
57006	 => std_logic_vector(to_unsigned(47,8) ,
57007	 => std_logic_vector(to_unsigned(51,8) ,
57008	 => std_logic_vector(to_unsigned(48,8) ,
57009	 => std_logic_vector(to_unsigned(49,8) ,
57010	 => std_logic_vector(to_unsigned(55,8) ,
57011	 => std_logic_vector(to_unsigned(62,8) ,
57012	 => std_logic_vector(to_unsigned(61,8) ,
57013	 => std_logic_vector(to_unsigned(64,8) ,
57014	 => std_logic_vector(to_unsigned(56,8) ,
57015	 => std_logic_vector(to_unsigned(44,8) ,
57016	 => std_logic_vector(to_unsigned(59,8) ,
57017	 => std_logic_vector(to_unsigned(71,8) ,
57018	 => std_logic_vector(to_unsigned(58,8) ,
57019	 => std_logic_vector(to_unsigned(48,8) ,
57020	 => std_logic_vector(to_unsigned(57,8) ,
57021	 => std_logic_vector(to_unsigned(65,8) ,
57022	 => std_logic_vector(to_unsigned(52,8) ,
57023	 => std_logic_vector(to_unsigned(82,8) ,
57024	 => std_logic_vector(to_unsigned(103,8) ,
57025	 => std_logic_vector(to_unsigned(99,8) ,
57026	 => std_logic_vector(to_unsigned(112,8) ,
57027	 => std_logic_vector(to_unsigned(86,8) ,
57028	 => std_logic_vector(to_unsigned(96,8) ,
57029	 => std_logic_vector(to_unsigned(111,8) ,
57030	 => std_logic_vector(to_unsigned(96,8) ,
57031	 => std_logic_vector(to_unsigned(114,8) ,
57032	 => std_logic_vector(to_unsigned(108,8) ,
57033	 => std_logic_vector(to_unsigned(97,8) ,
57034	 => std_logic_vector(to_unsigned(109,8) ,
57035	 => std_logic_vector(to_unsigned(130,8) ,
57036	 => std_logic_vector(to_unsigned(130,8) ,
57037	 => std_logic_vector(to_unsigned(130,8) ,
57038	 => std_logic_vector(to_unsigned(136,8) ,
57039	 => std_logic_vector(to_unsigned(127,8) ,
57040	 => std_logic_vector(to_unsigned(121,8) ,
57041	 => std_logic_vector(to_unsigned(115,8) ,
57042	 => std_logic_vector(to_unsigned(81,8) ,
57043	 => std_logic_vector(to_unsigned(71,8) ,
57044	 => std_logic_vector(to_unsigned(97,8) ,
57045	 => std_logic_vector(to_unsigned(90,8) ,
57046	 => std_logic_vector(to_unsigned(44,8) ,
57047	 => std_logic_vector(to_unsigned(33,8) ,
57048	 => std_logic_vector(to_unsigned(34,8) ,
57049	 => std_logic_vector(to_unsigned(32,8) ,
57050	 => std_logic_vector(to_unsigned(34,8) ,
57051	 => std_logic_vector(to_unsigned(40,8) ,
57052	 => std_logic_vector(to_unsigned(40,8) ,
57053	 => std_logic_vector(to_unsigned(39,8) ,
57054	 => std_logic_vector(to_unsigned(46,8) ,
57055	 => std_logic_vector(to_unsigned(52,8) ,
57056	 => std_logic_vector(to_unsigned(58,8) ,
57057	 => std_logic_vector(to_unsigned(50,8) ,
57058	 => std_logic_vector(to_unsigned(45,8) ,
57059	 => std_logic_vector(to_unsigned(53,8) ,
57060	 => std_logic_vector(to_unsigned(51,8) ,
57061	 => std_logic_vector(to_unsigned(50,8) ,
57062	 => std_logic_vector(to_unsigned(54,8) ,
57063	 => std_logic_vector(to_unsigned(57,8) ,
57064	 => std_logic_vector(to_unsigned(58,8) ,
57065	 => std_logic_vector(to_unsigned(51,8) ,
57066	 => std_logic_vector(to_unsigned(59,8) ,
57067	 => std_logic_vector(to_unsigned(72,8) ,
57068	 => std_logic_vector(to_unsigned(79,8) ,
57069	 => std_logic_vector(to_unsigned(78,8) ,
57070	 => std_logic_vector(to_unsigned(93,8) ,
57071	 => std_logic_vector(to_unsigned(108,8) ,
57072	 => std_logic_vector(to_unsigned(115,8) ,
57073	 => std_logic_vector(to_unsigned(79,8) ,
57074	 => std_logic_vector(to_unsigned(53,8) ,
57075	 => std_logic_vector(to_unsigned(57,8) ,
57076	 => std_logic_vector(to_unsigned(76,8) ,
57077	 => std_logic_vector(to_unsigned(53,8) ,
57078	 => std_logic_vector(to_unsigned(63,8) ,
57079	 => std_logic_vector(to_unsigned(47,8) ,
57080	 => std_logic_vector(to_unsigned(30,8) ,
57081	 => std_logic_vector(to_unsigned(39,8) ,
57082	 => std_logic_vector(to_unsigned(48,8) ,
57083	 => std_logic_vector(to_unsigned(52,8) ,
57084	 => std_logic_vector(to_unsigned(63,8) ,
57085	 => std_logic_vector(to_unsigned(71,8) ,
57086	 => std_logic_vector(to_unsigned(66,8) ,
57087	 => std_logic_vector(to_unsigned(66,8) ,
57088	 => std_logic_vector(to_unsigned(61,8) ,
57089	 => std_logic_vector(to_unsigned(49,8) ,
57090	 => std_logic_vector(to_unsigned(37,8) ,
57091	 => std_logic_vector(to_unsigned(35,8) ,
57092	 => std_logic_vector(to_unsigned(39,8) ,
57093	 => std_logic_vector(to_unsigned(44,8) ,
57094	 => std_logic_vector(to_unsigned(41,8) ,
57095	 => std_logic_vector(to_unsigned(38,8) ,
57096	 => std_logic_vector(to_unsigned(41,8) ,
57097	 => std_logic_vector(to_unsigned(41,8) ,
57098	 => std_logic_vector(to_unsigned(44,8) ,
57099	 => std_logic_vector(to_unsigned(61,8) ,
57100	 => std_logic_vector(to_unsigned(49,8) ,
57101	 => std_logic_vector(to_unsigned(14,8) ,
57102	 => std_logic_vector(to_unsigned(9,8) ,
57103	 => std_logic_vector(to_unsigned(15,8) ,
57104	 => std_logic_vector(to_unsigned(12,8) ,
57105	 => std_logic_vector(to_unsigned(31,8) ,
57106	 => std_logic_vector(to_unsigned(41,8) ,
57107	 => std_logic_vector(to_unsigned(12,8) ,
57108	 => std_logic_vector(to_unsigned(7,8) ,
57109	 => std_logic_vector(to_unsigned(8,8) ,
57110	 => std_logic_vector(to_unsigned(53,8) ,
57111	 => std_logic_vector(to_unsigned(54,8) ,
57112	 => std_logic_vector(to_unsigned(53,8) ,
57113	 => std_logic_vector(to_unsigned(71,8) ,
57114	 => std_logic_vector(to_unsigned(77,8) ,
57115	 => std_logic_vector(to_unsigned(36,8) ,
57116	 => std_logic_vector(to_unsigned(45,8) ,
57117	 => std_logic_vector(to_unsigned(48,8) ,
57118	 => std_logic_vector(to_unsigned(6,8) ,
57119	 => std_logic_vector(to_unsigned(5,8) ,
57120	 => std_logic_vector(to_unsigned(8,8) ,
57121	 => std_logic_vector(to_unsigned(32,8) ,
57122	 => std_logic_vector(to_unsigned(36,8) ,
57123	 => std_logic_vector(to_unsigned(26,8) ,
57124	 => std_logic_vector(to_unsigned(28,8) ,
57125	 => std_logic_vector(to_unsigned(32,8) ,
57126	 => std_logic_vector(to_unsigned(43,8) ,
57127	 => std_logic_vector(to_unsigned(42,8) ,
57128	 => std_logic_vector(to_unsigned(37,8) ,
57129	 => std_logic_vector(to_unsigned(29,8) ,
57130	 => std_logic_vector(to_unsigned(24,8) ,
57131	 => std_logic_vector(to_unsigned(22,8) ,
57132	 => std_logic_vector(to_unsigned(22,8) ,
57133	 => std_logic_vector(to_unsigned(17,8) ,
57134	 => std_logic_vector(to_unsigned(11,8) ,
57135	 => std_logic_vector(to_unsigned(14,8) ,
57136	 => std_logic_vector(to_unsigned(17,8) ,
57137	 => std_logic_vector(to_unsigned(16,8) ,
57138	 => std_logic_vector(to_unsigned(22,8) ,
57139	 => std_logic_vector(to_unsigned(34,8) ,
57140	 => std_logic_vector(to_unsigned(43,8) ,
57141	 => std_logic_vector(to_unsigned(50,8) ,
57142	 => std_logic_vector(to_unsigned(48,8) ,
57143	 => std_logic_vector(to_unsigned(22,8) ,
57144	 => std_logic_vector(to_unsigned(19,8) ,
57145	 => std_logic_vector(to_unsigned(28,8) ,
57146	 => std_logic_vector(to_unsigned(25,8) ,
57147	 => std_logic_vector(to_unsigned(20,8) ,
57148	 => std_logic_vector(to_unsigned(26,8) ,
57149	 => std_logic_vector(to_unsigned(40,8) ,
57150	 => std_logic_vector(to_unsigned(56,8) ,
57151	 => std_logic_vector(to_unsigned(26,8) ,
57152	 => std_logic_vector(to_unsigned(18,8) ,
57153	 => std_logic_vector(to_unsigned(24,8) ,
57154	 => std_logic_vector(to_unsigned(20,8) ,
57155	 => std_logic_vector(to_unsigned(28,8) ,
57156	 => std_logic_vector(to_unsigned(30,8) ,
57157	 => std_logic_vector(to_unsigned(23,8) ,
57158	 => std_logic_vector(to_unsigned(23,8) ,
57159	 => std_logic_vector(to_unsigned(17,8) ,
57160	 => std_logic_vector(to_unsigned(22,8) ,
57161	 => std_logic_vector(to_unsigned(17,8) ,
57162	 => std_logic_vector(to_unsigned(12,8) ,
57163	 => std_logic_vector(to_unsigned(14,8) ,
57164	 => std_logic_vector(to_unsigned(29,8) ,
57165	 => std_logic_vector(to_unsigned(30,8) ,
57166	 => std_logic_vector(to_unsigned(9,8) ,
57167	 => std_logic_vector(to_unsigned(3,8) ,
57168	 => std_logic_vector(to_unsigned(8,8) ,
57169	 => std_logic_vector(to_unsigned(27,8) ,
57170	 => std_logic_vector(to_unsigned(25,8) ,
57171	 => std_logic_vector(to_unsigned(15,8) ,
57172	 => std_logic_vector(to_unsigned(11,8) ,
57173	 => std_logic_vector(to_unsigned(12,8) ,
57174	 => std_logic_vector(to_unsigned(17,8) ,
57175	 => std_logic_vector(to_unsigned(17,8) ,
57176	 => std_logic_vector(to_unsigned(16,8) ,
57177	 => std_logic_vector(to_unsigned(15,8) ,
57178	 => std_logic_vector(to_unsigned(11,8) ,
57179	 => std_logic_vector(to_unsigned(42,8) ,
57180	 => std_logic_vector(to_unsigned(130,8) ,
57181	 => std_logic_vector(to_unsigned(149,8) ,
57182	 => std_logic_vector(to_unsigned(138,8) ,
57183	 => std_logic_vector(to_unsigned(99,8) ,
57184	 => std_logic_vector(to_unsigned(30,8) ,
57185	 => std_logic_vector(to_unsigned(16,8) ,
57186	 => std_logic_vector(to_unsigned(10,8) ,
57187	 => std_logic_vector(to_unsigned(10,8) ,
57188	 => std_logic_vector(to_unsigned(14,8) ,
57189	 => std_logic_vector(to_unsigned(13,8) ,
57190	 => std_logic_vector(to_unsigned(7,8) ,
57191	 => std_logic_vector(to_unsigned(5,8) ,
57192	 => std_logic_vector(to_unsigned(9,8) ,
57193	 => std_logic_vector(to_unsigned(14,8) ,
57194	 => std_logic_vector(to_unsigned(17,8) ,
57195	 => std_logic_vector(to_unsigned(24,8) ,
57196	 => std_logic_vector(to_unsigned(24,8) ,
57197	 => std_logic_vector(to_unsigned(20,8) ,
57198	 => std_logic_vector(to_unsigned(24,8) ,
57199	 => std_logic_vector(to_unsigned(41,8) ,
57200	 => std_logic_vector(to_unsigned(41,8) ,
57201	 => std_logic_vector(to_unsigned(43,8) ,
57202	 => std_logic_vector(to_unsigned(25,8) ,
57203	 => std_logic_vector(to_unsigned(12,8) ,
57204	 => std_logic_vector(to_unsigned(13,8) ,
57205	 => std_logic_vector(to_unsigned(11,8) ,
57206	 => std_logic_vector(to_unsigned(12,8) ,
57207	 => std_logic_vector(to_unsigned(13,8) ,
57208	 => std_logic_vector(to_unsigned(11,8) ,
57209	 => std_logic_vector(to_unsigned(8,8) ,
57210	 => std_logic_vector(to_unsigned(9,8) ,
57211	 => std_logic_vector(to_unsigned(10,8) ,
57212	 => std_logic_vector(to_unsigned(10,8) ,
57213	 => std_logic_vector(to_unsigned(10,8) ,
57214	 => std_logic_vector(to_unsigned(11,8) ,
57215	 => std_logic_vector(to_unsigned(11,8) ,
57216	 => std_logic_vector(to_unsigned(13,8) ,
57217	 => std_logic_vector(to_unsigned(13,8) ,
57218	 => std_logic_vector(to_unsigned(14,8) ,
57219	 => std_logic_vector(to_unsigned(14,8) ,
57220	 => std_logic_vector(to_unsigned(12,8) ,
57221	 => std_logic_vector(to_unsigned(9,8) ,
57222	 => std_logic_vector(to_unsigned(1,8) ,
57223	 => std_logic_vector(to_unsigned(0,8) ,
57224	 => std_logic_vector(to_unsigned(6,8) ,
57225	 => std_logic_vector(to_unsigned(27,8) ,
57226	 => std_logic_vector(to_unsigned(27,8) ,
57227	 => std_logic_vector(to_unsigned(18,8) ,
57228	 => std_logic_vector(to_unsigned(13,8) ,
57229	 => std_logic_vector(to_unsigned(24,8) ,
57230	 => std_logic_vector(to_unsigned(32,8) ,
57231	 => std_logic_vector(to_unsigned(23,8) ,
57232	 => std_logic_vector(to_unsigned(16,8) ,
57233	 => std_logic_vector(to_unsigned(9,8) ,
57234	 => std_logic_vector(to_unsigned(7,8) ,
57235	 => std_logic_vector(to_unsigned(8,8) ,
57236	 => std_logic_vector(to_unsigned(7,8) ,
57237	 => std_logic_vector(to_unsigned(7,8) ,
57238	 => std_logic_vector(to_unsigned(8,8) ,
57239	 => std_logic_vector(to_unsigned(15,8) ,
57240	 => std_logic_vector(to_unsigned(21,8) ,
57241	 => std_logic_vector(to_unsigned(11,8) ,
57242	 => std_logic_vector(to_unsigned(1,8) ,
57243	 => std_logic_vector(to_unsigned(0,8) ,
57244	 => std_logic_vector(to_unsigned(0,8) ,
57245	 => std_logic_vector(to_unsigned(0,8) ,
57246	 => std_logic_vector(to_unsigned(1,8) ,
57247	 => std_logic_vector(to_unsigned(8,8) ,
57248	 => std_logic_vector(to_unsigned(5,8) ,
57249	 => std_logic_vector(to_unsigned(5,8) ,
57250	 => std_logic_vector(to_unsigned(13,8) ,
57251	 => std_logic_vector(to_unsigned(17,8) ,
57252	 => std_logic_vector(to_unsigned(13,8) ,
57253	 => std_logic_vector(to_unsigned(17,8) ,
57254	 => std_logic_vector(to_unsigned(15,8) ,
57255	 => std_logic_vector(to_unsigned(17,8) ,
57256	 => std_logic_vector(to_unsigned(17,8) ,
57257	 => std_logic_vector(to_unsigned(14,8) ,
57258	 => std_logic_vector(to_unsigned(11,8) ,
57259	 => std_logic_vector(to_unsigned(9,8) ,
57260	 => std_logic_vector(to_unsigned(9,8) ,
57261	 => std_logic_vector(to_unsigned(7,8) ,
57262	 => std_logic_vector(to_unsigned(8,8) ,
57263	 => std_logic_vector(to_unsigned(8,8) ,
57264	 => std_logic_vector(to_unsigned(7,8) ,
57265	 => std_logic_vector(to_unsigned(6,8) ,
57266	 => std_logic_vector(to_unsigned(4,8) ,
57267	 => std_logic_vector(to_unsigned(4,8) ,
57268	 => std_logic_vector(to_unsigned(6,8) ,
57269	 => std_logic_vector(to_unsigned(6,8) ,
57270	 => std_logic_vector(to_unsigned(8,8) ,
57271	 => std_logic_vector(to_unsigned(6,8) ,
57272	 => std_logic_vector(to_unsigned(10,8) ,
57273	 => std_logic_vector(to_unsigned(14,8) ,
57274	 => std_logic_vector(to_unsigned(12,8) ,
57275	 => std_logic_vector(to_unsigned(14,8) ,
57276	 => std_logic_vector(to_unsigned(14,8) ,
57277	 => std_logic_vector(to_unsigned(14,8) ,
57278	 => std_logic_vector(to_unsigned(17,8) ,
57279	 => std_logic_vector(to_unsigned(10,8) ,
57280	 => std_logic_vector(to_unsigned(7,8) ,
57281	 => std_logic_vector(to_unsigned(95,8) ,
57282	 => std_logic_vector(to_unsigned(82,8) ,
57283	 => std_logic_vector(to_unsigned(72,8) ,
57284	 => std_logic_vector(to_unsigned(72,8) ,
57285	 => std_logic_vector(to_unsigned(62,8) ,
57286	 => std_logic_vector(to_unsigned(37,8) ,
57287	 => std_logic_vector(to_unsigned(33,8) ,
57288	 => std_logic_vector(to_unsigned(55,8) ,
57289	 => std_logic_vector(to_unsigned(45,8) ,
57290	 => std_logic_vector(to_unsigned(77,8) ,
57291	 => std_logic_vector(to_unsigned(67,8) ,
57292	 => std_logic_vector(to_unsigned(37,8) ,
57293	 => std_logic_vector(to_unsigned(70,8) ,
57294	 => std_logic_vector(to_unsigned(95,8) ,
57295	 => std_logic_vector(to_unsigned(66,8) ,
57296	 => std_logic_vector(to_unsigned(66,8) ,
57297	 => std_logic_vector(to_unsigned(87,8) ,
57298	 => std_logic_vector(to_unsigned(63,8) ,
57299	 => std_logic_vector(to_unsigned(81,8) ,
57300	 => std_logic_vector(to_unsigned(87,8) ,
57301	 => std_logic_vector(to_unsigned(51,8) ,
57302	 => std_logic_vector(to_unsigned(38,8) ,
57303	 => std_logic_vector(to_unsigned(29,8) ,
57304	 => std_logic_vector(to_unsigned(67,8) ,
57305	 => std_logic_vector(to_unsigned(91,8) ,
57306	 => std_logic_vector(to_unsigned(68,8) ,
57307	 => std_logic_vector(to_unsigned(85,8) ,
57308	 => std_logic_vector(to_unsigned(58,8) ,
57309	 => std_logic_vector(to_unsigned(55,8) ,
57310	 => std_logic_vector(to_unsigned(73,8) ,
57311	 => std_logic_vector(to_unsigned(91,8) ,
57312	 => std_logic_vector(to_unsigned(73,8) ,
57313	 => std_logic_vector(to_unsigned(57,8) ,
57314	 => std_logic_vector(to_unsigned(23,8) ,
57315	 => std_logic_vector(to_unsigned(17,8) ,
57316	 => std_logic_vector(to_unsigned(27,8) ,
57317	 => std_logic_vector(to_unsigned(72,8) ,
57318	 => std_logic_vector(to_unsigned(46,8) ,
57319	 => std_logic_vector(to_unsigned(37,8) ,
57320	 => std_logic_vector(to_unsigned(51,8) ,
57321	 => std_logic_vector(to_unsigned(34,8) ,
57322	 => std_logic_vector(to_unsigned(25,8) ,
57323	 => std_logic_vector(to_unsigned(32,8) ,
57324	 => std_logic_vector(to_unsigned(38,8) ,
57325	 => std_logic_vector(to_unsigned(33,8) ,
57326	 => std_logic_vector(to_unsigned(50,8) ,
57327	 => std_logic_vector(to_unsigned(60,8) ,
57328	 => std_logic_vector(to_unsigned(59,8) ,
57329	 => std_logic_vector(to_unsigned(42,8) ,
57330	 => std_logic_vector(to_unsigned(43,8) ,
57331	 => std_logic_vector(to_unsigned(59,8) ,
57332	 => std_logic_vector(to_unsigned(68,8) ,
57333	 => std_logic_vector(to_unsigned(76,8) ,
57334	 => std_logic_vector(to_unsigned(74,8) ,
57335	 => std_logic_vector(to_unsigned(69,8) ,
57336	 => std_logic_vector(to_unsigned(65,8) ,
57337	 => std_logic_vector(to_unsigned(69,8) ,
57338	 => std_logic_vector(to_unsigned(67,8) ,
57339	 => std_logic_vector(to_unsigned(57,8) ,
57340	 => std_logic_vector(to_unsigned(58,8) ,
57341	 => std_logic_vector(to_unsigned(56,8) ,
57342	 => std_logic_vector(to_unsigned(60,8) ,
57343	 => std_logic_vector(to_unsigned(77,8) ,
57344	 => std_logic_vector(to_unsigned(84,8) ,
57345	 => std_logic_vector(to_unsigned(82,8) ,
57346	 => std_logic_vector(to_unsigned(84,8) ,
57347	 => std_logic_vector(to_unsigned(82,8) ,
57348	 => std_logic_vector(to_unsigned(87,8) ,
57349	 => std_logic_vector(to_unsigned(96,8) ,
57350	 => std_logic_vector(to_unsigned(90,8) ,
57351	 => std_logic_vector(to_unsigned(114,8) ,
57352	 => std_logic_vector(to_unsigned(105,8) ,
57353	 => std_logic_vector(to_unsigned(93,8) ,
57354	 => std_logic_vector(to_unsigned(134,8) ,
57355	 => std_logic_vector(to_unsigned(151,8) ,
57356	 => std_logic_vector(to_unsigned(138,8) ,
57357	 => std_logic_vector(to_unsigned(134,8) ,
57358	 => std_logic_vector(to_unsigned(125,8) ,
57359	 => std_logic_vector(to_unsigned(125,8) ,
57360	 => std_logic_vector(to_unsigned(125,8) ,
57361	 => std_logic_vector(to_unsigned(124,8) ,
57362	 => std_logic_vector(to_unsigned(101,8) ,
57363	 => std_logic_vector(to_unsigned(99,8) ,
57364	 => std_logic_vector(to_unsigned(112,8) ,
57365	 => std_logic_vector(to_unsigned(105,8) ,
57366	 => std_logic_vector(to_unsigned(66,8) ,
57367	 => std_logic_vector(to_unsigned(37,8) ,
57368	 => std_logic_vector(to_unsigned(36,8) ,
57369	 => std_logic_vector(to_unsigned(34,8) ,
57370	 => std_logic_vector(to_unsigned(37,8) ,
57371	 => std_logic_vector(to_unsigned(44,8) ,
57372	 => std_logic_vector(to_unsigned(43,8) ,
57373	 => std_logic_vector(to_unsigned(48,8) ,
57374	 => std_logic_vector(to_unsigned(47,8) ,
57375	 => std_logic_vector(to_unsigned(41,8) ,
57376	 => std_logic_vector(to_unsigned(50,8) ,
57377	 => std_logic_vector(to_unsigned(52,8) ,
57378	 => std_logic_vector(to_unsigned(47,8) ,
57379	 => std_logic_vector(to_unsigned(46,8) ,
57380	 => std_logic_vector(to_unsigned(47,8) ,
57381	 => std_logic_vector(to_unsigned(51,8) ,
57382	 => std_logic_vector(to_unsigned(54,8) ,
57383	 => std_logic_vector(to_unsigned(55,8) ,
57384	 => std_logic_vector(to_unsigned(51,8) ,
57385	 => std_logic_vector(to_unsigned(37,8) ,
57386	 => std_logic_vector(to_unsigned(35,8) ,
57387	 => std_logic_vector(to_unsigned(44,8) ,
57388	 => std_logic_vector(to_unsigned(40,8) ,
57389	 => std_logic_vector(to_unsigned(66,8) ,
57390	 => std_logic_vector(to_unsigned(114,8) ,
57391	 => std_logic_vector(to_unsigned(87,8) ,
57392	 => std_logic_vector(to_unsigned(91,8) ,
57393	 => std_logic_vector(to_unsigned(69,8) ,
57394	 => std_logic_vector(to_unsigned(54,8) ,
57395	 => std_logic_vector(to_unsigned(63,8) ,
57396	 => std_logic_vector(to_unsigned(79,8) ,
57397	 => std_logic_vector(to_unsigned(54,8) ,
57398	 => std_logic_vector(to_unsigned(61,8) ,
57399	 => std_logic_vector(to_unsigned(45,8) ,
57400	 => std_logic_vector(to_unsigned(41,8) ,
57401	 => std_logic_vector(to_unsigned(51,8) ,
57402	 => std_logic_vector(to_unsigned(41,8) ,
57403	 => std_logic_vector(to_unsigned(45,8) ,
57404	 => std_logic_vector(to_unsigned(54,8) ,
57405	 => std_logic_vector(to_unsigned(68,8) ,
57406	 => std_logic_vector(to_unsigned(64,8) ,
57407	 => std_logic_vector(to_unsigned(62,8) ,
57408	 => std_logic_vector(to_unsigned(55,8) ,
57409	 => std_logic_vector(to_unsigned(49,8) ,
57410	 => std_logic_vector(to_unsigned(51,8) ,
57411	 => std_logic_vector(to_unsigned(49,8) ,
57412	 => std_logic_vector(to_unsigned(48,8) ,
57413	 => std_logic_vector(to_unsigned(44,8) ,
57414	 => std_logic_vector(to_unsigned(43,8) ,
57415	 => std_logic_vector(to_unsigned(47,8) ,
57416	 => std_logic_vector(to_unsigned(44,8) ,
57417	 => std_logic_vector(to_unsigned(51,8) ,
57418	 => std_logic_vector(to_unsigned(63,8) ,
57419	 => std_logic_vector(to_unsigned(35,8) ,
57420	 => std_logic_vector(to_unsigned(13,8) ,
57421	 => std_logic_vector(to_unsigned(11,8) ,
57422	 => std_logic_vector(to_unsigned(15,8) ,
57423	 => std_logic_vector(to_unsigned(13,8) ,
57424	 => std_logic_vector(to_unsigned(10,8) ,
57425	 => std_logic_vector(to_unsigned(25,8) ,
57426	 => std_logic_vector(to_unsigned(45,8) ,
57427	 => std_logic_vector(to_unsigned(42,8) ,
57428	 => std_logic_vector(to_unsigned(38,8) ,
57429	 => std_logic_vector(to_unsigned(30,8) ,
57430	 => std_logic_vector(to_unsigned(51,8) ,
57431	 => std_logic_vector(to_unsigned(30,8) ,
57432	 => std_logic_vector(to_unsigned(37,8) ,
57433	 => std_logic_vector(to_unsigned(65,8) ,
57434	 => std_logic_vector(to_unsigned(65,8) ,
57435	 => std_logic_vector(to_unsigned(29,8) ,
57436	 => std_logic_vector(to_unsigned(28,8) ,
57437	 => std_logic_vector(to_unsigned(42,8) ,
57438	 => std_logic_vector(to_unsigned(7,8) ,
57439	 => std_logic_vector(to_unsigned(4,8) ,
57440	 => std_logic_vector(to_unsigned(20,8) ,
57441	 => std_logic_vector(to_unsigned(111,8) ,
57442	 => std_logic_vector(to_unsigned(88,8) ,
57443	 => std_logic_vector(to_unsigned(64,8) ,
57444	 => std_logic_vector(to_unsigned(49,8) ,
57445	 => std_logic_vector(to_unsigned(51,8) ,
57446	 => std_logic_vector(to_unsigned(105,8) ,
57447	 => std_logic_vector(to_unsigned(43,8) ,
57448	 => std_logic_vector(to_unsigned(22,8) ,
57449	 => std_logic_vector(to_unsigned(35,8) ,
57450	 => std_logic_vector(to_unsigned(33,8) ,
57451	 => std_logic_vector(to_unsigned(32,8) ,
57452	 => std_logic_vector(to_unsigned(27,8) ,
57453	 => std_logic_vector(to_unsigned(20,8) ,
57454	 => std_logic_vector(to_unsigned(12,8) ,
57455	 => std_logic_vector(to_unsigned(10,8) ,
57456	 => std_logic_vector(to_unsigned(9,8) ,
57457	 => std_logic_vector(to_unsigned(8,8) ,
57458	 => std_logic_vector(to_unsigned(10,8) ,
57459	 => std_logic_vector(to_unsigned(9,8) ,
57460	 => std_logic_vector(to_unsigned(15,8) ,
57461	 => std_logic_vector(to_unsigned(28,8) ,
57462	 => std_logic_vector(to_unsigned(44,8) ,
57463	 => std_logic_vector(to_unsigned(21,8) ,
57464	 => std_logic_vector(to_unsigned(22,8) ,
57465	 => std_logic_vector(to_unsigned(41,8) ,
57466	 => std_logic_vector(to_unsigned(38,8) ,
57467	 => std_logic_vector(to_unsigned(41,8) ,
57468	 => std_logic_vector(to_unsigned(53,8) ,
57469	 => std_logic_vector(to_unsigned(58,8) ,
57470	 => std_logic_vector(to_unsigned(30,8) ,
57471	 => std_logic_vector(to_unsigned(16,8) ,
57472	 => std_logic_vector(to_unsigned(17,8) ,
57473	 => std_logic_vector(to_unsigned(35,8) ,
57474	 => std_logic_vector(to_unsigned(40,8) ,
57475	 => std_logic_vector(to_unsigned(37,8) ,
57476	 => std_logic_vector(to_unsigned(30,8) ,
57477	 => std_logic_vector(to_unsigned(15,8) ,
57478	 => std_logic_vector(to_unsigned(18,8) ,
57479	 => std_logic_vector(to_unsigned(19,8) ,
57480	 => std_logic_vector(to_unsigned(16,8) ,
57481	 => std_logic_vector(to_unsigned(26,8) ,
57482	 => std_logic_vector(to_unsigned(37,8) ,
57483	 => std_logic_vector(to_unsigned(32,8) ,
57484	 => std_logic_vector(to_unsigned(29,8) ,
57485	 => std_logic_vector(to_unsigned(33,8) ,
57486	 => std_logic_vector(to_unsigned(25,8) ,
57487	 => std_logic_vector(to_unsigned(15,8) ,
57488	 => std_logic_vector(to_unsigned(13,8) ,
57489	 => std_logic_vector(to_unsigned(24,8) ,
57490	 => std_logic_vector(to_unsigned(23,8) ,
57491	 => std_logic_vector(to_unsigned(13,8) ,
57492	 => std_logic_vector(to_unsigned(6,8) ,
57493	 => std_logic_vector(to_unsigned(6,8) ,
57494	 => std_logic_vector(to_unsigned(14,8) ,
57495	 => std_logic_vector(to_unsigned(9,8) ,
57496	 => std_logic_vector(to_unsigned(4,8) ,
57497	 => std_logic_vector(to_unsigned(8,8) ,
57498	 => std_logic_vector(to_unsigned(10,8) ,
57499	 => std_logic_vector(to_unsigned(4,8) ,
57500	 => std_logic_vector(to_unsigned(18,8) ,
57501	 => std_logic_vector(to_unsigned(82,8) ,
57502	 => std_logic_vector(to_unsigned(144,8) ,
57503	 => std_logic_vector(to_unsigned(58,8) ,
57504	 => std_logic_vector(to_unsigned(11,8) ,
57505	 => std_logic_vector(to_unsigned(22,8) ,
57506	 => std_logic_vector(to_unsigned(13,8) ,
57507	 => std_logic_vector(to_unsigned(13,8) ,
57508	 => std_logic_vector(to_unsigned(17,8) ,
57509	 => std_logic_vector(to_unsigned(15,8) ,
57510	 => std_logic_vector(to_unsigned(12,8) ,
57511	 => std_logic_vector(to_unsigned(8,8) ,
57512	 => std_logic_vector(to_unsigned(7,8) ,
57513	 => std_logic_vector(to_unsigned(11,8) ,
57514	 => std_logic_vector(to_unsigned(22,8) ,
57515	 => std_logic_vector(to_unsigned(21,8) ,
57516	 => std_logic_vector(to_unsigned(17,8) ,
57517	 => std_logic_vector(to_unsigned(9,8) ,
57518	 => std_logic_vector(to_unsigned(9,8) ,
57519	 => std_logic_vector(to_unsigned(29,8) ,
57520	 => std_logic_vector(to_unsigned(27,8) ,
57521	 => std_logic_vector(to_unsigned(28,8) ,
57522	 => std_logic_vector(to_unsigned(22,8) ,
57523	 => std_logic_vector(to_unsigned(17,8) ,
57524	 => std_logic_vector(to_unsigned(28,8) ,
57525	 => std_logic_vector(to_unsigned(28,8) ,
57526	 => std_logic_vector(to_unsigned(17,8) ,
57527	 => std_logic_vector(to_unsigned(12,8) ,
57528	 => std_logic_vector(to_unsigned(12,8) ,
57529	 => std_logic_vector(to_unsigned(9,8) ,
57530	 => std_logic_vector(to_unsigned(10,8) ,
57531	 => std_logic_vector(to_unsigned(13,8) ,
57532	 => std_logic_vector(to_unsigned(11,8) ,
57533	 => std_logic_vector(to_unsigned(10,8) ,
57534	 => std_logic_vector(to_unsigned(10,8) ,
57535	 => std_logic_vector(to_unsigned(10,8) ,
57536	 => std_logic_vector(to_unsigned(10,8) ,
57537	 => std_logic_vector(to_unsigned(11,8) ,
57538	 => std_logic_vector(to_unsigned(13,8) ,
57539	 => std_logic_vector(to_unsigned(12,8) ,
57540	 => std_logic_vector(to_unsigned(13,8) ,
57541	 => std_logic_vector(to_unsigned(11,8) ,
57542	 => std_logic_vector(to_unsigned(1,8) ,
57543	 => std_logic_vector(to_unsigned(0,8) ,
57544	 => std_logic_vector(to_unsigned(2,8) ,
57545	 => std_logic_vector(to_unsigned(22,8) ,
57546	 => std_logic_vector(to_unsigned(23,8) ,
57547	 => std_logic_vector(to_unsigned(17,8) ,
57548	 => std_logic_vector(to_unsigned(13,8) ,
57549	 => std_logic_vector(to_unsigned(19,8) ,
57550	 => std_logic_vector(to_unsigned(23,8) ,
57551	 => std_logic_vector(to_unsigned(18,8) ,
57552	 => std_logic_vector(to_unsigned(12,8) ,
57553	 => std_logic_vector(to_unsigned(13,8) ,
57554	 => std_logic_vector(to_unsigned(13,8) ,
57555	 => std_logic_vector(to_unsigned(9,8) ,
57556	 => std_logic_vector(to_unsigned(8,8) ,
57557	 => std_logic_vector(to_unsigned(9,8) ,
57558	 => std_logic_vector(to_unsigned(10,8) ,
57559	 => std_logic_vector(to_unsigned(16,8) ,
57560	 => std_logic_vector(to_unsigned(13,8) ,
57561	 => std_logic_vector(to_unsigned(10,8) ,
57562	 => std_logic_vector(to_unsigned(3,8) ,
57563	 => std_logic_vector(to_unsigned(0,8) ,
57564	 => std_logic_vector(to_unsigned(0,8) ,
57565	 => std_logic_vector(to_unsigned(0,8) ,
57566	 => std_logic_vector(to_unsigned(0,8) ,
57567	 => std_logic_vector(to_unsigned(3,8) ,
57568	 => std_logic_vector(to_unsigned(10,8) ,
57569	 => std_logic_vector(to_unsigned(5,8) ,
57570	 => std_logic_vector(to_unsigned(7,8) ,
57571	 => std_logic_vector(to_unsigned(10,8) ,
57572	 => std_logic_vector(to_unsigned(9,8) ,
57573	 => std_logic_vector(to_unsigned(10,8) ,
57574	 => std_logic_vector(to_unsigned(14,8) ,
57575	 => std_logic_vector(to_unsigned(19,8) ,
57576	 => std_logic_vector(to_unsigned(15,8) ,
57577	 => std_logic_vector(to_unsigned(14,8) ,
57578	 => std_logic_vector(to_unsigned(16,8) ,
57579	 => std_logic_vector(to_unsigned(13,8) ,
57580	 => std_logic_vector(to_unsigned(20,8) ,
57581	 => std_logic_vector(to_unsigned(19,8) ,
57582	 => std_logic_vector(to_unsigned(17,8) ,
57583	 => std_logic_vector(to_unsigned(17,8) ,
57584	 => std_logic_vector(to_unsigned(14,8) ,
57585	 => std_logic_vector(to_unsigned(8,8) ,
57586	 => std_logic_vector(to_unsigned(9,8) ,
57587	 => std_logic_vector(to_unsigned(9,8) ,
57588	 => std_logic_vector(to_unsigned(7,8) ,
57589	 => std_logic_vector(to_unsigned(4,8) ,
57590	 => std_logic_vector(to_unsigned(8,8) ,
57591	 => std_logic_vector(to_unsigned(12,8) ,
57592	 => std_logic_vector(to_unsigned(11,8) ,
57593	 => std_logic_vector(to_unsigned(12,8) ,
57594	 => std_logic_vector(to_unsigned(21,8) ,
57595	 => std_logic_vector(to_unsigned(35,8) ,
57596	 => std_logic_vector(to_unsigned(35,8) ,
57597	 => std_logic_vector(to_unsigned(22,8) ,
57598	 => std_logic_vector(to_unsigned(10,8) ,
57599	 => std_logic_vector(to_unsigned(7,8) ,
57600	 => std_logic_vector(to_unsigned(9,8) ,
57601	 => std_logic_vector(to_unsigned(84,8) ,
57602	 => std_logic_vector(to_unsigned(96,8) ,
57603	 => std_logic_vector(to_unsigned(101,8) ,
57604	 => std_logic_vector(to_unsigned(72,8) ,
57605	 => std_logic_vector(to_unsigned(55,8) ,
57606	 => std_logic_vector(to_unsigned(37,8) ,
57607	 => std_logic_vector(to_unsigned(25,8) ,
57608	 => std_logic_vector(to_unsigned(64,8) ,
57609	 => std_logic_vector(to_unsigned(87,8) ,
57610	 => std_logic_vector(to_unsigned(71,8) ,
57611	 => std_logic_vector(to_unsigned(62,8) ,
57612	 => std_logic_vector(to_unsigned(58,8) ,
57613	 => std_logic_vector(to_unsigned(74,8) ,
57614	 => std_logic_vector(to_unsigned(87,8) ,
57615	 => std_logic_vector(to_unsigned(92,8) ,
57616	 => std_logic_vector(to_unsigned(128,8) ,
57617	 => std_logic_vector(to_unsigned(93,8) ,
57618	 => std_logic_vector(to_unsigned(57,8) ,
57619	 => std_logic_vector(to_unsigned(55,8) ,
57620	 => std_logic_vector(to_unsigned(71,8) ,
57621	 => std_logic_vector(to_unsigned(32,8) ,
57622	 => std_logic_vector(to_unsigned(26,8) ,
57623	 => std_logic_vector(to_unsigned(32,8) ,
57624	 => std_logic_vector(to_unsigned(70,8) ,
57625	 => std_logic_vector(to_unsigned(97,8) ,
57626	 => std_logic_vector(to_unsigned(72,8) ,
57627	 => std_logic_vector(to_unsigned(92,8) ,
57628	 => std_logic_vector(to_unsigned(74,8) ,
57629	 => std_logic_vector(to_unsigned(65,8) ,
57630	 => std_logic_vector(to_unsigned(70,8) ,
57631	 => std_logic_vector(to_unsigned(96,8) ,
57632	 => std_logic_vector(to_unsigned(73,8) ,
57633	 => std_logic_vector(to_unsigned(53,8) ,
57634	 => std_logic_vector(to_unsigned(22,8) ,
57635	 => std_logic_vector(to_unsigned(16,8) ,
57636	 => std_logic_vector(to_unsigned(24,8) ,
57637	 => std_logic_vector(to_unsigned(64,8) ,
57638	 => std_logic_vector(to_unsigned(79,8) ,
57639	 => std_logic_vector(to_unsigned(69,8) ,
57640	 => std_logic_vector(to_unsigned(41,8) ,
57641	 => std_logic_vector(to_unsigned(29,8) ,
57642	 => std_logic_vector(to_unsigned(26,8) ,
57643	 => std_logic_vector(to_unsigned(26,8) ,
57644	 => std_logic_vector(to_unsigned(29,8) ,
57645	 => std_logic_vector(to_unsigned(26,8) ,
57646	 => std_logic_vector(to_unsigned(36,8) ,
57647	 => std_logic_vector(to_unsigned(47,8) ,
57648	 => std_logic_vector(to_unsigned(63,8) ,
57649	 => std_logic_vector(to_unsigned(51,8) ,
57650	 => std_logic_vector(to_unsigned(51,8) ,
57651	 => std_logic_vector(to_unsigned(59,8) ,
57652	 => std_logic_vector(to_unsigned(72,8) ,
57653	 => std_logic_vector(to_unsigned(69,8) ,
57654	 => std_logic_vector(to_unsigned(59,8) ,
57655	 => std_logic_vector(to_unsigned(69,8) ,
57656	 => std_logic_vector(to_unsigned(73,8) ,
57657	 => std_logic_vector(to_unsigned(68,8) ,
57658	 => std_logic_vector(to_unsigned(53,8) ,
57659	 => std_logic_vector(to_unsigned(70,8) ,
57660	 => std_logic_vector(to_unsigned(63,8) ,
57661	 => std_logic_vector(to_unsigned(44,8) ,
57662	 => std_logic_vector(to_unsigned(39,8) ,
57663	 => std_logic_vector(to_unsigned(74,8) ,
57664	 => std_logic_vector(to_unsigned(81,8) ,
57665	 => std_logic_vector(to_unsigned(82,8) ,
57666	 => std_logic_vector(to_unsigned(90,8) ,
57667	 => std_logic_vector(to_unsigned(86,8) ,
57668	 => std_logic_vector(to_unsigned(87,8) ,
57669	 => std_logic_vector(to_unsigned(90,8) ,
57670	 => std_logic_vector(to_unsigned(92,8) ,
57671	 => std_logic_vector(to_unsigned(97,8) ,
57672	 => std_logic_vector(to_unsigned(90,8) ,
57673	 => std_logic_vector(to_unsigned(87,8) ,
57674	 => std_logic_vector(to_unsigned(133,8) ,
57675	 => std_logic_vector(to_unsigned(151,8) ,
57676	 => std_logic_vector(to_unsigned(131,8) ,
57677	 => std_logic_vector(to_unsigned(133,8) ,
57678	 => std_logic_vector(to_unsigned(131,8) ,
57679	 => std_logic_vector(to_unsigned(131,8) ,
57680	 => std_logic_vector(to_unsigned(127,8) ,
57681	 => std_logic_vector(to_unsigned(115,8) ,
57682	 => std_logic_vector(to_unsigned(100,8) ,
57683	 => std_logic_vector(to_unsigned(118,8) ,
57684	 => std_logic_vector(to_unsigned(116,8) ,
57685	 => std_logic_vector(to_unsigned(97,8) ,
57686	 => std_logic_vector(to_unsigned(64,8) ,
57687	 => std_logic_vector(to_unsigned(37,8) ,
57688	 => std_logic_vector(to_unsigned(40,8) ,
57689	 => std_logic_vector(to_unsigned(41,8) ,
57690	 => std_logic_vector(to_unsigned(44,8) ,
57691	 => std_logic_vector(to_unsigned(44,8) ,
57692	 => std_logic_vector(to_unsigned(53,8) ,
57693	 => std_logic_vector(to_unsigned(63,8) ,
57694	 => std_logic_vector(to_unsigned(60,8) ,
57695	 => std_logic_vector(to_unsigned(64,8) ,
57696	 => std_logic_vector(to_unsigned(58,8) ,
57697	 => std_logic_vector(to_unsigned(48,8) ,
57698	 => std_logic_vector(to_unsigned(36,8) ,
57699	 => std_logic_vector(to_unsigned(43,8) ,
57700	 => std_logic_vector(to_unsigned(50,8) ,
57701	 => std_logic_vector(to_unsigned(47,8) ,
57702	 => std_logic_vector(to_unsigned(50,8) ,
57703	 => std_logic_vector(to_unsigned(52,8) ,
57704	 => std_logic_vector(to_unsigned(51,8) ,
57705	 => std_logic_vector(to_unsigned(43,8) ,
57706	 => std_logic_vector(to_unsigned(35,8) ,
57707	 => std_logic_vector(to_unsigned(35,8) ,
57708	 => std_logic_vector(to_unsigned(27,8) ,
57709	 => std_logic_vector(to_unsigned(60,8) ,
57710	 => std_logic_vector(to_unsigned(104,8) ,
57711	 => std_logic_vector(to_unsigned(61,8) ,
57712	 => std_logic_vector(to_unsigned(84,8) ,
57713	 => std_logic_vector(to_unsigned(76,8) ,
57714	 => std_logic_vector(to_unsigned(59,8) ,
57715	 => std_logic_vector(to_unsigned(65,8) ,
57716	 => std_logic_vector(to_unsigned(82,8) ,
57717	 => std_logic_vector(to_unsigned(53,8) ,
57718	 => std_logic_vector(to_unsigned(58,8) ,
57719	 => std_logic_vector(to_unsigned(53,8) ,
57720	 => std_logic_vector(to_unsigned(37,8) ,
57721	 => std_logic_vector(to_unsigned(52,8) ,
57722	 => std_logic_vector(to_unsigned(49,8) ,
57723	 => std_logic_vector(to_unsigned(53,8) ,
57724	 => std_logic_vector(to_unsigned(62,8) ,
57725	 => std_logic_vector(to_unsigned(61,8) ,
57726	 => std_logic_vector(to_unsigned(41,8) ,
57727	 => std_logic_vector(to_unsigned(54,8) ,
57728	 => std_logic_vector(to_unsigned(56,8) ,
57729	 => std_logic_vector(to_unsigned(51,8) ,
57730	 => std_logic_vector(to_unsigned(41,8) ,
57731	 => std_logic_vector(to_unsigned(43,8) ,
57732	 => std_logic_vector(to_unsigned(50,8) ,
57733	 => std_logic_vector(to_unsigned(44,8) ,
57734	 => std_logic_vector(to_unsigned(46,8) ,
57735	 => std_logic_vector(to_unsigned(51,8) ,
57736	 => std_logic_vector(to_unsigned(58,8) ,
57737	 => std_logic_vector(to_unsigned(60,8) ,
57738	 => std_logic_vector(to_unsigned(29,8) ,
57739	 => std_logic_vector(to_unsigned(12,8) ,
57740	 => std_logic_vector(to_unsigned(17,8) ,
57741	 => std_logic_vector(to_unsigned(16,8) ,
57742	 => std_logic_vector(to_unsigned(13,8) ,
57743	 => std_logic_vector(to_unsigned(12,8) ,
57744	 => std_logic_vector(to_unsigned(11,8) ,
57745	 => std_logic_vector(to_unsigned(25,8) ,
57746	 => std_logic_vector(to_unsigned(55,8) ,
57747	 => std_logic_vector(to_unsigned(38,8) ,
57748	 => std_logic_vector(to_unsigned(36,8) ,
57749	 => std_logic_vector(to_unsigned(71,8) ,
57750	 => std_logic_vector(to_unsigned(73,8) ,
57751	 => std_logic_vector(to_unsigned(36,8) ,
57752	 => std_logic_vector(to_unsigned(33,8) ,
57753	 => std_logic_vector(to_unsigned(64,8) ,
57754	 => std_logic_vector(to_unsigned(76,8) ,
57755	 => std_logic_vector(to_unsigned(35,8) ,
57756	 => std_logic_vector(to_unsigned(31,8) ,
57757	 => std_logic_vector(to_unsigned(50,8) ,
57758	 => std_logic_vector(to_unsigned(14,8) ,
57759	 => std_logic_vector(to_unsigned(8,8) ,
57760	 => std_logic_vector(to_unsigned(29,8) ,
57761	 => std_logic_vector(to_unsigned(149,8) ,
57762	 => std_logic_vector(to_unsigned(163,8) ,
57763	 => std_logic_vector(to_unsigned(161,8) ,
57764	 => std_logic_vector(to_unsigned(136,8) ,
57765	 => std_logic_vector(to_unsigned(146,8) ,
57766	 => std_logic_vector(to_unsigned(142,8) ,
57767	 => std_logic_vector(to_unsigned(23,8) ,
57768	 => std_logic_vector(to_unsigned(6,8) ,
57769	 => std_logic_vector(to_unsigned(12,8) ,
57770	 => std_logic_vector(to_unsigned(13,8) ,
57771	 => std_logic_vector(to_unsigned(12,8) ,
57772	 => std_logic_vector(to_unsigned(16,8) ,
57773	 => std_logic_vector(to_unsigned(19,8) ,
57774	 => std_logic_vector(to_unsigned(18,8) ,
57775	 => std_logic_vector(to_unsigned(15,8) ,
57776	 => std_logic_vector(to_unsigned(17,8) ,
57777	 => std_logic_vector(to_unsigned(18,8) ,
57778	 => std_logic_vector(to_unsigned(21,8) ,
57779	 => std_logic_vector(to_unsigned(16,8) ,
57780	 => std_logic_vector(to_unsigned(18,8) ,
57781	 => std_logic_vector(to_unsigned(21,8) ,
57782	 => std_logic_vector(to_unsigned(44,8) ,
57783	 => std_logic_vector(to_unsigned(44,8) ,
57784	 => std_logic_vector(to_unsigned(41,8) ,
57785	 => std_logic_vector(to_unsigned(51,8) ,
57786	 => std_logic_vector(to_unsigned(51,8) ,
57787	 => std_logic_vector(to_unsigned(56,8) ,
57788	 => std_logic_vector(to_unsigned(65,8) ,
57789	 => std_logic_vector(to_unsigned(40,8) ,
57790	 => std_logic_vector(to_unsigned(14,8) ,
57791	 => std_logic_vector(to_unsigned(23,8) ,
57792	 => std_logic_vector(to_unsigned(20,8) ,
57793	 => std_logic_vector(to_unsigned(23,8) ,
57794	 => std_logic_vector(to_unsigned(35,8) ,
57795	 => std_logic_vector(to_unsigned(23,8) ,
57796	 => std_logic_vector(to_unsigned(18,8) ,
57797	 => std_logic_vector(to_unsigned(22,8) ,
57798	 => std_logic_vector(to_unsigned(33,8) ,
57799	 => std_logic_vector(to_unsigned(29,8) ,
57800	 => std_logic_vector(to_unsigned(19,8) ,
57801	 => std_logic_vector(to_unsigned(23,8) ,
57802	 => std_logic_vector(to_unsigned(28,8) ,
57803	 => std_logic_vector(to_unsigned(29,8) ,
57804	 => std_logic_vector(to_unsigned(29,8) ,
57805	 => std_logic_vector(to_unsigned(29,8) ,
57806	 => std_logic_vector(to_unsigned(34,8) ,
57807	 => std_logic_vector(to_unsigned(44,8) ,
57808	 => std_logic_vector(to_unsigned(36,8) ,
57809	 => std_logic_vector(to_unsigned(24,8) ,
57810	 => std_logic_vector(to_unsigned(21,8) ,
57811	 => std_logic_vector(to_unsigned(24,8) ,
57812	 => std_logic_vector(to_unsigned(25,8) ,
57813	 => std_logic_vector(to_unsigned(17,8) ,
57814	 => std_logic_vector(to_unsigned(14,8) ,
57815	 => std_logic_vector(to_unsigned(11,8) ,
57816	 => std_logic_vector(to_unsigned(8,8) ,
57817	 => std_logic_vector(to_unsigned(11,8) ,
57818	 => std_logic_vector(to_unsigned(12,8) ,
57819	 => std_logic_vector(to_unsigned(5,8) ,
57820	 => std_logic_vector(to_unsigned(1,8) ,
57821	 => std_logic_vector(to_unsigned(6,8) ,
57822	 => std_logic_vector(to_unsigned(37,8) ,
57823	 => std_logic_vector(to_unsigned(23,8) ,
57824	 => std_logic_vector(to_unsigned(18,8) ,
57825	 => std_logic_vector(to_unsigned(28,8) ,
57826	 => std_logic_vector(to_unsigned(22,8) ,
57827	 => std_logic_vector(to_unsigned(21,8) ,
57828	 => std_logic_vector(to_unsigned(14,8) ,
57829	 => std_logic_vector(to_unsigned(12,8) ,
57830	 => std_logic_vector(to_unsigned(12,8) ,
57831	 => std_logic_vector(to_unsigned(12,8) ,
57832	 => std_logic_vector(to_unsigned(14,8) ,
57833	 => std_logic_vector(to_unsigned(17,8) ,
57834	 => std_logic_vector(to_unsigned(18,8) ,
57835	 => std_logic_vector(to_unsigned(13,8) ,
57836	 => std_logic_vector(to_unsigned(8,8) ,
57837	 => std_logic_vector(to_unsigned(5,8) ,
57838	 => std_logic_vector(to_unsigned(12,8) ,
57839	 => std_logic_vector(to_unsigned(43,8) ,
57840	 => std_logic_vector(to_unsigned(41,8) ,
57841	 => std_logic_vector(to_unsigned(32,8) ,
57842	 => std_logic_vector(to_unsigned(20,8) ,
57843	 => std_logic_vector(to_unsigned(30,8) ,
57844	 => std_logic_vector(to_unsigned(41,8) ,
57845	 => std_logic_vector(to_unsigned(43,8) ,
57846	 => std_logic_vector(to_unsigned(25,8) ,
57847	 => std_logic_vector(to_unsigned(13,8) ,
57848	 => std_logic_vector(to_unsigned(24,8) ,
57849	 => std_logic_vector(to_unsigned(11,8) ,
57850	 => std_logic_vector(to_unsigned(8,8) ,
57851	 => std_logic_vector(to_unsigned(12,8) ,
57852	 => std_logic_vector(to_unsigned(12,8) ,
57853	 => std_logic_vector(to_unsigned(9,8) ,
57854	 => std_logic_vector(to_unsigned(9,8) ,
57855	 => std_logic_vector(to_unsigned(8,8) ,
57856	 => std_logic_vector(to_unsigned(8,8) ,
57857	 => std_logic_vector(to_unsigned(8,8) ,
57858	 => std_logic_vector(to_unsigned(9,8) ,
57859	 => std_logic_vector(to_unsigned(13,8) ,
57860	 => std_logic_vector(to_unsigned(14,8) ,
57861	 => std_logic_vector(to_unsigned(8,8) ,
57862	 => std_logic_vector(to_unsigned(2,8) ,
57863	 => std_logic_vector(to_unsigned(0,8) ,
57864	 => std_logic_vector(to_unsigned(1,8) ,
57865	 => std_logic_vector(to_unsigned(12,8) ,
57866	 => std_logic_vector(to_unsigned(19,8) ,
57867	 => std_logic_vector(to_unsigned(14,8) ,
57868	 => std_logic_vector(to_unsigned(23,8) ,
57869	 => std_logic_vector(to_unsigned(27,8) ,
57870	 => std_logic_vector(to_unsigned(25,8) ,
57871	 => std_logic_vector(to_unsigned(29,8) ,
57872	 => std_logic_vector(to_unsigned(22,8) ,
57873	 => std_logic_vector(to_unsigned(16,8) ,
57874	 => std_logic_vector(to_unsigned(12,8) ,
57875	 => std_logic_vector(to_unsigned(6,8) ,
57876	 => std_logic_vector(to_unsigned(9,8) ,
57877	 => std_logic_vector(to_unsigned(9,8) ,
57878	 => std_logic_vector(to_unsigned(10,8) ,
57879	 => std_logic_vector(to_unsigned(15,8) ,
57880	 => std_logic_vector(to_unsigned(8,8) ,
57881	 => std_logic_vector(to_unsigned(5,8) ,
57882	 => std_logic_vector(to_unsigned(4,8) ,
57883	 => std_logic_vector(to_unsigned(1,8) ,
57884	 => std_logic_vector(to_unsigned(0,8) ,
57885	 => std_logic_vector(to_unsigned(0,8) ,
57886	 => std_logic_vector(to_unsigned(0,8) ,
57887	 => std_logic_vector(to_unsigned(4,8) ,
57888	 => std_logic_vector(to_unsigned(6,8) ,
57889	 => std_logic_vector(to_unsigned(2,8) ,
57890	 => std_logic_vector(to_unsigned(2,8) ,
57891	 => std_logic_vector(to_unsigned(1,8) ,
57892	 => std_logic_vector(to_unsigned(1,8) ,
57893	 => std_logic_vector(to_unsigned(3,8) ,
57894	 => std_logic_vector(to_unsigned(11,8) ,
57895	 => std_logic_vector(to_unsigned(15,8) ,
57896	 => std_logic_vector(to_unsigned(8,8) ,
57897	 => std_logic_vector(to_unsigned(8,8) ,
57898	 => std_logic_vector(to_unsigned(15,8) ,
57899	 => std_logic_vector(to_unsigned(19,8) ,
57900	 => std_logic_vector(to_unsigned(22,8) ,
57901	 => std_logic_vector(to_unsigned(25,8) ,
57902	 => std_logic_vector(to_unsigned(35,8) ,
57903	 => std_logic_vector(to_unsigned(30,8) ,
57904	 => std_logic_vector(to_unsigned(24,8) ,
57905	 => std_logic_vector(to_unsigned(23,8) ,
57906	 => std_logic_vector(to_unsigned(13,8) ,
57907	 => std_logic_vector(to_unsigned(10,8) ,
57908	 => std_logic_vector(to_unsigned(9,8) ,
57909	 => std_logic_vector(to_unsigned(5,8) ,
57910	 => std_logic_vector(to_unsigned(6,8) ,
57911	 => std_logic_vector(to_unsigned(10,8) ,
57912	 => std_logic_vector(to_unsigned(13,8) ,
57913	 => std_logic_vector(to_unsigned(17,8) ,
57914	 => std_logic_vector(to_unsigned(14,8) ,
57915	 => std_logic_vector(to_unsigned(12,8) ,
57916	 => std_logic_vector(to_unsigned(24,8) ,
57917	 => std_logic_vector(to_unsigned(20,8) ,
57918	 => std_logic_vector(to_unsigned(5,8) ,
57919	 => std_logic_vector(to_unsigned(8,8) ,
57920	 => std_logic_vector(to_unsigned(17,8) ,
57921	 => std_logic_vector(to_unsigned(85,8) ,
57922	 => std_logic_vector(to_unsigned(81,8) ,
57923	 => std_logic_vector(to_unsigned(80,8) ,
57924	 => std_logic_vector(to_unsigned(80,8) ,
57925	 => std_logic_vector(to_unsigned(47,8) ,
57926	 => std_logic_vector(to_unsigned(29,8) ,
57927	 => std_logic_vector(to_unsigned(27,8) ,
57928	 => std_logic_vector(to_unsigned(70,8) ,
57929	 => std_logic_vector(to_unsigned(114,8) ,
57930	 => std_logic_vector(to_unsigned(53,8) ,
57931	 => std_logic_vector(to_unsigned(69,8) ,
57932	 => std_logic_vector(to_unsigned(119,8) ,
57933	 => std_logic_vector(to_unsigned(85,8) ,
57934	 => std_logic_vector(to_unsigned(87,8) ,
57935	 => std_logic_vector(to_unsigned(81,8) ,
57936	 => std_logic_vector(to_unsigned(105,8) ,
57937	 => std_logic_vector(to_unsigned(93,8) ,
57938	 => std_logic_vector(to_unsigned(66,8) ,
57939	 => std_logic_vector(to_unsigned(49,8) ,
57940	 => std_logic_vector(to_unsigned(56,8) ,
57941	 => std_logic_vector(to_unsigned(50,8) ,
57942	 => std_logic_vector(to_unsigned(35,8) ,
57943	 => std_logic_vector(to_unsigned(34,8) ,
57944	 => std_logic_vector(to_unsigned(65,8) ,
57945	 => std_logic_vector(to_unsigned(92,8) ,
57946	 => std_logic_vector(to_unsigned(73,8) ,
57947	 => std_logic_vector(to_unsigned(82,8) ,
57948	 => std_logic_vector(to_unsigned(72,8) ,
57949	 => std_logic_vector(to_unsigned(57,8) ,
57950	 => std_logic_vector(to_unsigned(65,8) ,
57951	 => std_logic_vector(to_unsigned(79,8) ,
57952	 => std_logic_vector(to_unsigned(67,8) ,
57953	 => std_logic_vector(to_unsigned(69,8) ,
57954	 => std_logic_vector(to_unsigned(32,8) ,
57955	 => std_logic_vector(to_unsigned(22,8) ,
57956	 => std_logic_vector(to_unsigned(45,8) ,
57957	 => std_logic_vector(to_unsigned(58,8) ,
57958	 => std_logic_vector(to_unsigned(63,8) ,
57959	 => std_logic_vector(to_unsigned(67,8) ,
57960	 => std_logic_vector(to_unsigned(53,8) ,
57961	 => std_logic_vector(to_unsigned(30,8) ,
57962	 => std_logic_vector(to_unsigned(22,8) ,
57963	 => std_logic_vector(to_unsigned(31,8) ,
57964	 => std_logic_vector(to_unsigned(41,8) ,
57965	 => std_logic_vector(to_unsigned(29,8) ,
57966	 => std_logic_vector(to_unsigned(20,8) ,
57967	 => std_logic_vector(to_unsigned(37,8) ,
57968	 => std_logic_vector(to_unsigned(61,8) ,
57969	 => std_logic_vector(to_unsigned(49,8) ,
57970	 => std_logic_vector(to_unsigned(51,8) ,
57971	 => std_logic_vector(to_unsigned(60,8) ,
57972	 => std_logic_vector(to_unsigned(70,8) ,
57973	 => std_logic_vector(to_unsigned(64,8) ,
57974	 => std_logic_vector(to_unsigned(44,8) ,
57975	 => std_logic_vector(to_unsigned(58,8) ,
57976	 => std_logic_vector(to_unsigned(62,8) ,
57977	 => std_logic_vector(to_unsigned(48,8) ,
57978	 => std_logic_vector(to_unsigned(41,8) ,
57979	 => std_logic_vector(to_unsigned(41,8) ,
57980	 => std_logic_vector(to_unsigned(49,8) ,
57981	 => std_logic_vector(to_unsigned(63,8) ,
57982	 => std_logic_vector(to_unsigned(37,8) ,
57983	 => std_logic_vector(to_unsigned(63,8) ,
57984	 => std_logic_vector(to_unsigned(96,8) ,
57985	 => std_logic_vector(to_unsigned(96,8) ,
57986	 => std_logic_vector(to_unsigned(97,8) ,
57987	 => std_logic_vector(to_unsigned(76,8) ,
57988	 => std_logic_vector(to_unsigned(99,8) ,
57989	 => std_logic_vector(to_unsigned(100,8) ,
57990	 => std_logic_vector(to_unsigned(81,8) ,
57991	 => std_logic_vector(to_unsigned(108,8) ,
57992	 => std_logic_vector(to_unsigned(101,8) ,
57993	 => std_logic_vector(to_unsigned(103,8) ,
57994	 => std_logic_vector(to_unsigned(130,8) ,
57995	 => std_logic_vector(to_unsigned(149,8) ,
57996	 => std_logic_vector(to_unsigned(133,8) ,
57997	 => std_logic_vector(to_unsigned(134,8) ,
57998	 => std_logic_vector(to_unsigned(131,8) ,
57999	 => std_logic_vector(to_unsigned(115,8) ,
58000	 => std_logic_vector(to_unsigned(115,8) ,
58001	 => std_logic_vector(to_unsigned(130,8) ,
58002	 => std_logic_vector(to_unsigned(119,8) ,
58003	 => std_logic_vector(to_unsigned(109,8) ,
58004	 => std_logic_vector(to_unsigned(109,8) ,
58005	 => std_logic_vector(to_unsigned(103,8) ,
58006	 => std_logic_vector(to_unsigned(67,8) ,
58007	 => std_logic_vector(to_unsigned(40,8) ,
58008	 => std_logic_vector(to_unsigned(41,8) ,
58009	 => std_logic_vector(to_unsigned(37,8) ,
58010	 => std_logic_vector(to_unsigned(34,8) ,
58011	 => std_logic_vector(to_unsigned(32,8) ,
58012	 => std_logic_vector(to_unsigned(43,8) ,
58013	 => std_logic_vector(to_unsigned(47,8) ,
58014	 => std_logic_vector(to_unsigned(52,8) ,
58015	 => std_logic_vector(to_unsigned(71,8) ,
58016	 => std_logic_vector(to_unsigned(67,8) ,
58017	 => std_logic_vector(to_unsigned(47,8) ,
58018	 => std_logic_vector(to_unsigned(43,8) ,
58019	 => std_logic_vector(to_unsigned(48,8) ,
58020	 => std_logic_vector(to_unsigned(43,8) ,
58021	 => std_logic_vector(to_unsigned(41,8) ,
58022	 => std_logic_vector(to_unsigned(41,8) ,
58023	 => std_logic_vector(to_unsigned(44,8) ,
58024	 => std_logic_vector(to_unsigned(48,8) ,
58025	 => std_logic_vector(to_unsigned(41,8) ,
58026	 => std_logic_vector(to_unsigned(33,8) ,
58027	 => std_logic_vector(to_unsigned(32,8) ,
58028	 => std_logic_vector(to_unsigned(31,8) ,
58029	 => std_logic_vector(to_unsigned(77,8) ,
58030	 => std_logic_vector(to_unsigned(116,8) ,
58031	 => std_logic_vector(to_unsigned(63,8) ,
58032	 => std_logic_vector(to_unsigned(76,8) ,
58033	 => std_logic_vector(to_unsigned(78,8) ,
58034	 => std_logic_vector(to_unsigned(54,8) ,
58035	 => std_logic_vector(to_unsigned(54,8) ,
58036	 => std_logic_vector(to_unsigned(65,8) ,
58037	 => std_logic_vector(to_unsigned(51,8) ,
58038	 => std_logic_vector(to_unsigned(58,8) ,
58039	 => std_logic_vector(to_unsigned(32,8) ,
58040	 => std_logic_vector(to_unsigned(19,8) ,
58041	 => std_logic_vector(to_unsigned(32,8) ,
58042	 => std_logic_vector(to_unsigned(29,8) ,
58043	 => std_logic_vector(to_unsigned(34,8) ,
58044	 => std_logic_vector(to_unsigned(43,8) ,
58045	 => std_logic_vector(to_unsigned(35,8) ,
58046	 => std_logic_vector(to_unsigned(25,8) ,
58047	 => std_logic_vector(to_unsigned(41,8) ,
58048	 => std_logic_vector(to_unsigned(57,8) ,
58049	 => std_logic_vector(to_unsigned(65,8) ,
58050	 => std_logic_vector(to_unsigned(59,8) ,
58051	 => std_logic_vector(to_unsigned(46,8) ,
58052	 => std_logic_vector(to_unsigned(42,8) ,
58053	 => std_logic_vector(to_unsigned(48,8) ,
58054	 => std_logic_vector(to_unsigned(46,8) ,
58055	 => std_logic_vector(to_unsigned(59,8) ,
58056	 => std_logic_vector(to_unsigned(63,8) ,
58057	 => std_logic_vector(to_unsigned(19,8) ,
58058	 => std_logic_vector(to_unsigned(8,8) ,
58059	 => std_logic_vector(to_unsigned(14,8) ,
58060	 => std_logic_vector(to_unsigned(16,8) ,
58061	 => std_logic_vector(to_unsigned(9,8) ,
58062	 => std_logic_vector(to_unsigned(11,8) ,
58063	 => std_logic_vector(to_unsigned(14,8) ,
58064	 => std_logic_vector(to_unsigned(12,8) ,
58065	 => std_logic_vector(to_unsigned(24,8) ,
58066	 => std_logic_vector(to_unsigned(63,8) ,
58067	 => std_logic_vector(to_unsigned(22,8) ,
58068	 => std_logic_vector(to_unsigned(6,8) ,
58069	 => std_logic_vector(to_unsigned(47,8) ,
58070	 => std_logic_vector(to_unsigned(81,8) ,
58071	 => std_logic_vector(to_unsigned(36,8) ,
58072	 => std_logic_vector(to_unsigned(40,8) ,
58073	 => std_logic_vector(to_unsigned(82,8) ,
58074	 => std_logic_vector(to_unsigned(107,8) ,
58075	 => std_logic_vector(to_unsigned(79,8) ,
58076	 => std_logic_vector(to_unsigned(63,8) ,
58077	 => std_logic_vector(to_unsigned(60,8) ,
58078	 => std_logic_vector(to_unsigned(42,8) ,
58079	 => std_logic_vector(to_unsigned(34,8) ,
58080	 => std_logic_vector(to_unsigned(66,8) ,
58081	 => std_logic_vector(to_unsigned(138,8) ,
58082	 => std_logic_vector(to_unsigned(103,8) ,
58083	 => std_logic_vector(to_unsigned(87,8) ,
58084	 => std_logic_vector(to_unsigned(147,8) ,
58085	 => std_logic_vector(to_unsigned(131,8) ,
58086	 => std_logic_vector(to_unsigned(90,8) ,
58087	 => std_logic_vector(to_unsigned(23,8) ,
58088	 => std_logic_vector(to_unsigned(6,8) ,
58089	 => std_logic_vector(to_unsigned(6,8) ,
58090	 => std_logic_vector(to_unsigned(3,8) ,
58091	 => std_logic_vector(to_unsigned(5,8) ,
58092	 => std_logic_vector(to_unsigned(5,8) ,
58093	 => std_logic_vector(to_unsigned(8,8) ,
58094	 => std_logic_vector(to_unsigned(5,8) ,
58095	 => std_logic_vector(to_unsigned(6,8) ,
58096	 => std_logic_vector(to_unsigned(7,8) ,
58097	 => std_logic_vector(to_unsigned(10,8) ,
58098	 => std_logic_vector(to_unsigned(13,8) ,
58099	 => std_logic_vector(to_unsigned(17,8) ,
58100	 => std_logic_vector(to_unsigned(17,8) ,
58101	 => std_logic_vector(to_unsigned(17,8) ,
58102	 => std_logic_vector(to_unsigned(25,8) ,
58103	 => std_logic_vector(to_unsigned(35,8) ,
58104	 => std_logic_vector(to_unsigned(48,8) ,
58105	 => std_logic_vector(to_unsigned(47,8) ,
58106	 => std_logic_vector(to_unsigned(58,8) ,
58107	 => std_logic_vector(to_unsigned(74,8) ,
58108	 => std_logic_vector(to_unsigned(37,8) ,
58109	 => std_logic_vector(to_unsigned(14,8) ,
58110	 => std_logic_vector(to_unsigned(13,8) ,
58111	 => std_logic_vector(to_unsigned(29,8) ,
58112	 => std_logic_vector(to_unsigned(24,8) ,
58113	 => std_logic_vector(to_unsigned(25,8) ,
58114	 => std_logic_vector(to_unsigned(41,8) ,
58115	 => std_logic_vector(to_unsigned(30,8) ,
58116	 => std_logic_vector(to_unsigned(18,8) ,
58117	 => std_logic_vector(to_unsigned(22,8) ,
58118	 => std_logic_vector(to_unsigned(28,8) ,
58119	 => std_logic_vector(to_unsigned(27,8) ,
58120	 => std_logic_vector(to_unsigned(23,8) ,
58121	 => std_logic_vector(to_unsigned(40,8) ,
58122	 => std_logic_vector(to_unsigned(54,8) ,
58123	 => std_logic_vector(to_unsigned(37,8) ,
58124	 => std_logic_vector(to_unsigned(25,8) ,
58125	 => std_logic_vector(to_unsigned(35,8) ,
58126	 => std_logic_vector(to_unsigned(15,8) ,
58127	 => std_logic_vector(to_unsigned(18,8) ,
58128	 => std_logic_vector(to_unsigned(28,8) ,
58129	 => std_logic_vector(to_unsigned(27,8) ,
58130	 => std_logic_vector(to_unsigned(24,8) ,
58131	 => std_logic_vector(to_unsigned(20,8) ,
58132	 => std_logic_vector(to_unsigned(27,8) ,
58133	 => std_logic_vector(to_unsigned(23,8) ,
58134	 => std_logic_vector(to_unsigned(6,8) ,
58135	 => std_logic_vector(to_unsigned(13,8) ,
58136	 => std_logic_vector(to_unsigned(17,8) ,
58137	 => std_logic_vector(to_unsigned(10,8) ,
58138	 => std_logic_vector(to_unsigned(10,8) ,
58139	 => std_logic_vector(to_unsigned(6,8) ,
58140	 => std_logic_vector(to_unsigned(5,8) ,
58141	 => std_logic_vector(to_unsigned(6,8) ,
58142	 => std_logic_vector(to_unsigned(6,8) ,
58143	 => std_logic_vector(to_unsigned(29,8) ,
58144	 => std_logic_vector(to_unsigned(41,8) ,
58145	 => std_logic_vector(to_unsigned(27,8) ,
58146	 => std_logic_vector(to_unsigned(19,8) ,
58147	 => std_logic_vector(to_unsigned(12,8) ,
58148	 => std_logic_vector(to_unsigned(15,8) ,
58149	 => std_logic_vector(to_unsigned(16,8) ,
58150	 => std_logic_vector(to_unsigned(14,8) ,
58151	 => std_logic_vector(to_unsigned(16,8) ,
58152	 => std_logic_vector(to_unsigned(15,8) ,
58153	 => std_logic_vector(to_unsigned(16,8) ,
58154	 => std_logic_vector(to_unsigned(23,8) ,
58155	 => std_logic_vector(to_unsigned(24,8) ,
58156	 => std_logic_vector(to_unsigned(16,8) ,
58157	 => std_logic_vector(to_unsigned(21,8) ,
58158	 => std_logic_vector(to_unsigned(32,8) ,
58159	 => std_logic_vector(to_unsigned(46,8) ,
58160	 => std_logic_vector(to_unsigned(88,8) ,
58161	 => std_logic_vector(to_unsigned(69,8) ,
58162	 => std_logic_vector(to_unsigned(27,8) ,
58163	 => std_logic_vector(to_unsigned(38,8) ,
58164	 => std_logic_vector(to_unsigned(46,8) ,
58165	 => std_logic_vector(to_unsigned(47,8) ,
58166	 => std_logic_vector(to_unsigned(34,8) ,
58167	 => std_logic_vector(to_unsigned(13,8) ,
58168	 => std_logic_vector(to_unsigned(15,8) ,
58169	 => std_logic_vector(to_unsigned(10,8) ,
58170	 => std_logic_vector(to_unsigned(10,8) ,
58171	 => std_logic_vector(to_unsigned(8,8) ,
58172	 => std_logic_vector(to_unsigned(5,8) ,
58173	 => std_logic_vector(to_unsigned(6,8) ,
58174	 => std_logic_vector(to_unsigned(7,8) ,
58175	 => std_logic_vector(to_unsigned(8,8) ,
58176	 => std_logic_vector(to_unsigned(6,8) ,
58177	 => std_logic_vector(to_unsigned(7,8) ,
58178	 => std_logic_vector(to_unsigned(11,8) ,
58179	 => std_logic_vector(to_unsigned(10,8) ,
58180	 => std_logic_vector(to_unsigned(12,8) ,
58181	 => std_logic_vector(to_unsigned(10,8) ,
58182	 => std_logic_vector(to_unsigned(6,8) ,
58183	 => std_logic_vector(to_unsigned(1,8) ,
58184	 => std_logic_vector(to_unsigned(0,8) ,
58185	 => std_logic_vector(to_unsigned(8,8) ,
58186	 => std_logic_vector(to_unsigned(20,8) ,
58187	 => std_logic_vector(to_unsigned(16,8) ,
58188	 => std_logic_vector(to_unsigned(35,8) ,
58189	 => std_logic_vector(to_unsigned(32,8) ,
58190	 => std_logic_vector(to_unsigned(43,8) ,
58191	 => std_logic_vector(to_unsigned(30,8) ,
58192	 => std_logic_vector(to_unsigned(41,8) ,
58193	 => std_logic_vector(to_unsigned(23,8) ,
58194	 => std_logic_vector(to_unsigned(12,8) ,
58195	 => std_logic_vector(to_unsigned(7,8) ,
58196	 => std_logic_vector(to_unsigned(10,8) ,
58197	 => std_logic_vector(to_unsigned(8,8) ,
58198	 => std_logic_vector(to_unsigned(7,8) ,
58199	 => std_logic_vector(to_unsigned(12,8) ,
58200	 => std_logic_vector(to_unsigned(9,8) ,
58201	 => std_logic_vector(to_unsigned(7,8) ,
58202	 => std_logic_vector(to_unsigned(6,8) ,
58203	 => std_logic_vector(to_unsigned(1,8) ,
58204	 => std_logic_vector(to_unsigned(0,8) ,
58205	 => std_logic_vector(to_unsigned(1,8) ,
58206	 => std_logic_vector(to_unsigned(1,8) ,
58207	 => std_logic_vector(to_unsigned(6,8) ,
58208	 => std_logic_vector(to_unsigned(3,8) ,
58209	 => std_logic_vector(to_unsigned(0,8) ,
58210	 => std_logic_vector(to_unsigned(0,8) ,
58211	 => std_logic_vector(to_unsigned(1,8) ,
58212	 => std_logic_vector(to_unsigned(1,8) ,
58213	 => std_logic_vector(to_unsigned(2,8) ,
58214	 => std_logic_vector(to_unsigned(15,8) ,
58215	 => std_logic_vector(to_unsigned(18,8) ,
58216	 => std_logic_vector(to_unsigned(7,8) ,
58217	 => std_logic_vector(to_unsigned(7,8) ,
58218	 => std_logic_vector(to_unsigned(13,8) ,
58219	 => std_logic_vector(to_unsigned(19,8) ,
58220	 => std_logic_vector(to_unsigned(12,8) ,
58221	 => std_logic_vector(to_unsigned(11,8) ,
58222	 => std_logic_vector(to_unsigned(22,8) ,
58223	 => std_logic_vector(to_unsigned(22,8) ,
58224	 => std_logic_vector(to_unsigned(25,8) ,
58225	 => std_logic_vector(to_unsigned(49,8) ,
58226	 => std_logic_vector(to_unsigned(13,8) ,
58227	 => std_logic_vector(to_unsigned(7,8) ,
58228	 => std_logic_vector(to_unsigned(13,8) ,
58229	 => std_logic_vector(to_unsigned(13,8) ,
58230	 => std_logic_vector(to_unsigned(6,8) ,
58231	 => std_logic_vector(to_unsigned(8,8) ,
58232	 => std_logic_vector(to_unsigned(19,8) ,
58233	 => std_logic_vector(to_unsigned(30,8) ,
58234	 => std_logic_vector(to_unsigned(15,8) ,
58235	 => std_logic_vector(to_unsigned(6,8) ,
58236	 => std_logic_vector(to_unsigned(15,8) ,
58237	 => std_logic_vector(to_unsigned(18,8) ,
58238	 => std_logic_vector(to_unsigned(6,8) ,
58239	 => std_logic_vector(to_unsigned(12,8) ,
58240	 => std_logic_vector(to_unsigned(18,8) ,
58241	 => std_logic_vector(to_unsigned(97,8) ,
58242	 => std_logic_vector(to_unsigned(93,8) ,
58243	 => std_logic_vector(to_unsigned(70,8) ,
58244	 => std_logic_vector(to_unsigned(79,8) ,
58245	 => std_logic_vector(to_unsigned(49,8) ,
58246	 => std_logic_vector(to_unsigned(29,8) ,
58247	 => std_logic_vector(to_unsigned(32,8) ,
58248	 => std_logic_vector(to_unsigned(58,8) ,
58249	 => std_logic_vector(to_unsigned(52,8) ,
58250	 => std_logic_vector(to_unsigned(50,8) ,
58251	 => std_logic_vector(to_unsigned(76,8) ,
58252	 => std_logic_vector(to_unsigned(77,8) ,
58253	 => std_logic_vector(to_unsigned(67,8) ,
58254	 => std_logic_vector(to_unsigned(93,8) ,
58255	 => std_logic_vector(to_unsigned(69,8) ,
58256	 => std_logic_vector(to_unsigned(48,8) ,
58257	 => std_logic_vector(to_unsigned(85,8) ,
58258	 => std_logic_vector(to_unsigned(57,8) ,
58259	 => std_logic_vector(to_unsigned(41,8) ,
58260	 => std_logic_vector(to_unsigned(62,8) ,
58261	 => std_logic_vector(to_unsigned(60,8) ,
58262	 => std_logic_vector(to_unsigned(36,8) ,
58263	 => std_logic_vector(to_unsigned(32,8) ,
58264	 => std_logic_vector(to_unsigned(64,8) ,
58265	 => std_logic_vector(to_unsigned(95,8) ,
58266	 => std_logic_vector(to_unsigned(69,8) ,
58267	 => std_logic_vector(to_unsigned(76,8) ,
58268	 => std_logic_vector(to_unsigned(61,8) ,
58269	 => std_logic_vector(to_unsigned(52,8) ,
58270	 => std_logic_vector(to_unsigned(52,8) ,
58271	 => std_logic_vector(to_unsigned(44,8) ,
58272	 => std_logic_vector(to_unsigned(47,8) ,
58273	 => std_logic_vector(to_unsigned(53,8) ,
58274	 => std_logic_vector(to_unsigned(53,8) ,
58275	 => std_logic_vector(to_unsigned(39,8) ,
58276	 => std_logic_vector(to_unsigned(37,8) ,
58277	 => std_logic_vector(to_unsigned(51,8) ,
58278	 => std_logic_vector(to_unsigned(57,8) ,
58279	 => std_logic_vector(to_unsigned(61,8) ,
58280	 => std_logic_vector(to_unsigned(45,8) ,
58281	 => std_logic_vector(to_unsigned(26,8) ,
58282	 => std_logic_vector(to_unsigned(24,8) ,
58283	 => std_logic_vector(to_unsigned(33,8) ,
58284	 => std_logic_vector(to_unsigned(40,8) ,
58285	 => std_logic_vector(to_unsigned(32,8) ,
58286	 => std_logic_vector(to_unsigned(27,8) ,
58287	 => std_logic_vector(to_unsigned(51,8) ,
58288	 => std_logic_vector(to_unsigned(70,8) ,
58289	 => std_logic_vector(to_unsigned(50,8) ,
58290	 => std_logic_vector(to_unsigned(47,8) ,
58291	 => std_logic_vector(to_unsigned(57,8) ,
58292	 => std_logic_vector(to_unsigned(67,8) ,
58293	 => std_logic_vector(to_unsigned(62,8) ,
58294	 => std_logic_vector(to_unsigned(55,8) ,
58295	 => std_logic_vector(to_unsigned(56,8) ,
58296	 => std_logic_vector(to_unsigned(45,8) ,
58297	 => std_logic_vector(to_unsigned(48,8) ,
58298	 => std_logic_vector(to_unsigned(57,8) ,
58299	 => std_logic_vector(to_unsigned(49,8) ,
58300	 => std_logic_vector(to_unsigned(48,8) ,
58301	 => std_logic_vector(to_unsigned(68,8) ,
58302	 => std_logic_vector(to_unsigned(49,8) ,
58303	 => std_logic_vector(to_unsigned(69,8) ,
58304	 => std_logic_vector(to_unsigned(99,8) ,
58305	 => std_logic_vector(to_unsigned(95,8) ,
58306	 => std_logic_vector(to_unsigned(90,8) ,
58307	 => std_logic_vector(to_unsigned(77,8) ,
58308	 => std_logic_vector(to_unsigned(90,8) ,
58309	 => std_logic_vector(to_unsigned(91,8) ,
58310	 => std_logic_vector(to_unsigned(78,8) ,
58311	 => std_logic_vector(to_unsigned(109,8) ,
58312	 => std_logic_vector(to_unsigned(119,8) ,
58313	 => std_logic_vector(to_unsigned(121,8) ,
58314	 => std_logic_vector(to_unsigned(139,8) ,
58315	 => std_logic_vector(to_unsigned(147,8) ,
58316	 => std_logic_vector(to_unsigned(136,8) ,
58317	 => std_logic_vector(to_unsigned(131,8) ,
58318	 => std_logic_vector(to_unsigned(122,8) ,
58319	 => std_logic_vector(to_unsigned(118,8) ,
58320	 => std_logic_vector(to_unsigned(131,8) ,
58321	 => std_logic_vector(to_unsigned(127,8) ,
58322	 => std_logic_vector(to_unsigned(107,8) ,
58323	 => std_logic_vector(to_unsigned(114,8) ,
58324	 => std_logic_vector(to_unsigned(109,8) ,
58325	 => std_logic_vector(to_unsigned(121,8) ,
58326	 => std_logic_vector(to_unsigned(79,8) ,
58327	 => std_logic_vector(to_unsigned(34,8) ,
58328	 => std_logic_vector(to_unsigned(37,8) ,
58329	 => std_logic_vector(to_unsigned(39,8) ,
58330	 => std_logic_vector(to_unsigned(41,8) ,
58331	 => std_logic_vector(to_unsigned(44,8) ,
58332	 => std_logic_vector(to_unsigned(45,8) ,
58333	 => std_logic_vector(to_unsigned(42,8) ,
58334	 => std_logic_vector(to_unsigned(43,8) ,
58335	 => std_logic_vector(to_unsigned(51,8) ,
58336	 => std_logic_vector(to_unsigned(53,8) ,
58337	 => std_logic_vector(to_unsigned(59,8) ,
58338	 => std_logic_vector(to_unsigned(70,8) ,
58339	 => std_logic_vector(to_unsigned(55,8) ,
58340	 => std_logic_vector(to_unsigned(47,8) ,
58341	 => std_logic_vector(to_unsigned(44,8) ,
58342	 => std_logic_vector(to_unsigned(44,8) ,
58343	 => std_logic_vector(to_unsigned(48,8) ,
58344	 => std_logic_vector(to_unsigned(50,8) ,
58345	 => std_logic_vector(to_unsigned(45,8) ,
58346	 => std_logic_vector(to_unsigned(41,8) ,
58347	 => std_logic_vector(to_unsigned(32,8) ,
58348	 => std_logic_vector(to_unsigned(45,8) ,
58349	 => std_logic_vector(to_unsigned(86,8) ,
58350	 => std_logic_vector(to_unsigned(85,8) ,
58351	 => std_logic_vector(to_unsigned(65,8) ,
58352	 => std_logic_vector(to_unsigned(73,8) ,
58353	 => std_logic_vector(to_unsigned(71,8) ,
58354	 => std_logic_vector(to_unsigned(51,8) ,
58355	 => std_logic_vector(to_unsigned(48,8) ,
58356	 => std_logic_vector(to_unsigned(65,8) ,
58357	 => std_logic_vector(to_unsigned(51,8) ,
58358	 => std_logic_vector(to_unsigned(44,8) ,
58359	 => std_logic_vector(to_unsigned(31,8) ,
58360	 => std_logic_vector(to_unsigned(47,8) ,
58361	 => std_logic_vector(to_unsigned(71,8) ,
58362	 => std_logic_vector(to_unsigned(66,8) ,
58363	 => std_logic_vector(to_unsigned(54,8) ,
58364	 => std_logic_vector(to_unsigned(50,8) ,
58365	 => std_logic_vector(to_unsigned(30,8) ,
58366	 => std_logic_vector(to_unsigned(21,8) ,
58367	 => std_logic_vector(to_unsigned(22,8) ,
58368	 => std_logic_vector(to_unsigned(19,8) ,
58369	 => std_logic_vector(to_unsigned(34,8) ,
58370	 => std_logic_vector(to_unsigned(74,8) ,
58371	 => std_logic_vector(to_unsigned(47,8) ,
58372	 => std_logic_vector(to_unsigned(47,8) ,
58373	 => std_logic_vector(to_unsigned(33,8) ,
58374	 => std_logic_vector(to_unsigned(33,8) ,
58375	 => std_logic_vector(to_unsigned(45,8) ,
58376	 => std_logic_vector(to_unsigned(21,8) ,
58377	 => std_logic_vector(to_unsigned(9,8) ,
58378	 => std_logic_vector(to_unsigned(12,8) ,
58379	 => std_logic_vector(to_unsigned(12,8) ,
58380	 => std_logic_vector(to_unsigned(10,8) ,
58381	 => std_logic_vector(to_unsigned(12,8) ,
58382	 => std_logic_vector(to_unsigned(14,8) ,
58383	 => std_logic_vector(to_unsigned(12,8) ,
58384	 => std_logic_vector(to_unsigned(14,8) ,
58385	 => std_logic_vector(to_unsigned(41,8) ,
58386	 => std_logic_vector(to_unsigned(64,8) ,
58387	 => std_logic_vector(to_unsigned(19,8) ,
58388	 => std_logic_vector(to_unsigned(3,8) ,
58389	 => std_logic_vector(to_unsigned(29,8) ,
58390	 => std_logic_vector(to_unsigned(88,8) ,
58391	 => std_logic_vector(to_unsigned(27,8) ,
58392	 => std_logic_vector(to_unsigned(32,8) ,
58393	 => std_logic_vector(to_unsigned(50,8) ,
58394	 => std_logic_vector(to_unsigned(44,8) ,
58395	 => std_logic_vector(to_unsigned(33,8) ,
58396	 => std_logic_vector(to_unsigned(29,8) ,
58397	 => std_logic_vector(to_unsigned(30,8) ,
58398	 => std_logic_vector(to_unsigned(35,8) ,
58399	 => std_logic_vector(to_unsigned(30,8) ,
58400	 => std_logic_vector(to_unsigned(59,8) ,
58401	 => std_logic_vector(to_unsigned(151,8) ,
58402	 => std_logic_vector(to_unsigned(74,8) ,
58403	 => std_logic_vector(to_unsigned(41,8) ,
58404	 => std_logic_vector(to_unsigned(134,8) ,
58405	 => std_logic_vector(to_unsigned(131,8) ,
58406	 => std_logic_vector(to_unsigned(103,8) ,
58407	 => std_logic_vector(to_unsigned(51,8) ,
58408	 => std_logic_vector(to_unsigned(21,8) ,
58409	 => std_logic_vector(to_unsigned(25,8) ,
58410	 => std_logic_vector(to_unsigned(18,8) ,
58411	 => std_logic_vector(to_unsigned(11,8) ,
58412	 => std_logic_vector(to_unsigned(8,8) ,
58413	 => std_logic_vector(to_unsigned(7,8) ,
58414	 => std_logic_vector(to_unsigned(5,8) ,
58415	 => std_logic_vector(to_unsigned(5,8) ,
58416	 => std_logic_vector(to_unsigned(6,8) ,
58417	 => std_logic_vector(to_unsigned(6,8) ,
58418	 => std_logic_vector(to_unsigned(5,8) ,
58419	 => std_logic_vector(to_unsigned(8,8) ,
58420	 => std_logic_vector(to_unsigned(9,8) ,
58421	 => std_logic_vector(to_unsigned(11,8) ,
58422	 => std_logic_vector(to_unsigned(8,8) ,
58423	 => std_logic_vector(to_unsigned(10,8) ,
58424	 => std_logic_vector(to_unsigned(16,8) ,
58425	 => std_logic_vector(to_unsigned(16,8) ,
58426	 => std_logic_vector(to_unsigned(25,8) ,
58427	 => std_logic_vector(to_unsigned(30,8) ,
58428	 => std_logic_vector(to_unsigned(18,8) ,
58429	 => std_logic_vector(to_unsigned(22,8) ,
58430	 => std_logic_vector(to_unsigned(26,8) ,
58431	 => std_logic_vector(to_unsigned(30,8) ,
58432	 => std_logic_vector(to_unsigned(30,8) ,
58433	 => std_logic_vector(to_unsigned(53,8) ,
58434	 => std_logic_vector(to_unsigned(81,8) ,
58435	 => std_logic_vector(to_unsigned(74,8) ,
58436	 => std_logic_vector(to_unsigned(33,8) ,
58437	 => std_logic_vector(to_unsigned(26,8) ,
58438	 => std_logic_vector(to_unsigned(31,8) ,
58439	 => std_logic_vector(to_unsigned(28,8) ,
58440	 => std_logic_vector(to_unsigned(19,8) ,
58441	 => std_logic_vector(to_unsigned(45,8) ,
58442	 => std_logic_vector(to_unsigned(57,8) ,
58443	 => std_logic_vector(to_unsigned(36,8) ,
58444	 => std_logic_vector(to_unsigned(26,8) ,
58445	 => std_logic_vector(to_unsigned(27,8) ,
58446	 => std_logic_vector(to_unsigned(25,8) ,
58447	 => std_logic_vector(to_unsigned(11,8) ,
58448	 => std_logic_vector(to_unsigned(9,8) ,
58449	 => std_logic_vector(to_unsigned(25,8) ,
58450	 => std_logic_vector(to_unsigned(19,8) ,
58451	 => std_logic_vector(to_unsigned(11,8) ,
58452	 => std_logic_vector(to_unsigned(7,8) ,
58453	 => std_logic_vector(to_unsigned(12,8) ,
58454	 => std_logic_vector(to_unsigned(15,8) ,
58455	 => std_logic_vector(to_unsigned(22,8) ,
58456	 => std_logic_vector(to_unsigned(24,8) ,
58457	 => std_logic_vector(to_unsigned(20,8) ,
58458	 => std_logic_vector(to_unsigned(23,8) ,
58459	 => std_logic_vector(to_unsigned(12,8) ,
58460	 => std_logic_vector(to_unsigned(12,8) ,
58461	 => std_logic_vector(to_unsigned(13,8) ,
58462	 => std_logic_vector(to_unsigned(22,8) ,
58463	 => std_logic_vector(to_unsigned(41,8) ,
58464	 => std_logic_vector(to_unsigned(27,8) ,
58465	 => std_logic_vector(to_unsigned(24,8) ,
58466	 => std_logic_vector(to_unsigned(18,8) ,
58467	 => std_logic_vector(to_unsigned(7,8) ,
58468	 => std_logic_vector(to_unsigned(14,8) ,
58469	 => std_logic_vector(to_unsigned(16,8) ,
58470	 => std_logic_vector(to_unsigned(16,8) ,
58471	 => std_logic_vector(to_unsigned(18,8) ,
58472	 => std_logic_vector(to_unsigned(13,8) ,
58473	 => std_logic_vector(to_unsigned(17,8) ,
58474	 => std_logic_vector(to_unsigned(27,8) ,
58475	 => std_logic_vector(to_unsigned(27,8) ,
58476	 => std_logic_vector(to_unsigned(22,8) ,
58477	 => std_logic_vector(to_unsigned(37,8) ,
58478	 => std_logic_vector(to_unsigned(30,8) ,
58479	 => std_logic_vector(to_unsigned(38,8) ,
58480	 => std_logic_vector(to_unsigned(85,8) ,
58481	 => std_logic_vector(to_unsigned(87,8) ,
58482	 => std_logic_vector(to_unsigned(50,8) ,
58483	 => std_logic_vector(to_unsigned(35,8) ,
58484	 => std_logic_vector(to_unsigned(33,8) ,
58485	 => std_logic_vector(to_unsigned(44,8) ,
58486	 => std_logic_vector(to_unsigned(35,8) ,
58487	 => std_logic_vector(to_unsigned(20,8) ,
58488	 => std_logic_vector(to_unsigned(12,8) ,
58489	 => std_logic_vector(to_unsigned(11,8) ,
58490	 => std_logic_vector(to_unsigned(47,8) ,
58491	 => std_logic_vector(to_unsigned(58,8) ,
58492	 => std_logic_vector(to_unsigned(37,8) ,
58493	 => std_logic_vector(to_unsigned(14,8) ,
58494	 => std_logic_vector(to_unsigned(8,8) ,
58495	 => std_logic_vector(to_unsigned(7,8) ,
58496	 => std_logic_vector(to_unsigned(6,8) ,
58497	 => std_logic_vector(to_unsigned(6,8) ,
58498	 => std_logic_vector(to_unsigned(9,8) ,
58499	 => std_logic_vector(to_unsigned(7,8) ,
58500	 => std_logic_vector(to_unsigned(8,8) ,
58501	 => std_logic_vector(to_unsigned(6,8) ,
58502	 => std_logic_vector(to_unsigned(11,8) ,
58503	 => std_logic_vector(to_unsigned(3,8) ,
58504	 => std_logic_vector(to_unsigned(0,8) ,
58505	 => std_logic_vector(to_unsigned(3,8) ,
58506	 => std_logic_vector(to_unsigned(25,8) ,
58507	 => std_logic_vector(to_unsigned(25,8) ,
58508	 => std_logic_vector(to_unsigned(42,8) ,
58509	 => std_logic_vector(to_unsigned(44,8) ,
58510	 => std_logic_vector(to_unsigned(42,8) ,
58511	 => std_logic_vector(to_unsigned(25,8) ,
58512	 => std_logic_vector(to_unsigned(46,8) ,
58513	 => std_logic_vector(to_unsigned(33,8) ,
58514	 => std_logic_vector(to_unsigned(15,8) ,
58515	 => std_logic_vector(to_unsigned(14,8) ,
58516	 => std_logic_vector(to_unsigned(14,8) ,
58517	 => std_logic_vector(to_unsigned(9,8) ,
58518	 => std_logic_vector(to_unsigned(8,8) ,
58519	 => std_logic_vector(to_unsigned(9,8) ,
58520	 => std_logic_vector(to_unsigned(6,8) ,
58521	 => std_logic_vector(to_unsigned(8,8) ,
58522	 => std_logic_vector(to_unsigned(3,8) ,
58523	 => std_logic_vector(to_unsigned(0,8) ,
58524	 => std_logic_vector(to_unsigned(0,8) ,
58525	 => std_logic_vector(to_unsigned(0,8) ,
58526	 => std_logic_vector(to_unsigned(0,8) ,
58527	 => std_logic_vector(to_unsigned(2,8) ,
58528	 => std_logic_vector(to_unsigned(3,8) ,
58529	 => std_logic_vector(to_unsigned(3,8) ,
58530	 => std_logic_vector(to_unsigned(2,8) ,
58531	 => std_logic_vector(to_unsigned(6,8) ,
58532	 => std_logic_vector(to_unsigned(14,8) ,
58533	 => std_logic_vector(to_unsigned(9,8) ,
58534	 => std_logic_vector(to_unsigned(13,8) ,
58535	 => std_logic_vector(to_unsigned(17,8) ,
58536	 => std_logic_vector(to_unsigned(13,8) ,
58537	 => std_logic_vector(to_unsigned(7,8) ,
58538	 => std_logic_vector(to_unsigned(16,8) ,
58539	 => std_logic_vector(to_unsigned(26,8) ,
58540	 => std_logic_vector(to_unsigned(17,8) ,
58541	 => std_logic_vector(to_unsigned(14,8) ,
58542	 => std_logic_vector(to_unsigned(13,8) ,
58543	 => std_logic_vector(to_unsigned(12,8) ,
58544	 => std_logic_vector(to_unsigned(17,8) ,
58545	 => std_logic_vector(to_unsigned(27,8) ,
58546	 => std_logic_vector(to_unsigned(13,8) ,
58547	 => std_logic_vector(to_unsigned(9,8) ,
58548	 => std_logic_vector(to_unsigned(10,8) ,
58549	 => std_logic_vector(to_unsigned(9,8) ,
58550	 => std_logic_vector(to_unsigned(5,8) ,
58551	 => std_logic_vector(to_unsigned(7,8) ,
58552	 => std_logic_vector(to_unsigned(12,8) ,
58553	 => std_logic_vector(to_unsigned(11,8) ,
58554	 => std_logic_vector(to_unsigned(13,8) ,
58555	 => std_logic_vector(to_unsigned(9,8) ,
58556	 => std_logic_vector(to_unsigned(14,8) ,
58557	 => std_logic_vector(to_unsigned(11,8) ,
58558	 => std_logic_vector(to_unsigned(4,8) ,
58559	 => std_logic_vector(to_unsigned(10,8) ,
58560	 => std_logic_vector(to_unsigned(11,8) ,
58561	 => std_logic_vector(to_unsigned(96,8) ,
58562	 => std_logic_vector(to_unsigned(97,8) ,
58563	 => std_logic_vector(to_unsigned(66,8) ,
58564	 => std_logic_vector(to_unsigned(76,8) ,
58565	 => std_logic_vector(to_unsigned(63,8) ,
58566	 => std_logic_vector(to_unsigned(37,8) ,
58567	 => std_logic_vector(to_unsigned(25,8) ,
58568	 => std_logic_vector(to_unsigned(48,8) ,
58569	 => std_logic_vector(to_unsigned(48,8) ,
58570	 => std_logic_vector(to_unsigned(53,8) ,
58571	 => std_logic_vector(to_unsigned(62,8) ,
58572	 => std_logic_vector(to_unsigned(34,8) ,
58573	 => std_logic_vector(to_unsigned(49,8) ,
58574	 => std_logic_vector(to_unsigned(96,8) ,
58575	 => std_logic_vector(to_unsigned(77,8) ,
58576	 => std_logic_vector(to_unsigned(45,8) ,
58577	 => std_logic_vector(to_unsigned(77,8) ,
58578	 => std_logic_vector(to_unsigned(64,8) ,
58579	 => std_logic_vector(to_unsigned(53,8) ,
58580	 => std_logic_vector(to_unsigned(68,8) ,
58581	 => std_logic_vector(to_unsigned(53,8) ,
58582	 => std_logic_vector(to_unsigned(32,8) ,
58583	 => std_logic_vector(to_unsigned(33,8) ,
58584	 => std_logic_vector(to_unsigned(61,8) ,
58585	 => std_logic_vector(to_unsigned(87,8) ,
58586	 => std_logic_vector(to_unsigned(56,8) ,
58587	 => std_logic_vector(to_unsigned(64,8) ,
58588	 => std_logic_vector(to_unsigned(60,8) ,
58589	 => std_logic_vector(to_unsigned(62,8) ,
58590	 => std_logic_vector(to_unsigned(27,8) ,
58591	 => std_logic_vector(to_unsigned(18,8) ,
58592	 => std_logic_vector(to_unsigned(51,8) ,
58593	 => std_logic_vector(to_unsigned(59,8) ,
58594	 => std_logic_vector(to_unsigned(57,8) ,
58595	 => std_logic_vector(to_unsigned(51,8) ,
58596	 => std_logic_vector(to_unsigned(32,8) ,
58597	 => std_logic_vector(to_unsigned(39,8) ,
58598	 => std_logic_vector(to_unsigned(52,8) ,
58599	 => std_logic_vector(to_unsigned(60,8) ,
58600	 => std_logic_vector(to_unsigned(51,8) ,
58601	 => std_logic_vector(to_unsigned(38,8) ,
58602	 => std_logic_vector(to_unsigned(41,8) ,
58603	 => std_logic_vector(to_unsigned(51,8) ,
58604	 => std_logic_vector(to_unsigned(45,8) ,
58605	 => std_logic_vector(to_unsigned(41,8) ,
58606	 => std_logic_vector(to_unsigned(51,8) ,
58607	 => std_logic_vector(to_unsigned(63,8) ,
58608	 => std_logic_vector(to_unsigned(68,8) ,
58609	 => std_logic_vector(to_unsigned(74,8) ,
58610	 => std_logic_vector(to_unsigned(80,8) ,
58611	 => std_logic_vector(to_unsigned(85,8) ,
58612	 => std_logic_vector(to_unsigned(79,8) ,
58613	 => std_logic_vector(to_unsigned(72,8) ,
58614	 => std_logic_vector(to_unsigned(86,8) ,
58615	 => std_logic_vector(to_unsigned(91,8) ,
58616	 => std_logic_vector(to_unsigned(82,8) ,
58617	 => std_logic_vector(to_unsigned(78,8) ,
58618	 => std_logic_vector(to_unsigned(56,8) ,
58619	 => std_logic_vector(to_unsigned(51,8) ,
58620	 => std_logic_vector(to_unsigned(51,8) ,
58621	 => std_logic_vector(to_unsigned(46,8) ,
58622	 => std_logic_vector(to_unsigned(37,8) ,
58623	 => std_logic_vector(to_unsigned(76,8) ,
58624	 => std_logic_vector(to_unsigned(69,8) ,
58625	 => std_logic_vector(to_unsigned(64,8) ,
58626	 => std_logic_vector(to_unsigned(96,8) ,
58627	 => std_logic_vector(to_unsigned(73,8) ,
58628	 => std_logic_vector(to_unsigned(92,8) ,
58629	 => std_logic_vector(to_unsigned(86,8) ,
58630	 => std_logic_vector(to_unsigned(86,8) ,
58631	 => std_logic_vector(to_unsigned(111,8) ,
58632	 => std_logic_vector(to_unsigned(111,8) ,
58633	 => std_logic_vector(to_unsigned(105,8) ,
58634	 => std_logic_vector(to_unsigned(136,8) ,
58635	 => std_logic_vector(to_unsigned(154,8) ,
58636	 => std_logic_vector(to_unsigned(125,8) ,
58637	 => std_logic_vector(to_unsigned(118,8) ,
58638	 => std_logic_vector(to_unsigned(127,8) ,
58639	 => std_logic_vector(to_unsigned(124,8) ,
58640	 => std_logic_vector(to_unsigned(119,8) ,
58641	 => std_logic_vector(to_unsigned(122,8) ,
58642	 => std_logic_vector(to_unsigned(116,8) ,
58643	 => std_logic_vector(to_unsigned(116,8) ,
58644	 => std_logic_vector(to_unsigned(111,8) ,
58645	 => std_logic_vector(to_unsigned(133,8) ,
58646	 => std_logic_vector(to_unsigned(86,8) ,
58647	 => std_logic_vector(to_unsigned(31,8) ,
58648	 => std_logic_vector(to_unsigned(35,8) ,
58649	 => std_logic_vector(to_unsigned(43,8) ,
58650	 => std_logic_vector(to_unsigned(42,8) ,
58651	 => std_logic_vector(to_unsigned(54,8) ,
58652	 => std_logic_vector(to_unsigned(52,8) ,
58653	 => std_logic_vector(to_unsigned(47,8) ,
58654	 => std_logic_vector(to_unsigned(48,8) ,
58655	 => std_logic_vector(to_unsigned(51,8) ,
58656	 => std_logic_vector(to_unsigned(57,8) ,
58657	 => std_logic_vector(to_unsigned(64,8) ,
58658	 => std_logic_vector(to_unsigned(68,8) ,
58659	 => std_logic_vector(to_unsigned(67,8) ,
58660	 => std_logic_vector(to_unsigned(69,8) ,
58661	 => std_logic_vector(to_unsigned(51,8) ,
58662	 => std_logic_vector(to_unsigned(47,8) ,
58663	 => std_logic_vector(to_unsigned(63,8) ,
58664	 => std_logic_vector(to_unsigned(62,8) ,
58665	 => std_logic_vector(to_unsigned(56,8) ,
58666	 => std_logic_vector(to_unsigned(51,8) ,
58667	 => std_logic_vector(to_unsigned(68,8) ,
58668	 => std_logic_vector(to_unsigned(107,8) ,
58669	 => std_logic_vector(to_unsigned(76,8) ,
58670	 => std_logic_vector(to_unsigned(61,8) ,
58671	 => std_logic_vector(to_unsigned(60,8) ,
58672	 => std_logic_vector(to_unsigned(62,8) ,
58673	 => std_logic_vector(to_unsigned(65,8) ,
58674	 => std_logic_vector(to_unsigned(49,8) ,
58675	 => std_logic_vector(to_unsigned(46,8) ,
58676	 => std_logic_vector(to_unsigned(65,8) ,
58677	 => std_logic_vector(to_unsigned(51,8) ,
58678	 => std_logic_vector(to_unsigned(44,8) ,
58679	 => std_logic_vector(to_unsigned(32,8) ,
58680	 => std_logic_vector(to_unsigned(23,8) ,
58681	 => std_logic_vector(to_unsigned(40,8) ,
58682	 => std_logic_vector(to_unsigned(43,8) ,
58683	 => std_logic_vector(to_unsigned(55,8) ,
58684	 => std_logic_vector(to_unsigned(65,8) ,
58685	 => std_logic_vector(to_unsigned(64,8) ,
58686	 => std_logic_vector(to_unsigned(49,8) ,
58687	 => std_logic_vector(to_unsigned(72,8) ,
58688	 => std_logic_vector(to_unsigned(71,8) ,
58689	 => std_logic_vector(to_unsigned(63,8) ,
58690	 => std_logic_vector(to_unsigned(51,8) ,
58691	 => std_logic_vector(to_unsigned(37,8) ,
58692	 => std_logic_vector(to_unsigned(33,8) ,
58693	 => std_logic_vector(to_unsigned(21,8) ,
58694	 => std_logic_vector(to_unsigned(23,8) ,
58695	 => std_logic_vector(to_unsigned(27,8) ,
58696	 => std_logic_vector(to_unsigned(15,8) ,
58697	 => std_logic_vector(to_unsigned(19,8) ,
58698	 => std_logic_vector(to_unsigned(13,8) ,
58699	 => std_logic_vector(to_unsigned(9,8) ,
58700	 => std_logic_vector(to_unsigned(15,8) ,
58701	 => std_logic_vector(to_unsigned(13,8) ,
58702	 => std_logic_vector(to_unsigned(13,8) ,
58703	 => std_logic_vector(to_unsigned(10,8) ,
58704	 => std_logic_vector(to_unsigned(19,8) ,
58705	 => std_logic_vector(to_unsigned(45,8) ,
58706	 => std_logic_vector(to_unsigned(41,8) ,
58707	 => std_logic_vector(to_unsigned(14,8) ,
58708	 => std_logic_vector(to_unsigned(8,8) ,
58709	 => std_logic_vector(to_unsigned(41,8) ,
58710	 => std_logic_vector(to_unsigned(72,8) ,
58711	 => std_logic_vector(to_unsigned(17,8) ,
58712	 => std_logic_vector(to_unsigned(27,8) ,
58713	 => std_logic_vector(to_unsigned(46,8) ,
58714	 => std_logic_vector(to_unsigned(30,8) ,
58715	 => std_logic_vector(to_unsigned(24,8) ,
58716	 => std_logic_vector(to_unsigned(27,8) ,
58717	 => std_logic_vector(to_unsigned(27,8) ,
58718	 => std_logic_vector(to_unsigned(29,8) ,
58719	 => std_logic_vector(to_unsigned(16,8) ,
58720	 => std_logic_vector(to_unsigned(34,8) ,
58721	 => std_logic_vector(to_unsigned(141,8) ,
58722	 => std_logic_vector(to_unsigned(144,8) ,
58723	 => std_logic_vector(to_unsigned(141,8) ,
58724	 => std_logic_vector(to_unsigned(139,8) ,
58725	 => std_logic_vector(to_unsigned(142,8) ,
58726	 => std_logic_vector(to_unsigned(152,8) ,
58727	 => std_logic_vector(to_unsigned(43,8) ,
58728	 => std_logic_vector(to_unsigned(32,8) ,
58729	 => std_logic_vector(to_unsigned(85,8) ,
58730	 => std_logic_vector(to_unsigned(74,8) ,
58731	 => std_logic_vector(to_unsigned(18,8) ,
58732	 => std_logic_vector(to_unsigned(9,8) ,
58733	 => std_logic_vector(to_unsigned(11,8) ,
58734	 => std_logic_vector(to_unsigned(11,8) ,
58735	 => std_logic_vector(to_unsigned(12,8) ,
58736	 => std_logic_vector(to_unsigned(11,8) ,
58737	 => std_logic_vector(to_unsigned(10,8) ,
58738	 => std_logic_vector(to_unsigned(12,8) ,
58739	 => std_logic_vector(to_unsigned(8,8) ,
58740	 => std_logic_vector(to_unsigned(8,8) ,
58741	 => std_logic_vector(to_unsigned(9,8) ,
58742	 => std_logic_vector(to_unsigned(8,8) ,
58743	 => std_logic_vector(to_unsigned(9,8) ,
58744	 => std_logic_vector(to_unsigned(9,8) ,
58745	 => std_logic_vector(to_unsigned(6,8) ,
58746	 => std_logic_vector(to_unsigned(10,8) ,
58747	 => std_logic_vector(to_unsigned(10,8) ,
58748	 => std_logic_vector(to_unsigned(25,8) ,
58749	 => std_logic_vector(to_unsigned(32,8) ,
58750	 => std_logic_vector(to_unsigned(15,8) ,
58751	 => std_logic_vector(to_unsigned(24,8) ,
58752	 => std_logic_vector(to_unsigned(26,8) ,
58753	 => std_logic_vector(to_unsigned(38,8) ,
58754	 => std_logic_vector(to_unsigned(64,8) ,
58755	 => std_logic_vector(to_unsigned(65,8) ,
58756	 => std_logic_vector(to_unsigned(37,8) ,
58757	 => std_logic_vector(to_unsigned(32,8) ,
58758	 => std_logic_vector(to_unsigned(39,8) ,
58759	 => std_logic_vector(to_unsigned(27,8) ,
58760	 => std_logic_vector(to_unsigned(16,8) ,
58761	 => std_logic_vector(to_unsigned(28,8) ,
58762	 => std_logic_vector(to_unsigned(37,8) ,
58763	 => std_logic_vector(to_unsigned(25,8) ,
58764	 => std_logic_vector(to_unsigned(24,8) ,
58765	 => std_logic_vector(to_unsigned(30,8) ,
58766	 => std_logic_vector(to_unsigned(45,8) ,
58767	 => std_logic_vector(to_unsigned(35,8) ,
58768	 => std_logic_vector(to_unsigned(18,8) ,
58769	 => std_logic_vector(to_unsigned(17,8) ,
58770	 => std_logic_vector(to_unsigned(16,8) ,
58771	 => std_logic_vector(to_unsigned(14,8) ,
58772	 => std_logic_vector(to_unsigned(6,8) ,
58773	 => std_logic_vector(to_unsigned(6,8) ,
58774	 => std_logic_vector(to_unsigned(18,8) ,
58775	 => std_logic_vector(to_unsigned(15,8) ,
58776	 => std_logic_vector(to_unsigned(26,8) ,
58777	 => std_logic_vector(to_unsigned(27,8) ,
58778	 => std_logic_vector(to_unsigned(21,8) ,
58779	 => std_logic_vector(to_unsigned(18,8) ,
58780	 => std_logic_vector(to_unsigned(19,8) ,
58781	 => std_logic_vector(to_unsigned(25,8) ,
58782	 => std_logic_vector(to_unsigned(31,8) ,
58783	 => std_logic_vector(to_unsigned(35,8) ,
58784	 => std_logic_vector(to_unsigned(30,8) ,
58785	 => std_logic_vector(to_unsigned(20,8) ,
58786	 => std_logic_vector(to_unsigned(14,8) ,
58787	 => std_logic_vector(to_unsigned(12,8) ,
58788	 => std_logic_vector(to_unsigned(12,8) ,
58789	 => std_logic_vector(to_unsigned(12,8) ,
58790	 => std_logic_vector(to_unsigned(15,8) ,
58791	 => std_logic_vector(to_unsigned(15,8) ,
58792	 => std_logic_vector(to_unsigned(17,8) ,
58793	 => std_logic_vector(to_unsigned(12,8) ,
58794	 => std_logic_vector(to_unsigned(14,8) ,
58795	 => std_logic_vector(to_unsigned(18,8) ,
58796	 => std_logic_vector(to_unsigned(31,8) ,
58797	 => std_logic_vector(to_unsigned(35,8) ,
58798	 => std_logic_vector(to_unsigned(38,8) ,
58799	 => std_logic_vector(to_unsigned(45,8) ,
58800	 => std_logic_vector(to_unsigned(51,8) ,
58801	 => std_logic_vector(to_unsigned(63,8) ,
58802	 => std_logic_vector(to_unsigned(56,8) ,
58803	 => std_logic_vector(to_unsigned(43,8) ,
58804	 => std_logic_vector(to_unsigned(43,8) ,
58805	 => std_logic_vector(to_unsigned(41,8) ,
58806	 => std_logic_vector(to_unsigned(45,8) ,
58807	 => std_logic_vector(to_unsigned(45,8) ,
58808	 => std_logic_vector(to_unsigned(35,8) ,
58809	 => std_logic_vector(to_unsigned(32,8) ,
58810	 => std_logic_vector(to_unsigned(76,8) ,
58811	 => std_logic_vector(to_unsigned(90,8) ,
58812	 => std_logic_vector(to_unsigned(57,8) ,
58813	 => std_logic_vector(to_unsigned(20,8) ,
58814	 => std_logic_vector(to_unsigned(12,8) ,
58815	 => std_logic_vector(to_unsigned(5,8) ,
58816	 => std_logic_vector(to_unsigned(6,8) ,
58817	 => std_logic_vector(to_unsigned(6,8) ,
58818	 => std_logic_vector(to_unsigned(8,8) ,
58819	 => std_logic_vector(to_unsigned(16,8) ,
58820	 => std_logic_vector(to_unsigned(10,8) ,
58821	 => std_logic_vector(to_unsigned(6,8) ,
58822	 => std_logic_vector(to_unsigned(12,8) ,
58823	 => std_logic_vector(to_unsigned(9,8) ,
58824	 => std_logic_vector(to_unsigned(0,8) ,
58825	 => std_logic_vector(to_unsigned(2,8) ,
58826	 => std_logic_vector(to_unsigned(14,8) ,
58827	 => std_logic_vector(to_unsigned(28,8) ,
58828	 => std_logic_vector(to_unsigned(45,8) ,
58829	 => std_logic_vector(to_unsigned(57,8) ,
58830	 => std_logic_vector(to_unsigned(35,8) ,
58831	 => std_logic_vector(to_unsigned(25,8) ,
58832	 => std_logic_vector(to_unsigned(27,8) ,
58833	 => std_logic_vector(to_unsigned(17,8) ,
58834	 => std_logic_vector(to_unsigned(17,8) ,
58835	 => std_logic_vector(to_unsigned(18,8) ,
58836	 => std_logic_vector(to_unsigned(14,8) ,
58837	 => std_logic_vector(to_unsigned(10,8) ,
58838	 => std_logic_vector(to_unsigned(9,8) ,
58839	 => std_logic_vector(to_unsigned(7,8) ,
58840	 => std_logic_vector(to_unsigned(5,8) ,
58841	 => std_logic_vector(to_unsigned(6,8) ,
58842	 => std_logic_vector(to_unsigned(2,8) ,
58843	 => std_logic_vector(to_unsigned(0,8) ,
58844	 => std_logic_vector(to_unsigned(1,8) ,
58845	 => std_logic_vector(to_unsigned(0,8) ,
58846	 => std_logic_vector(to_unsigned(0,8) ,
58847	 => std_logic_vector(to_unsigned(2,8) ,
58848	 => std_logic_vector(to_unsigned(11,8) ,
58849	 => std_logic_vector(to_unsigned(10,8) ,
58850	 => std_logic_vector(to_unsigned(3,8) ,
58851	 => std_logic_vector(to_unsigned(2,8) ,
58852	 => std_logic_vector(to_unsigned(3,8) ,
58853	 => std_logic_vector(to_unsigned(7,8) ,
58854	 => std_logic_vector(to_unsigned(8,8) ,
58855	 => std_logic_vector(to_unsigned(9,8) ,
58856	 => std_logic_vector(to_unsigned(10,8) ,
58857	 => std_logic_vector(to_unsigned(7,8) ,
58858	 => std_logic_vector(to_unsigned(12,8) ,
58859	 => std_logic_vector(to_unsigned(17,8) ,
58860	 => std_logic_vector(to_unsigned(16,8) ,
58861	 => std_logic_vector(to_unsigned(14,8) ,
58862	 => std_logic_vector(to_unsigned(10,8) ,
58863	 => std_logic_vector(to_unsigned(8,8) ,
58864	 => std_logic_vector(to_unsigned(14,8) ,
58865	 => std_logic_vector(to_unsigned(12,8) ,
58866	 => std_logic_vector(to_unsigned(12,8) ,
58867	 => std_logic_vector(to_unsigned(12,8) ,
58868	 => std_logic_vector(to_unsigned(9,8) ,
58869	 => std_logic_vector(to_unsigned(6,8) ,
58870	 => std_logic_vector(to_unsigned(4,8) ,
58871	 => std_logic_vector(to_unsigned(7,8) ,
58872	 => std_logic_vector(to_unsigned(8,8) ,
58873	 => std_logic_vector(to_unsigned(5,8) ,
58874	 => std_logic_vector(to_unsigned(6,8) ,
58875	 => std_logic_vector(to_unsigned(13,8) ,
58876	 => std_logic_vector(to_unsigned(20,8) ,
58877	 => std_logic_vector(to_unsigned(8,8) ,
58878	 => std_logic_vector(to_unsigned(4,8) ,
58879	 => std_logic_vector(to_unsigned(9,8) ,
58880	 => std_logic_vector(to_unsigned(8,8) ,
58881	 => std_logic_vector(to_unsigned(88,8) ,
58882	 => std_logic_vector(to_unsigned(91,8) ,
58883	 => std_logic_vector(to_unsigned(68,8) ,
58884	 => std_logic_vector(to_unsigned(79,8) ,
58885	 => std_logic_vector(to_unsigned(74,8) ,
58886	 => std_logic_vector(to_unsigned(47,8) ,
58887	 => std_logic_vector(to_unsigned(27,8) ,
58888	 => std_logic_vector(to_unsigned(43,8) ,
58889	 => std_logic_vector(to_unsigned(63,8) ,
58890	 => std_logic_vector(to_unsigned(59,8) ,
58891	 => std_logic_vector(to_unsigned(63,8) ,
58892	 => std_logic_vector(to_unsigned(45,8) ,
58893	 => std_logic_vector(to_unsigned(48,8) ,
58894	 => std_logic_vector(to_unsigned(92,8) ,
58895	 => std_logic_vector(to_unsigned(88,8) ,
58896	 => std_logic_vector(to_unsigned(61,8) ,
58897	 => std_logic_vector(to_unsigned(79,8) ,
58898	 => std_logic_vector(to_unsigned(77,8) ,
58899	 => std_logic_vector(to_unsigned(65,8) ,
58900	 => std_logic_vector(to_unsigned(68,8) ,
58901	 => std_logic_vector(to_unsigned(49,8) ,
58902	 => std_logic_vector(to_unsigned(35,8) ,
58903	 => std_logic_vector(to_unsigned(33,8) ,
58904	 => std_logic_vector(to_unsigned(45,8) ,
58905	 => std_logic_vector(to_unsigned(77,8) ,
58906	 => std_logic_vector(to_unsigned(58,8) ,
58907	 => std_logic_vector(to_unsigned(60,8) ,
58908	 => std_logic_vector(to_unsigned(54,8) ,
58909	 => std_logic_vector(to_unsigned(46,8) ,
58910	 => std_logic_vector(to_unsigned(40,8) ,
58911	 => std_logic_vector(to_unsigned(38,8) ,
58912	 => std_logic_vector(to_unsigned(65,8) ,
58913	 => std_logic_vector(to_unsigned(74,8) ,
58914	 => std_logic_vector(to_unsigned(72,8) ,
58915	 => std_logic_vector(to_unsigned(50,8) ,
58916	 => std_logic_vector(to_unsigned(35,8) ,
58917	 => std_logic_vector(to_unsigned(34,8) ,
58918	 => std_logic_vector(to_unsigned(22,8) ,
58919	 => std_logic_vector(to_unsigned(39,8) ,
58920	 => std_logic_vector(to_unsigned(53,8) ,
58921	 => std_logic_vector(to_unsigned(51,8) ,
58922	 => std_logic_vector(to_unsigned(59,8) ,
58923	 => std_logic_vector(to_unsigned(68,8) ,
58924	 => std_logic_vector(to_unsigned(64,8) ,
58925	 => std_logic_vector(to_unsigned(51,8) ,
58926	 => std_logic_vector(to_unsigned(63,8) ,
58927	 => std_logic_vector(to_unsigned(66,8) ,
58928	 => std_logic_vector(to_unsigned(66,8) ,
58929	 => std_logic_vector(to_unsigned(74,8) ,
58930	 => std_logic_vector(to_unsigned(72,8) ,
58931	 => std_logic_vector(to_unsigned(85,8) ,
58932	 => std_logic_vector(to_unsigned(88,8) ,
58933	 => std_logic_vector(to_unsigned(91,8) ,
58934	 => std_logic_vector(to_unsigned(67,8) ,
58935	 => std_logic_vector(to_unsigned(84,8) ,
58936	 => std_logic_vector(to_unsigned(107,8) ,
58937	 => std_logic_vector(to_unsigned(90,8) ,
58938	 => std_logic_vector(to_unsigned(51,8) ,
58939	 => std_logic_vector(to_unsigned(48,8) ,
58940	 => std_logic_vector(to_unsigned(45,8) ,
58941	 => std_logic_vector(to_unsigned(23,8) ,
58942	 => std_logic_vector(to_unsigned(19,8) ,
58943	 => std_logic_vector(to_unsigned(55,8) ,
58944	 => std_logic_vector(to_unsigned(56,8) ,
58945	 => std_logic_vector(to_unsigned(56,8) ,
58946	 => std_logic_vector(to_unsigned(97,8) ,
58947	 => std_logic_vector(to_unsigned(80,8) ,
58948	 => std_logic_vector(to_unsigned(103,8) ,
58949	 => std_logic_vector(to_unsigned(84,8) ,
58950	 => std_logic_vector(to_unsigned(72,8) ,
58951	 => std_logic_vector(to_unsigned(114,8) ,
58952	 => std_logic_vector(to_unsigned(95,8) ,
58953	 => std_logic_vector(to_unsigned(91,8) ,
58954	 => std_logic_vector(to_unsigned(130,8) ,
58955	 => std_logic_vector(to_unsigned(144,8) ,
58956	 => std_logic_vector(to_unsigned(138,8) ,
58957	 => std_logic_vector(to_unsigned(125,8) ,
58958	 => std_logic_vector(to_unsigned(119,8) ,
58959	 => std_logic_vector(to_unsigned(112,8) ,
58960	 => std_logic_vector(to_unsigned(118,8) ,
58961	 => std_logic_vector(to_unsigned(125,8) ,
58962	 => std_logic_vector(to_unsigned(119,8) ,
58963	 => std_logic_vector(to_unsigned(111,8) ,
58964	 => std_logic_vector(to_unsigned(109,8) ,
58965	 => std_logic_vector(to_unsigned(127,8) ,
58966	 => std_logic_vector(to_unsigned(91,8) ,
58967	 => std_logic_vector(to_unsigned(30,8) ,
58968	 => std_logic_vector(to_unsigned(30,8) ,
58969	 => std_logic_vector(to_unsigned(34,8) ,
58970	 => std_logic_vector(to_unsigned(30,8) ,
58971	 => std_logic_vector(to_unsigned(39,8) ,
58972	 => std_logic_vector(to_unsigned(43,8) ,
58973	 => std_logic_vector(to_unsigned(48,8) ,
58974	 => std_logic_vector(to_unsigned(51,8) ,
58975	 => std_logic_vector(to_unsigned(51,8) ,
58976	 => std_logic_vector(to_unsigned(55,8) ,
58977	 => std_logic_vector(to_unsigned(61,8) ,
58978	 => std_logic_vector(to_unsigned(62,8) ,
58979	 => std_logic_vector(to_unsigned(69,8) ,
58980	 => std_logic_vector(to_unsigned(61,8) ,
58981	 => std_logic_vector(to_unsigned(55,8) ,
58982	 => std_logic_vector(to_unsigned(59,8) ,
58983	 => std_logic_vector(to_unsigned(61,8) ,
58984	 => std_logic_vector(to_unsigned(53,8) ,
58985	 => std_logic_vector(to_unsigned(51,8) ,
58986	 => std_logic_vector(to_unsigned(48,8) ,
58987	 => std_logic_vector(to_unsigned(93,8) ,
58988	 => std_logic_vector(to_unsigned(100,8) ,
58989	 => std_logic_vector(to_unsigned(52,8) ,
58990	 => std_logic_vector(to_unsigned(55,8) ,
58991	 => std_logic_vector(to_unsigned(55,8) ,
58992	 => std_logic_vector(to_unsigned(61,8) ,
58993	 => std_logic_vector(to_unsigned(66,8) ,
58994	 => std_logic_vector(to_unsigned(46,8) ,
58995	 => std_logic_vector(to_unsigned(48,8) ,
58996	 => std_logic_vector(to_unsigned(60,8) ,
58997	 => std_logic_vector(to_unsigned(47,8) ,
58998	 => std_logic_vector(to_unsigned(41,8) ,
58999	 => std_logic_vector(to_unsigned(28,8) ,
59000	 => std_logic_vector(to_unsigned(29,8) ,
59001	 => std_logic_vector(to_unsigned(37,8) ,
59002	 => std_logic_vector(to_unsigned(22,8) ,
59003	 => std_logic_vector(to_unsigned(19,8) ,
59004	 => std_logic_vector(to_unsigned(20,8) ,
59005	 => std_logic_vector(to_unsigned(22,8) ,
59006	 => std_logic_vector(to_unsigned(22,8) ,
59007	 => std_logic_vector(to_unsigned(35,8) ,
59008	 => std_logic_vector(to_unsigned(52,8) ,
59009	 => std_logic_vector(to_unsigned(79,8) ,
59010	 => std_logic_vector(to_unsigned(57,8) ,
59011	 => std_logic_vector(to_unsigned(33,8) ,
59012	 => std_logic_vector(to_unsigned(33,8) ,
59013	 => std_logic_vector(to_unsigned(39,8) ,
59014	 => std_logic_vector(to_unsigned(48,8) ,
59015	 => std_logic_vector(to_unsigned(29,8) ,
59016	 => std_logic_vector(to_unsigned(18,8) ,
59017	 => std_logic_vector(to_unsigned(15,8) ,
59018	 => std_logic_vector(to_unsigned(11,8) ,
59019	 => std_logic_vector(to_unsigned(12,8) ,
59020	 => std_logic_vector(to_unsigned(14,8) ,
59021	 => std_logic_vector(to_unsigned(10,8) ,
59022	 => std_logic_vector(to_unsigned(12,8) ,
59023	 => std_logic_vector(to_unsigned(18,8) ,
59024	 => std_logic_vector(to_unsigned(16,8) ,
59025	 => std_logic_vector(to_unsigned(14,8) ,
59026	 => std_logic_vector(to_unsigned(20,8) ,
59027	 => std_logic_vector(to_unsigned(18,8) ,
59028	 => std_logic_vector(to_unsigned(22,8) ,
59029	 => std_logic_vector(to_unsigned(48,8) ,
59030	 => std_logic_vector(to_unsigned(46,8) ,
59031	 => std_logic_vector(to_unsigned(15,8) ,
59032	 => std_logic_vector(to_unsigned(28,8) ,
59033	 => std_logic_vector(to_unsigned(39,8) ,
59034	 => std_logic_vector(to_unsigned(56,8) ,
59035	 => std_logic_vector(to_unsigned(20,8) ,
59036	 => std_logic_vector(to_unsigned(7,8) ,
59037	 => std_logic_vector(to_unsigned(13,8) ,
59038	 => std_logic_vector(to_unsigned(18,8) ,
59039	 => std_logic_vector(to_unsigned(4,8) ,
59040	 => std_logic_vector(to_unsigned(23,8) ,
59041	 => std_logic_vector(to_unsigned(114,8) ,
59042	 => std_logic_vector(to_unsigned(69,8) ,
59043	 => std_logic_vector(to_unsigned(99,8) ,
59044	 => std_logic_vector(to_unsigned(99,8) ,
59045	 => std_logic_vector(to_unsigned(131,8) ,
59046	 => std_logic_vector(to_unsigned(108,8) ,
59047	 => std_logic_vector(to_unsigned(23,8) ,
59048	 => std_logic_vector(to_unsigned(28,8) ,
59049	 => std_logic_vector(to_unsigned(84,8) ,
59050	 => std_logic_vector(to_unsigned(76,8) ,
59051	 => std_logic_vector(to_unsigned(30,8) ,
59052	 => std_logic_vector(to_unsigned(16,8) ,
59053	 => std_logic_vector(to_unsigned(13,8) ,
59054	 => std_logic_vector(to_unsigned(10,8) ,
59055	 => std_logic_vector(to_unsigned(9,8) ,
59056	 => std_logic_vector(to_unsigned(6,8) ,
59057	 => std_logic_vector(to_unsigned(9,8) ,
59058	 => std_logic_vector(to_unsigned(10,8) ,
59059	 => std_logic_vector(to_unsigned(11,8) ,
59060	 => std_logic_vector(to_unsigned(9,8) ,
59061	 => std_logic_vector(to_unsigned(11,8) ,
59062	 => std_logic_vector(to_unsigned(11,8) ,
59063	 => std_logic_vector(to_unsigned(11,8) ,
59064	 => std_logic_vector(to_unsigned(12,8) ,
59065	 => std_logic_vector(to_unsigned(10,8) ,
59066	 => std_logic_vector(to_unsigned(11,8) ,
59067	 => std_logic_vector(to_unsigned(22,8) ,
59068	 => std_logic_vector(to_unsigned(27,8) ,
59069	 => std_logic_vector(to_unsigned(23,8) ,
59070	 => std_logic_vector(to_unsigned(22,8) ,
59071	 => std_logic_vector(to_unsigned(22,8) ,
59072	 => std_logic_vector(to_unsigned(23,8) ,
59073	 => std_logic_vector(to_unsigned(25,8) ,
59074	 => std_logic_vector(to_unsigned(34,8) ,
59075	 => std_logic_vector(to_unsigned(30,8) ,
59076	 => std_logic_vector(to_unsigned(23,8) ,
59077	 => std_logic_vector(to_unsigned(29,8) ,
59078	 => std_logic_vector(to_unsigned(29,8) ,
59079	 => std_logic_vector(to_unsigned(24,8) ,
59080	 => std_logic_vector(to_unsigned(20,8) ,
59081	 => std_logic_vector(to_unsigned(33,8) ,
59082	 => std_logic_vector(to_unsigned(39,8) ,
59083	 => std_logic_vector(to_unsigned(29,8) ,
59084	 => std_logic_vector(to_unsigned(20,8) ,
59085	 => std_logic_vector(to_unsigned(29,8) ,
59086	 => std_logic_vector(to_unsigned(33,8) ,
59087	 => std_logic_vector(to_unsigned(37,8) ,
59088	 => std_logic_vector(to_unsigned(30,8) ,
59089	 => std_logic_vector(to_unsigned(19,8) ,
59090	 => std_logic_vector(to_unsigned(16,8) ,
59091	 => std_logic_vector(to_unsigned(13,8) ,
59092	 => std_logic_vector(to_unsigned(10,8) ,
59093	 => std_logic_vector(to_unsigned(11,8) ,
59094	 => std_logic_vector(to_unsigned(14,8) ,
59095	 => std_logic_vector(to_unsigned(16,8) ,
59096	 => std_logic_vector(to_unsigned(21,8) ,
59097	 => std_logic_vector(to_unsigned(26,8) ,
59098	 => std_logic_vector(to_unsigned(16,8) ,
59099	 => std_logic_vector(to_unsigned(14,8) ,
59100	 => std_logic_vector(to_unsigned(23,8) ,
59101	 => std_logic_vector(to_unsigned(24,8) ,
59102	 => std_logic_vector(to_unsigned(28,8) ,
59103	 => std_logic_vector(to_unsigned(35,8) ,
59104	 => std_logic_vector(to_unsigned(37,8) ,
59105	 => std_logic_vector(to_unsigned(27,8) ,
59106	 => std_logic_vector(to_unsigned(23,8) ,
59107	 => std_logic_vector(to_unsigned(19,8) ,
59108	 => std_logic_vector(to_unsigned(13,8) ,
59109	 => std_logic_vector(to_unsigned(12,8) ,
59110	 => std_logic_vector(to_unsigned(13,8) ,
59111	 => std_logic_vector(to_unsigned(19,8) ,
59112	 => std_logic_vector(to_unsigned(29,8) ,
59113	 => std_logic_vector(to_unsigned(14,8) ,
59114	 => std_logic_vector(to_unsigned(7,8) ,
59115	 => std_logic_vector(to_unsigned(19,8) ,
59116	 => std_logic_vector(to_unsigned(35,8) ,
59117	 => std_logic_vector(to_unsigned(30,8) ,
59118	 => std_logic_vector(to_unsigned(68,8) ,
59119	 => std_logic_vector(to_unsigned(84,8) ,
59120	 => std_logic_vector(to_unsigned(59,8) ,
59121	 => std_logic_vector(to_unsigned(35,8) ,
59122	 => std_logic_vector(to_unsigned(35,8) ,
59123	 => std_logic_vector(to_unsigned(48,8) ,
59124	 => std_logic_vector(to_unsigned(51,8) ,
59125	 => std_logic_vector(to_unsigned(49,8) ,
59126	 => std_logic_vector(to_unsigned(55,8) ,
59127	 => std_logic_vector(to_unsigned(48,8) ,
59128	 => std_logic_vector(to_unsigned(32,8) ,
59129	 => std_logic_vector(to_unsigned(55,8) ,
59130	 => std_logic_vector(to_unsigned(84,8) ,
59131	 => std_logic_vector(to_unsigned(78,8) ,
59132	 => std_logic_vector(to_unsigned(24,8) ,
59133	 => std_logic_vector(to_unsigned(16,8) ,
59134	 => std_logic_vector(to_unsigned(11,8) ,
59135	 => std_logic_vector(to_unsigned(5,8) ,
59136	 => std_logic_vector(to_unsigned(8,8) ,
59137	 => std_logic_vector(to_unsigned(13,8) ,
59138	 => std_logic_vector(to_unsigned(22,8) ,
59139	 => std_logic_vector(to_unsigned(17,8) ,
59140	 => std_logic_vector(to_unsigned(12,8) ,
59141	 => std_logic_vector(to_unsigned(15,8) ,
59142	 => std_logic_vector(to_unsigned(18,8) ,
59143	 => std_logic_vector(to_unsigned(10,8) ,
59144	 => std_logic_vector(to_unsigned(1,8) ,
59145	 => std_logic_vector(to_unsigned(1,8) ,
59146	 => std_logic_vector(to_unsigned(3,8) ,
59147	 => std_logic_vector(to_unsigned(19,8) ,
59148	 => std_logic_vector(to_unsigned(23,8) ,
59149	 => std_logic_vector(to_unsigned(20,8) ,
59150	 => std_logic_vector(to_unsigned(25,8) ,
59151	 => std_logic_vector(to_unsigned(14,8) ,
59152	 => std_logic_vector(to_unsigned(16,8) ,
59153	 => std_logic_vector(to_unsigned(12,8) ,
59154	 => std_logic_vector(to_unsigned(12,8) ,
59155	 => std_logic_vector(to_unsigned(13,8) ,
59156	 => std_logic_vector(to_unsigned(13,8) ,
59157	 => std_logic_vector(to_unsigned(10,8) ,
59158	 => std_logic_vector(to_unsigned(7,8) ,
59159	 => std_logic_vector(to_unsigned(8,8) ,
59160	 => std_logic_vector(to_unsigned(7,8) ,
59161	 => std_logic_vector(to_unsigned(6,8) ,
59162	 => std_logic_vector(to_unsigned(7,8) ,
59163	 => std_logic_vector(to_unsigned(2,8) ,
59164	 => std_logic_vector(to_unsigned(0,8) ,
59165	 => std_logic_vector(to_unsigned(0,8) ,
59166	 => std_logic_vector(to_unsigned(0,8) ,
59167	 => std_logic_vector(to_unsigned(2,8) ,
59168	 => std_logic_vector(to_unsigned(4,8) ,
59169	 => std_logic_vector(to_unsigned(1,8) ,
59170	 => std_logic_vector(to_unsigned(0,8) ,
59171	 => std_logic_vector(to_unsigned(1,8) ,
59172	 => std_logic_vector(to_unsigned(2,8) ,
59173	 => std_logic_vector(to_unsigned(7,8) ,
59174	 => std_logic_vector(to_unsigned(8,8) ,
59175	 => std_logic_vector(to_unsigned(7,8) ,
59176	 => std_logic_vector(to_unsigned(5,8) ,
59177	 => std_logic_vector(to_unsigned(5,8) ,
59178	 => std_logic_vector(to_unsigned(8,8) ,
59179	 => std_logic_vector(to_unsigned(8,8) ,
59180	 => std_logic_vector(to_unsigned(10,8) ,
59181	 => std_logic_vector(to_unsigned(10,8) ,
59182	 => std_logic_vector(to_unsigned(10,8) ,
59183	 => std_logic_vector(to_unsigned(10,8) ,
59184	 => std_logic_vector(to_unsigned(19,8) ,
59185	 => std_logic_vector(to_unsigned(20,8) ,
59186	 => std_logic_vector(to_unsigned(13,8) ,
59187	 => std_logic_vector(to_unsigned(11,8) ,
59188	 => std_logic_vector(to_unsigned(10,8) ,
59189	 => std_logic_vector(to_unsigned(6,8) ,
59190	 => std_logic_vector(to_unsigned(4,8) ,
59191	 => std_logic_vector(to_unsigned(5,8) ,
59192	 => std_logic_vector(to_unsigned(8,8) ,
59193	 => std_logic_vector(to_unsigned(9,8) ,
59194	 => std_logic_vector(to_unsigned(9,8) ,
59195	 => std_logic_vector(to_unsigned(8,8) ,
59196	 => std_logic_vector(to_unsigned(13,8) ,
59197	 => std_logic_vector(to_unsigned(9,8) ,
59198	 => std_logic_vector(to_unsigned(6,8) ,
59199	 => std_logic_vector(to_unsigned(10,8) ,
59200	 => std_logic_vector(to_unsigned(10,8) ,
59201	 => std_logic_vector(to_unsigned(81,8) ,
59202	 => std_logic_vector(to_unsigned(88,8) ,
59203	 => std_logic_vector(to_unsigned(71,8) ,
59204	 => std_logic_vector(to_unsigned(74,8) ,
59205	 => std_logic_vector(to_unsigned(72,8) ,
59206	 => std_logic_vector(to_unsigned(52,8) ,
59207	 => std_logic_vector(to_unsigned(35,8) ,
59208	 => std_logic_vector(to_unsigned(47,8) ,
59209	 => std_logic_vector(to_unsigned(57,8) ,
59210	 => std_logic_vector(to_unsigned(56,8) ,
59211	 => std_logic_vector(to_unsigned(70,8) ,
59212	 => std_logic_vector(to_unsigned(60,8) ,
59213	 => std_logic_vector(to_unsigned(62,8) ,
59214	 => std_logic_vector(to_unsigned(93,8) ,
59215	 => std_logic_vector(to_unsigned(93,8) ,
59216	 => std_logic_vector(to_unsigned(57,8) ,
59217	 => std_logic_vector(to_unsigned(80,8) ,
59218	 => std_logic_vector(to_unsigned(65,8) ,
59219	 => std_logic_vector(to_unsigned(41,8) ,
59220	 => std_logic_vector(to_unsigned(58,8) ,
59221	 => std_logic_vector(to_unsigned(41,8) ,
59222	 => std_logic_vector(to_unsigned(30,8) ,
59223	 => std_logic_vector(to_unsigned(26,8) ,
59224	 => std_logic_vector(to_unsigned(32,8) ,
59225	 => std_logic_vector(to_unsigned(76,8) ,
59226	 => std_logic_vector(to_unsigned(77,8) ,
59227	 => std_logic_vector(to_unsigned(61,8) ,
59228	 => std_logic_vector(to_unsigned(48,8) ,
59229	 => std_logic_vector(to_unsigned(58,8) ,
59230	 => std_logic_vector(to_unsigned(71,8) ,
59231	 => std_logic_vector(to_unsigned(47,8) ,
59232	 => std_logic_vector(to_unsigned(29,8) ,
59233	 => std_logic_vector(to_unsigned(27,8) ,
59234	 => std_logic_vector(to_unsigned(25,8) ,
59235	 => std_logic_vector(to_unsigned(17,8) ,
59236	 => std_logic_vector(to_unsigned(15,8) ,
59237	 => std_logic_vector(to_unsigned(42,8) ,
59238	 => std_logic_vector(to_unsigned(45,8) ,
59239	 => std_logic_vector(to_unsigned(38,8) ,
59240	 => std_logic_vector(to_unsigned(55,8) ,
59241	 => std_logic_vector(to_unsigned(57,8) ,
59242	 => std_logic_vector(to_unsigned(72,8) ,
59243	 => std_logic_vector(to_unsigned(80,8) ,
59244	 => std_logic_vector(to_unsigned(68,8) ,
59245	 => std_logic_vector(to_unsigned(78,8) ,
59246	 => std_logic_vector(to_unsigned(65,8) ,
59247	 => std_logic_vector(to_unsigned(61,8) ,
59248	 => std_logic_vector(to_unsigned(67,8) ,
59249	 => std_logic_vector(to_unsigned(58,8) ,
59250	 => std_logic_vector(to_unsigned(58,8) ,
59251	 => std_logic_vector(to_unsigned(58,8) ,
59252	 => std_logic_vector(to_unsigned(68,8) ,
59253	 => std_logic_vector(to_unsigned(72,8) ,
59254	 => std_logic_vector(to_unsigned(43,8) ,
59255	 => std_logic_vector(to_unsigned(66,8) ,
59256	 => std_logic_vector(to_unsigned(87,8) ,
59257	 => std_logic_vector(to_unsigned(73,8) ,
59258	 => std_logic_vector(to_unsigned(41,8) ,
59259	 => std_logic_vector(to_unsigned(58,8) ,
59260	 => std_logic_vector(to_unsigned(80,8) ,
59261	 => std_logic_vector(to_unsigned(26,8) ,
59262	 => std_logic_vector(to_unsigned(20,8) ,
59263	 => std_logic_vector(to_unsigned(63,8) ,
59264	 => std_logic_vector(to_unsigned(69,8) ,
59265	 => std_logic_vector(to_unsigned(76,8) ,
59266	 => std_logic_vector(to_unsigned(93,8) ,
59267	 => std_logic_vector(to_unsigned(95,8) ,
59268	 => std_logic_vector(to_unsigned(101,8) ,
59269	 => std_logic_vector(to_unsigned(101,8) ,
59270	 => std_logic_vector(to_unsigned(103,8) ,
59271	 => std_logic_vector(to_unsigned(103,8) ,
59272	 => std_logic_vector(to_unsigned(84,8) ,
59273	 => std_logic_vector(to_unsigned(92,8) ,
59274	 => std_logic_vector(to_unsigned(134,8) ,
59275	 => std_logic_vector(to_unsigned(146,8) ,
59276	 => std_logic_vector(to_unsigned(131,8) ,
59277	 => std_logic_vector(to_unsigned(118,8) ,
59278	 => std_logic_vector(to_unsigned(122,8) ,
59279	 => std_logic_vector(to_unsigned(125,8) ,
59280	 => std_logic_vector(to_unsigned(130,8) ,
59281	 => std_logic_vector(to_unsigned(127,8) ,
59282	 => std_logic_vector(to_unsigned(108,8) ,
59283	 => std_logic_vector(to_unsigned(111,8) ,
59284	 => std_logic_vector(to_unsigned(111,8) ,
59285	 => std_logic_vector(to_unsigned(130,8) ,
59286	 => std_logic_vector(to_unsigned(95,8) ,
59287	 => std_logic_vector(to_unsigned(25,8) ,
59288	 => std_logic_vector(to_unsigned(33,8) ,
59289	 => std_logic_vector(to_unsigned(43,8) ,
59290	 => std_logic_vector(to_unsigned(46,8) ,
59291	 => std_logic_vector(to_unsigned(43,8) ,
59292	 => std_logic_vector(to_unsigned(38,8) ,
59293	 => std_logic_vector(to_unsigned(47,8) ,
59294	 => std_logic_vector(to_unsigned(44,8) ,
59295	 => std_logic_vector(to_unsigned(48,8) ,
59296	 => std_logic_vector(to_unsigned(54,8) ,
59297	 => std_logic_vector(to_unsigned(57,8) ,
59298	 => std_logic_vector(to_unsigned(57,8) ,
59299	 => std_logic_vector(to_unsigned(63,8) ,
59300	 => std_logic_vector(to_unsigned(58,8) ,
59301	 => std_logic_vector(to_unsigned(57,8) ,
59302	 => std_logic_vector(to_unsigned(82,8) ,
59303	 => std_logic_vector(to_unsigned(76,8) ,
59304	 => std_logic_vector(to_unsigned(60,8) ,
59305	 => std_logic_vector(to_unsigned(60,8) ,
59306	 => std_logic_vector(to_unsigned(84,8) ,
59307	 => std_logic_vector(to_unsigned(103,8) ,
59308	 => std_logic_vector(to_unsigned(66,8) ,
59309	 => std_logic_vector(to_unsigned(44,8) ,
59310	 => std_logic_vector(to_unsigned(46,8) ,
59311	 => std_logic_vector(to_unsigned(51,8) ,
59312	 => std_logic_vector(to_unsigned(64,8) ,
59313	 => std_logic_vector(to_unsigned(67,8) ,
59314	 => std_logic_vector(to_unsigned(44,8) ,
59315	 => std_logic_vector(to_unsigned(47,8) ,
59316	 => std_logic_vector(to_unsigned(57,8) ,
59317	 => std_logic_vector(to_unsigned(45,8) ,
59318	 => std_logic_vector(to_unsigned(38,8) ,
59319	 => std_logic_vector(to_unsigned(27,8) ,
59320	 => std_logic_vector(to_unsigned(37,8) ,
59321	 => std_logic_vector(to_unsigned(85,8) ,
59322	 => std_logic_vector(to_unsigned(78,8) ,
59323	 => std_logic_vector(to_unsigned(56,8) ,
59324	 => std_logic_vector(to_unsigned(58,8) ,
59325	 => std_logic_vector(to_unsigned(48,8) ,
59326	 => std_logic_vector(to_unsigned(30,8) ,
59327	 => std_logic_vector(to_unsigned(30,8) ,
59328	 => std_logic_vector(to_unsigned(21,8) ,
59329	 => std_logic_vector(to_unsigned(33,8) ,
59330	 => std_logic_vector(to_unsigned(53,8) ,
59331	 => std_logic_vector(to_unsigned(28,8) ,
59332	 => std_logic_vector(to_unsigned(32,8) ,
59333	 => std_logic_vector(to_unsigned(23,8) ,
59334	 => std_logic_vector(to_unsigned(32,8) ,
59335	 => std_logic_vector(to_unsigned(30,8) ,
59336	 => std_logic_vector(to_unsigned(10,8) ,
59337	 => std_logic_vector(to_unsigned(13,8) ,
59338	 => std_logic_vector(to_unsigned(17,8) ,
59339	 => std_logic_vector(to_unsigned(10,8) ,
59340	 => std_logic_vector(to_unsigned(10,8) ,
59341	 => std_logic_vector(to_unsigned(14,8) ,
59342	 => std_logic_vector(to_unsigned(15,8) ,
59343	 => std_logic_vector(to_unsigned(20,8) ,
59344	 => std_logic_vector(to_unsigned(16,8) ,
59345	 => std_logic_vector(to_unsigned(22,8) ,
59346	 => std_logic_vector(to_unsigned(30,8) ,
59347	 => std_logic_vector(to_unsigned(22,8) ,
59348	 => std_logic_vector(to_unsigned(17,8) ,
59349	 => std_logic_vector(to_unsigned(20,8) ,
59350	 => std_logic_vector(to_unsigned(101,8) ,
59351	 => std_logic_vector(to_unsigned(48,8) ,
59352	 => std_logic_vector(to_unsigned(23,8) ,
59353	 => std_logic_vector(to_unsigned(37,8) ,
59354	 => std_logic_vector(to_unsigned(51,8) ,
59355	 => std_logic_vector(to_unsigned(23,8) ,
59356	 => std_logic_vector(to_unsigned(10,8) ,
59357	 => std_logic_vector(to_unsigned(13,8) ,
59358	 => std_logic_vector(to_unsigned(15,8) ,
59359	 => std_logic_vector(to_unsigned(10,8) ,
59360	 => std_logic_vector(to_unsigned(30,8) ,
59361	 => std_logic_vector(to_unsigned(108,8) ,
59362	 => std_logic_vector(to_unsigned(42,8) ,
59363	 => std_logic_vector(to_unsigned(44,8) ,
59364	 => std_logic_vector(to_unsigned(61,8) ,
59365	 => std_logic_vector(to_unsigned(130,8) ,
59366	 => std_logic_vector(to_unsigned(66,8) ,
59367	 => std_logic_vector(to_unsigned(77,8) ,
59368	 => std_logic_vector(to_unsigned(54,8) ,
59369	 => std_logic_vector(to_unsigned(54,8) ,
59370	 => std_logic_vector(to_unsigned(81,8) ,
59371	 => std_logic_vector(to_unsigned(25,8) ,
59372	 => std_logic_vector(to_unsigned(22,8) ,
59373	 => std_logic_vector(to_unsigned(32,8) ,
59374	 => std_logic_vector(to_unsigned(26,8) ,
59375	 => std_logic_vector(to_unsigned(21,8) ,
59376	 => std_logic_vector(to_unsigned(17,8) ,
59377	 => std_logic_vector(to_unsigned(9,8) ,
59378	 => std_logic_vector(to_unsigned(6,8) ,
59379	 => std_logic_vector(to_unsigned(7,8) ,
59380	 => std_logic_vector(to_unsigned(8,8) ,
59381	 => std_logic_vector(to_unsigned(10,8) ,
59382	 => std_logic_vector(to_unsigned(8,8) ,
59383	 => std_logic_vector(to_unsigned(8,8) ,
59384	 => std_logic_vector(to_unsigned(10,8) ,
59385	 => std_logic_vector(to_unsigned(12,8) ,
59386	 => std_logic_vector(to_unsigned(11,8) ,
59387	 => std_logic_vector(to_unsigned(20,8) ,
59388	 => std_logic_vector(to_unsigned(24,8) ,
59389	 => std_logic_vector(to_unsigned(29,8) ,
59390	 => std_logic_vector(to_unsigned(35,8) ,
59391	 => std_logic_vector(to_unsigned(33,8) ,
59392	 => std_logic_vector(to_unsigned(35,8) ,
59393	 => std_logic_vector(to_unsigned(49,8) ,
59394	 => std_logic_vector(to_unsigned(57,8) ,
59395	 => std_logic_vector(to_unsigned(60,8) ,
59396	 => std_logic_vector(to_unsigned(37,8) ,
59397	 => std_logic_vector(to_unsigned(30,8) ,
59398	 => std_logic_vector(to_unsigned(27,8) ,
59399	 => std_logic_vector(to_unsigned(24,8) ,
59400	 => std_logic_vector(to_unsigned(23,8) ,
59401	 => std_logic_vector(to_unsigned(42,8) ,
59402	 => std_logic_vector(to_unsigned(55,8) ,
59403	 => std_logic_vector(to_unsigned(41,8) ,
59404	 => std_logic_vector(to_unsigned(22,8) ,
59405	 => std_logic_vector(to_unsigned(24,8) ,
59406	 => std_logic_vector(to_unsigned(41,8) ,
59407	 => std_logic_vector(to_unsigned(44,8) ,
59408	 => std_logic_vector(to_unsigned(37,8) ,
59409	 => std_logic_vector(to_unsigned(22,8) ,
59410	 => std_logic_vector(to_unsigned(13,8) ,
59411	 => std_logic_vector(to_unsigned(17,8) ,
59412	 => std_logic_vector(to_unsigned(13,8) ,
59413	 => std_logic_vector(to_unsigned(17,8) ,
59414	 => std_logic_vector(to_unsigned(21,8) ,
59415	 => std_logic_vector(to_unsigned(23,8) ,
59416	 => std_logic_vector(to_unsigned(24,8) ,
59417	 => std_logic_vector(to_unsigned(27,8) ,
59418	 => std_logic_vector(to_unsigned(18,8) ,
59419	 => std_logic_vector(to_unsigned(15,8) ,
59420	 => std_logic_vector(to_unsigned(18,8) ,
59421	 => std_logic_vector(to_unsigned(25,8) ,
59422	 => std_logic_vector(to_unsigned(23,8) ,
59423	 => std_logic_vector(to_unsigned(29,8) ,
59424	 => std_logic_vector(to_unsigned(25,8) ,
59425	 => std_logic_vector(to_unsigned(28,8) ,
59426	 => std_logic_vector(to_unsigned(38,8) ,
59427	 => std_logic_vector(to_unsigned(19,8) ,
59428	 => std_logic_vector(to_unsigned(11,8) ,
59429	 => std_logic_vector(to_unsigned(12,8) ,
59430	 => std_logic_vector(to_unsigned(17,8) ,
59431	 => std_logic_vector(to_unsigned(40,8) ,
59432	 => std_logic_vector(to_unsigned(36,8) ,
59433	 => std_logic_vector(to_unsigned(12,8) ,
59434	 => std_logic_vector(to_unsigned(14,8) ,
59435	 => std_logic_vector(to_unsigned(38,8) ,
59436	 => std_logic_vector(to_unsigned(30,8) ,
59437	 => std_logic_vector(to_unsigned(27,8) ,
59438	 => std_logic_vector(to_unsigned(32,8) ,
59439	 => std_logic_vector(to_unsigned(49,8) ,
59440	 => std_logic_vector(to_unsigned(54,8) ,
59441	 => std_logic_vector(to_unsigned(40,8) ,
59442	 => std_logic_vector(to_unsigned(37,8) ,
59443	 => std_logic_vector(to_unsigned(36,8) ,
59444	 => std_logic_vector(to_unsigned(40,8) ,
59445	 => std_logic_vector(to_unsigned(51,8) ,
59446	 => std_logic_vector(to_unsigned(43,8) ,
59447	 => std_logic_vector(to_unsigned(57,8) ,
59448	 => std_logic_vector(to_unsigned(85,8) ,
59449	 => std_logic_vector(to_unsigned(73,8) ,
59450	 => std_logic_vector(to_unsigned(54,8) ,
59451	 => std_logic_vector(to_unsigned(29,8) ,
59452	 => std_logic_vector(to_unsigned(26,8) ,
59453	 => std_logic_vector(to_unsigned(15,8) ,
59454	 => std_logic_vector(to_unsigned(9,8) ,
59455	 => std_logic_vector(to_unsigned(13,8) ,
59456	 => std_logic_vector(to_unsigned(12,8) ,
59457	 => std_logic_vector(to_unsigned(18,8) ,
59458	 => std_logic_vector(to_unsigned(18,8) ,
59459	 => std_logic_vector(to_unsigned(12,8) ,
59460	 => std_logic_vector(to_unsigned(14,8) ,
59461	 => std_logic_vector(to_unsigned(24,8) ,
59462	 => std_logic_vector(to_unsigned(30,8) ,
59463	 => std_logic_vector(to_unsigned(14,8) ,
59464	 => std_logic_vector(to_unsigned(2,8) ,
59465	 => std_logic_vector(to_unsigned(0,8) ,
59466	 => std_logic_vector(to_unsigned(2,8) ,
59467	 => std_logic_vector(to_unsigned(23,8) ,
59468	 => std_logic_vector(to_unsigned(47,8) ,
59469	 => std_logic_vector(to_unsigned(30,8) ,
59470	 => std_logic_vector(to_unsigned(14,8) ,
59471	 => std_logic_vector(to_unsigned(20,8) ,
59472	 => std_logic_vector(to_unsigned(29,8) ,
59473	 => std_logic_vector(to_unsigned(16,8) ,
59474	 => std_logic_vector(to_unsigned(8,8) ,
59475	 => std_logic_vector(to_unsigned(8,8) ,
59476	 => std_logic_vector(to_unsigned(9,8) ,
59477	 => std_logic_vector(to_unsigned(8,8) ,
59478	 => std_logic_vector(to_unsigned(4,8) ,
59479	 => std_logic_vector(to_unsigned(5,8) ,
59480	 => std_logic_vector(to_unsigned(8,8) ,
59481	 => std_logic_vector(to_unsigned(9,8) ,
59482	 => std_logic_vector(to_unsigned(11,8) ,
59483	 => std_logic_vector(to_unsigned(7,8) ,
59484	 => std_logic_vector(to_unsigned(0,8) ,
59485	 => std_logic_vector(to_unsigned(0,8) ,
59486	 => std_logic_vector(to_unsigned(0,8) ,
59487	 => std_logic_vector(to_unsigned(0,8) ,
59488	 => std_logic_vector(to_unsigned(0,8) ,
59489	 => std_logic_vector(to_unsigned(2,8) ,
59490	 => std_logic_vector(to_unsigned(4,8) ,
59491	 => std_logic_vector(to_unsigned(13,8) ,
59492	 => std_logic_vector(to_unsigned(20,8) ,
59493	 => std_logic_vector(to_unsigned(12,8) ,
59494	 => std_logic_vector(to_unsigned(8,8) ,
59495	 => std_logic_vector(to_unsigned(9,8) ,
59496	 => std_logic_vector(to_unsigned(14,8) ,
59497	 => std_logic_vector(to_unsigned(6,8) ,
59498	 => std_logic_vector(to_unsigned(6,8) ,
59499	 => std_logic_vector(to_unsigned(6,8) ,
59500	 => std_logic_vector(to_unsigned(7,8) ,
59501	 => std_logic_vector(to_unsigned(8,8) ,
59502	 => std_logic_vector(to_unsigned(7,8) ,
59503	 => std_logic_vector(to_unsigned(10,8) ,
59504	 => std_logic_vector(to_unsigned(30,8) ,
59505	 => std_logic_vector(to_unsigned(32,8) ,
59506	 => std_logic_vector(to_unsigned(33,8) ,
59507	 => std_logic_vector(to_unsigned(35,8) ,
59508	 => std_logic_vector(to_unsigned(19,8) ,
59509	 => std_logic_vector(to_unsigned(8,8) ,
59510	 => std_logic_vector(to_unsigned(4,8) ,
59511	 => std_logic_vector(to_unsigned(4,8) ,
59512	 => std_logic_vector(to_unsigned(5,8) ,
59513	 => std_logic_vector(to_unsigned(8,8) ,
59514	 => std_logic_vector(to_unsigned(10,8) ,
59515	 => std_logic_vector(to_unsigned(8,8) ,
59516	 => std_logic_vector(to_unsigned(11,8) ,
59517	 => std_logic_vector(to_unsigned(12,8) ,
59518	 => std_logic_vector(to_unsigned(12,8) ,
59519	 => std_logic_vector(to_unsigned(15,8) ,
59520	 => std_logic_vector(to_unsigned(14,8) ,
59521	 => std_logic_vector(to_unsigned(79,8) ,
59522	 => std_logic_vector(to_unsigned(88,8) ,
59523	 => std_logic_vector(to_unsigned(60,8) ,
59524	 => std_logic_vector(to_unsigned(68,8) ,
59525	 => std_logic_vector(to_unsigned(66,8) ,
59526	 => std_logic_vector(to_unsigned(44,8) ,
59527	 => std_logic_vector(to_unsigned(34,8) ,
59528	 => std_logic_vector(to_unsigned(45,8) ,
59529	 => std_logic_vector(to_unsigned(52,8) ,
59530	 => std_logic_vector(to_unsigned(46,8) ,
59531	 => std_logic_vector(to_unsigned(69,8) ,
59532	 => std_logic_vector(to_unsigned(56,8) ,
59533	 => std_logic_vector(to_unsigned(63,8) ,
59534	 => std_logic_vector(to_unsigned(90,8) ,
59535	 => std_logic_vector(to_unsigned(92,8) ,
59536	 => std_logic_vector(to_unsigned(69,8) ,
59537	 => std_logic_vector(to_unsigned(77,8) ,
59538	 => std_logic_vector(to_unsigned(61,8) ,
59539	 => std_logic_vector(to_unsigned(44,8) ,
59540	 => std_logic_vector(to_unsigned(51,8) ,
59541	 => std_logic_vector(to_unsigned(44,8) ,
59542	 => std_logic_vector(to_unsigned(37,8) ,
59543	 => std_logic_vector(to_unsigned(30,8) ,
59544	 => std_logic_vector(to_unsigned(25,8) ,
59545	 => std_logic_vector(to_unsigned(67,8) ,
59546	 => std_logic_vector(to_unsigned(77,8) ,
59547	 => std_logic_vector(to_unsigned(56,8) ,
59548	 => std_logic_vector(to_unsigned(48,8) ,
59549	 => std_logic_vector(to_unsigned(52,8) ,
59550	 => std_logic_vector(to_unsigned(55,8) ,
59551	 => std_logic_vector(to_unsigned(45,8) ,
59552	 => std_logic_vector(to_unsigned(40,8) ,
59553	 => std_logic_vector(to_unsigned(35,8) ,
59554	 => std_logic_vector(to_unsigned(32,8) ,
59555	 => std_logic_vector(to_unsigned(34,8) ,
59556	 => std_logic_vector(to_unsigned(48,8) ,
59557	 => std_logic_vector(to_unsigned(66,8) ,
59558	 => std_logic_vector(to_unsigned(46,8) ,
59559	 => std_logic_vector(to_unsigned(32,8) ,
59560	 => std_logic_vector(to_unsigned(54,8) ,
59561	 => std_logic_vector(to_unsigned(68,8) ,
59562	 => std_logic_vector(to_unsigned(84,8) ,
59563	 => std_logic_vector(to_unsigned(95,8) ,
59564	 => std_logic_vector(to_unsigned(66,8) ,
59565	 => std_logic_vector(to_unsigned(95,8) ,
59566	 => std_logic_vector(to_unsigned(93,8) ,
59567	 => std_logic_vector(to_unsigned(52,8) ,
59568	 => std_logic_vector(to_unsigned(62,8) ,
59569	 => std_logic_vector(to_unsigned(86,8) ,
59570	 => std_logic_vector(to_unsigned(64,8) ,
59571	 => std_logic_vector(to_unsigned(41,8) ,
59572	 => std_logic_vector(to_unsigned(52,8) ,
59573	 => std_logic_vector(to_unsigned(60,8) ,
59574	 => std_logic_vector(to_unsigned(45,8) ,
59575	 => std_logic_vector(to_unsigned(65,8) ,
59576	 => std_logic_vector(to_unsigned(84,8) ,
59577	 => std_logic_vector(to_unsigned(82,8) ,
59578	 => std_logic_vector(to_unsigned(42,8) ,
59579	 => std_logic_vector(to_unsigned(56,8) ,
59580	 => std_logic_vector(to_unsigned(69,8) ,
59581	 => std_logic_vector(to_unsigned(37,8) ,
59582	 => std_logic_vector(to_unsigned(31,8) ,
59583	 => std_logic_vector(to_unsigned(70,8) ,
59584	 => std_logic_vector(to_unsigned(69,8) ,
59585	 => std_logic_vector(to_unsigned(79,8) ,
59586	 => std_logic_vector(to_unsigned(87,8) ,
59587	 => std_logic_vector(to_unsigned(73,8) ,
59588	 => std_logic_vector(to_unsigned(107,8) ,
59589	 => std_logic_vector(to_unsigned(100,8) ,
59590	 => std_logic_vector(to_unsigned(93,8) ,
59591	 => std_logic_vector(to_unsigned(107,8) ,
59592	 => std_logic_vector(to_unsigned(90,8) ,
59593	 => std_logic_vector(to_unsigned(99,8) ,
59594	 => std_logic_vector(to_unsigned(133,8) ,
59595	 => std_logic_vector(to_unsigned(149,8) ,
59596	 => std_logic_vector(to_unsigned(134,8) ,
59597	 => std_logic_vector(to_unsigned(121,8) ,
59598	 => std_logic_vector(to_unsigned(130,8) ,
59599	 => std_logic_vector(to_unsigned(127,8) ,
59600	 => std_logic_vector(to_unsigned(116,8) ,
59601	 => std_logic_vector(to_unsigned(122,8) ,
59602	 => std_logic_vector(to_unsigned(121,8) ,
59603	 => std_logic_vector(to_unsigned(115,8) ,
59604	 => std_logic_vector(to_unsigned(105,8) ,
59605	 => std_logic_vector(to_unsigned(128,8) ,
59606	 => std_logic_vector(to_unsigned(95,8) ,
59607	 => std_logic_vector(to_unsigned(35,8) ,
59608	 => std_logic_vector(to_unsigned(42,8) ,
59609	 => std_logic_vector(to_unsigned(45,8) ,
59610	 => std_logic_vector(to_unsigned(44,8) ,
59611	 => std_logic_vector(to_unsigned(41,8) ,
59612	 => std_logic_vector(to_unsigned(38,8) ,
59613	 => std_logic_vector(to_unsigned(49,8) ,
59614	 => std_logic_vector(to_unsigned(51,8) ,
59615	 => std_logic_vector(to_unsigned(53,8) ,
59616	 => std_logic_vector(to_unsigned(47,8) ,
59617	 => std_logic_vector(to_unsigned(66,8) ,
59618	 => std_logic_vector(to_unsigned(60,8) ,
59619	 => std_logic_vector(to_unsigned(51,8) ,
59620	 => std_logic_vector(to_unsigned(59,8) ,
59621	 => std_logic_vector(to_unsigned(68,8) ,
59622	 => std_logic_vector(to_unsigned(76,8) ,
59623	 => std_logic_vector(to_unsigned(68,8) ,
59624	 => std_logic_vector(to_unsigned(58,8) ,
59625	 => std_logic_vector(to_unsigned(66,8) ,
59626	 => std_logic_vector(to_unsigned(85,8) ,
59627	 => std_logic_vector(to_unsigned(96,8) ,
59628	 => std_logic_vector(to_unsigned(63,8) ,
59629	 => std_logic_vector(to_unsigned(43,8) ,
59630	 => std_logic_vector(to_unsigned(44,8) ,
59631	 => std_logic_vector(to_unsigned(49,8) ,
59632	 => std_logic_vector(to_unsigned(54,8) ,
59633	 => std_logic_vector(to_unsigned(64,8) ,
59634	 => std_logic_vector(to_unsigned(43,8) ,
59635	 => std_logic_vector(to_unsigned(41,8) ,
59636	 => std_logic_vector(to_unsigned(57,8) ,
59637	 => std_logic_vector(to_unsigned(50,8) ,
59638	 => std_logic_vector(to_unsigned(39,8) ,
59639	 => std_logic_vector(to_unsigned(20,8) ,
59640	 => std_logic_vector(to_unsigned(12,8) ,
59641	 => std_logic_vector(to_unsigned(37,8) ,
59642	 => std_logic_vector(to_unsigned(25,8) ,
59643	 => std_logic_vector(to_unsigned(45,8) ,
59644	 => std_logic_vector(to_unsigned(29,8) ,
59645	 => std_logic_vector(to_unsigned(27,8) ,
59646	 => std_logic_vector(to_unsigned(34,8) ,
59647	 => std_logic_vector(to_unsigned(54,8) ,
59648	 => std_logic_vector(to_unsigned(68,8) ,
59649	 => std_logic_vector(to_unsigned(67,8) ,
59650	 => std_logic_vector(to_unsigned(43,8) ,
59651	 => std_logic_vector(to_unsigned(17,8) ,
59652	 => std_logic_vector(to_unsigned(18,8) ,
59653	 => std_logic_vector(to_unsigned(17,8) ,
59654	 => std_logic_vector(to_unsigned(27,8) ,
59655	 => std_logic_vector(to_unsigned(30,8) ,
59656	 => std_logic_vector(to_unsigned(16,8) ,
59657	 => std_logic_vector(to_unsigned(16,8) ,
59658	 => std_logic_vector(to_unsigned(13,8) ,
59659	 => std_logic_vector(to_unsigned(12,8) ,
59660	 => std_logic_vector(to_unsigned(16,8) ,
59661	 => std_logic_vector(to_unsigned(20,8) ,
59662	 => std_logic_vector(to_unsigned(17,8) ,
59663	 => std_logic_vector(to_unsigned(17,8) ,
59664	 => std_logic_vector(to_unsigned(33,8) ,
59665	 => std_logic_vector(to_unsigned(45,8) ,
59666	 => std_logic_vector(to_unsigned(32,8) ,
59667	 => std_logic_vector(to_unsigned(30,8) ,
59668	 => std_logic_vector(to_unsigned(29,8) ,
59669	 => std_logic_vector(to_unsigned(23,8) ,
59670	 => std_logic_vector(to_unsigned(50,8) ,
59671	 => std_logic_vector(to_unsigned(23,8) ,
59672	 => std_logic_vector(to_unsigned(21,8) ,
59673	 => std_logic_vector(to_unsigned(32,8) ,
59674	 => std_logic_vector(to_unsigned(25,8) ,
59675	 => std_logic_vector(to_unsigned(31,8) ,
59676	 => std_logic_vector(to_unsigned(29,8) ,
59677	 => std_logic_vector(to_unsigned(25,8) ,
59678	 => std_logic_vector(to_unsigned(29,8) ,
59679	 => std_logic_vector(to_unsigned(23,8) ,
59680	 => std_logic_vector(to_unsigned(33,8) ,
59681	 => std_logic_vector(to_unsigned(122,8) ,
59682	 => std_logic_vector(to_unsigned(122,8) ,
59683	 => std_logic_vector(to_unsigned(99,8) ,
59684	 => std_logic_vector(to_unsigned(92,8) ,
59685	 => std_logic_vector(to_unsigned(100,8) ,
59686	 => std_logic_vector(to_unsigned(91,8) ,
59687	 => std_logic_vector(to_unsigned(95,8) ,
59688	 => std_logic_vector(to_unsigned(28,8) ,
59689	 => std_logic_vector(to_unsigned(34,8) ,
59690	 => std_logic_vector(to_unsigned(62,8) ,
59691	 => std_logic_vector(to_unsigned(27,8) ,
59692	 => std_logic_vector(to_unsigned(32,8) ,
59693	 => std_logic_vector(to_unsigned(44,8) ,
59694	 => std_logic_vector(to_unsigned(42,8) ,
59695	 => std_logic_vector(to_unsigned(41,8) ,
59696	 => std_logic_vector(to_unsigned(63,8) ,
59697	 => std_logic_vector(to_unsigned(34,8) ,
59698	 => std_logic_vector(to_unsigned(12,8) ,
59699	 => std_logic_vector(to_unsigned(7,8) ,
59700	 => std_logic_vector(to_unsigned(10,8) ,
59701	 => std_logic_vector(to_unsigned(8,8) ,
59702	 => std_logic_vector(to_unsigned(8,8) ,
59703	 => std_logic_vector(to_unsigned(9,8) ,
59704	 => std_logic_vector(to_unsigned(11,8) ,
59705	 => std_logic_vector(to_unsigned(9,8) ,
59706	 => std_logic_vector(to_unsigned(10,8) ,
59707	 => std_logic_vector(to_unsigned(17,8) ,
59708	 => std_logic_vector(to_unsigned(30,8) ,
59709	 => std_logic_vector(to_unsigned(26,8) ,
59710	 => std_logic_vector(to_unsigned(29,8) ,
59711	 => std_logic_vector(to_unsigned(39,8) ,
59712	 => std_logic_vector(to_unsigned(38,8) ,
59713	 => std_logic_vector(to_unsigned(33,8) ,
59714	 => std_logic_vector(to_unsigned(31,8) ,
59715	 => std_logic_vector(to_unsigned(45,8) ,
59716	 => std_logic_vector(to_unsigned(40,8) ,
59717	 => std_logic_vector(to_unsigned(33,8) ,
59718	 => std_logic_vector(to_unsigned(48,8) ,
59719	 => std_logic_vector(to_unsigned(46,8) ,
59720	 => std_logic_vector(to_unsigned(25,8) ,
59721	 => std_logic_vector(to_unsigned(30,8) ,
59722	 => std_logic_vector(to_unsigned(48,8) ,
59723	 => std_logic_vector(to_unsigned(37,8) ,
59724	 => std_logic_vector(to_unsigned(24,8) ,
59725	 => std_logic_vector(to_unsigned(30,8) ,
59726	 => std_logic_vector(to_unsigned(48,8) ,
59727	 => std_logic_vector(to_unsigned(65,8) ,
59728	 => std_logic_vector(to_unsigned(59,8) ,
59729	 => std_logic_vector(to_unsigned(21,8) ,
59730	 => std_logic_vector(to_unsigned(12,8) ,
59731	 => std_logic_vector(to_unsigned(25,8) ,
59732	 => std_logic_vector(to_unsigned(20,8) ,
59733	 => std_logic_vector(to_unsigned(16,8) ,
59734	 => std_logic_vector(to_unsigned(24,8) ,
59735	 => std_logic_vector(to_unsigned(29,8) ,
59736	 => std_logic_vector(to_unsigned(21,8) ,
59737	 => std_logic_vector(to_unsigned(16,8) ,
59738	 => std_logic_vector(to_unsigned(21,8) ,
59739	 => std_logic_vector(to_unsigned(26,8) ,
59740	 => std_logic_vector(to_unsigned(23,8) ,
59741	 => std_logic_vector(to_unsigned(32,8) ,
59742	 => std_logic_vector(to_unsigned(30,8) ,
59743	 => std_logic_vector(to_unsigned(25,8) ,
59744	 => std_logic_vector(to_unsigned(32,8) ,
59745	 => std_logic_vector(to_unsigned(41,8) ,
59746	 => std_logic_vector(to_unsigned(20,8) ,
59747	 => std_logic_vector(to_unsigned(16,8) ,
59748	 => std_logic_vector(to_unsigned(14,8) ,
59749	 => std_logic_vector(to_unsigned(38,8) ,
59750	 => std_logic_vector(to_unsigned(62,8) ,
59751	 => std_logic_vector(to_unsigned(45,8) ,
59752	 => std_logic_vector(to_unsigned(27,8) ,
59753	 => std_logic_vector(to_unsigned(11,8) ,
59754	 => std_logic_vector(to_unsigned(25,8) ,
59755	 => std_logic_vector(to_unsigned(70,8) ,
59756	 => std_logic_vector(to_unsigned(95,8) ,
59757	 => std_logic_vector(to_unsigned(80,8) ,
59758	 => std_logic_vector(to_unsigned(41,8) ,
59759	 => std_logic_vector(to_unsigned(30,8) ,
59760	 => std_logic_vector(to_unsigned(33,8) ,
59761	 => std_logic_vector(to_unsigned(38,8) ,
59762	 => std_logic_vector(to_unsigned(50,8) ,
59763	 => std_logic_vector(to_unsigned(52,8) ,
59764	 => std_logic_vector(to_unsigned(65,8) ,
59765	 => std_logic_vector(to_unsigned(104,8) ,
59766	 => std_logic_vector(to_unsigned(105,8) ,
59767	 => std_logic_vector(to_unsigned(90,8) ,
59768	 => std_logic_vector(to_unsigned(108,8) ,
59769	 => std_logic_vector(to_unsigned(76,8) ,
59770	 => std_logic_vector(to_unsigned(41,8) ,
59771	 => std_logic_vector(to_unsigned(17,8) ,
59772	 => std_logic_vector(to_unsigned(19,8) ,
59773	 => std_logic_vector(to_unsigned(14,8) ,
59774	 => std_logic_vector(to_unsigned(12,8) ,
59775	 => std_logic_vector(to_unsigned(13,8) ,
59776	 => std_logic_vector(to_unsigned(10,8) ,
59777	 => std_logic_vector(to_unsigned(12,8) ,
59778	 => std_logic_vector(to_unsigned(11,8) ,
59779	 => std_logic_vector(to_unsigned(11,8) ,
59780	 => std_logic_vector(to_unsigned(9,8) ,
59781	 => std_logic_vector(to_unsigned(23,8) ,
59782	 => std_logic_vector(to_unsigned(25,8) ,
59783	 => std_logic_vector(to_unsigned(17,8) ,
59784	 => std_logic_vector(to_unsigned(10,8) ,
59785	 => std_logic_vector(to_unsigned(1,8) ,
59786	 => std_logic_vector(to_unsigned(1,8) ,
59787	 => std_logic_vector(to_unsigned(17,8) ,
59788	 => std_logic_vector(to_unsigned(54,8) ,
59789	 => std_logic_vector(to_unsigned(25,8) ,
59790	 => std_logic_vector(to_unsigned(6,8) ,
59791	 => std_logic_vector(to_unsigned(8,8) ,
59792	 => std_logic_vector(to_unsigned(24,8) ,
59793	 => std_logic_vector(to_unsigned(18,8) ,
59794	 => std_logic_vector(to_unsigned(11,8) ,
59795	 => std_logic_vector(to_unsigned(8,8) ,
59796	 => std_logic_vector(to_unsigned(8,8) ,
59797	 => std_logic_vector(to_unsigned(6,8) ,
59798	 => std_logic_vector(to_unsigned(3,8) ,
59799	 => std_logic_vector(to_unsigned(11,8) ,
59800	 => std_logic_vector(to_unsigned(13,8) ,
59801	 => std_logic_vector(to_unsigned(10,8) ,
59802	 => std_logic_vector(to_unsigned(15,8) ,
59803	 => std_logic_vector(to_unsigned(14,8) ,
59804	 => std_logic_vector(to_unsigned(1,8) ,
59805	 => std_logic_vector(to_unsigned(0,8) ,
59806	 => std_logic_vector(to_unsigned(0,8) ,
59807	 => std_logic_vector(to_unsigned(0,8) ,
59808	 => std_logic_vector(to_unsigned(0,8) ,
59809	 => std_logic_vector(to_unsigned(10,8) ,
59810	 => std_logic_vector(to_unsigned(30,8) ,
59811	 => std_logic_vector(to_unsigned(27,8) ,
59812	 => std_logic_vector(to_unsigned(22,8) ,
59813	 => std_logic_vector(to_unsigned(14,8) ,
59814	 => std_logic_vector(to_unsigned(17,8) ,
59815	 => std_logic_vector(to_unsigned(18,8) ,
59816	 => std_logic_vector(to_unsigned(16,8) ,
59817	 => std_logic_vector(to_unsigned(8,8) ,
59818	 => std_logic_vector(to_unsigned(7,8) ,
59819	 => std_logic_vector(to_unsigned(7,8) ,
59820	 => std_logic_vector(to_unsigned(5,8) ,
59821	 => std_logic_vector(to_unsigned(8,8) ,
59822	 => std_logic_vector(to_unsigned(8,8) ,
59823	 => std_logic_vector(to_unsigned(7,8) ,
59824	 => std_logic_vector(to_unsigned(39,8) ,
59825	 => std_logic_vector(to_unsigned(43,8) ,
59826	 => std_logic_vector(to_unsigned(23,8) ,
59827	 => std_logic_vector(to_unsigned(34,8) ,
59828	 => std_logic_vector(to_unsigned(23,8) ,
59829	 => std_logic_vector(to_unsigned(10,8) ,
59830	 => std_logic_vector(to_unsigned(6,8) ,
59831	 => std_logic_vector(to_unsigned(6,8) ,
59832	 => std_logic_vector(to_unsigned(6,8) ,
59833	 => std_logic_vector(to_unsigned(8,8) ,
59834	 => std_logic_vector(to_unsigned(9,8) ,
59835	 => std_logic_vector(to_unsigned(10,8) ,
59836	 => std_logic_vector(to_unsigned(13,8) ,
59837	 => std_logic_vector(to_unsigned(17,8) ,
59838	 => std_logic_vector(to_unsigned(15,8) ,
59839	 => std_logic_vector(to_unsigned(16,8) ,
59840	 => std_logic_vector(to_unsigned(19,8) ,
59841	 => std_logic_vector(to_unsigned(78,8) ,
59842	 => std_logic_vector(to_unsigned(97,8) ,
59843	 => std_logic_vector(to_unsigned(70,8) ,
59844	 => std_logic_vector(to_unsigned(69,8) ,
59845	 => std_logic_vector(to_unsigned(62,8) ,
59846	 => std_logic_vector(to_unsigned(41,8) ,
59847	 => std_logic_vector(to_unsigned(35,8) ,
59848	 => std_logic_vector(to_unsigned(47,8) ,
59849	 => std_logic_vector(to_unsigned(51,8) ,
59850	 => std_logic_vector(to_unsigned(43,8) ,
59851	 => std_logic_vector(to_unsigned(62,8) ,
59852	 => std_logic_vector(to_unsigned(52,8) ,
59853	 => std_logic_vector(to_unsigned(55,8) ,
59854	 => std_logic_vector(to_unsigned(85,8) ,
59855	 => std_logic_vector(to_unsigned(88,8) ,
59856	 => std_logic_vector(to_unsigned(54,8) ,
59857	 => std_logic_vector(to_unsigned(59,8) ,
59858	 => std_logic_vector(to_unsigned(72,8) ,
59859	 => std_logic_vector(to_unsigned(58,8) ,
59860	 => std_logic_vector(to_unsigned(62,8) ,
59861	 => std_logic_vector(to_unsigned(52,8) ,
59862	 => std_logic_vector(to_unsigned(41,8) ,
59863	 => std_logic_vector(to_unsigned(34,8) ,
59864	 => std_logic_vector(to_unsigned(36,8) ,
59865	 => std_logic_vector(to_unsigned(68,8) ,
59866	 => std_logic_vector(to_unsigned(69,8) ,
59867	 => std_logic_vector(to_unsigned(54,8) ,
59868	 => std_logic_vector(to_unsigned(41,8) ,
59869	 => std_logic_vector(to_unsigned(39,8) ,
59870	 => std_logic_vector(to_unsigned(46,8) ,
59871	 => std_logic_vector(to_unsigned(41,8) ,
59872	 => std_logic_vector(to_unsigned(35,8) ,
59873	 => std_logic_vector(to_unsigned(45,8) ,
59874	 => std_logic_vector(to_unsigned(57,8) ,
59875	 => std_logic_vector(to_unsigned(52,8) ,
59876	 => std_logic_vector(to_unsigned(56,8) ,
59877	 => std_logic_vector(to_unsigned(60,8) ,
59878	 => std_logic_vector(to_unsigned(51,8) ,
59879	 => std_logic_vector(to_unsigned(53,8) ,
59880	 => std_logic_vector(to_unsigned(51,8) ,
59881	 => std_logic_vector(to_unsigned(62,8) ,
59882	 => std_logic_vector(to_unsigned(69,8) ,
59883	 => std_logic_vector(to_unsigned(65,8) ,
59884	 => std_logic_vector(to_unsigned(68,8) ,
59885	 => std_logic_vector(to_unsigned(74,8) ,
59886	 => std_logic_vector(to_unsigned(88,8) ,
59887	 => std_logic_vector(to_unsigned(66,8) ,
59888	 => std_logic_vector(to_unsigned(71,8) ,
59889	 => std_logic_vector(to_unsigned(86,8) ,
59890	 => std_logic_vector(to_unsigned(67,8) ,
59891	 => std_logic_vector(to_unsigned(45,8) ,
59892	 => std_logic_vector(to_unsigned(42,8) ,
59893	 => std_logic_vector(to_unsigned(56,8) ,
59894	 => std_logic_vector(to_unsigned(44,8) ,
59895	 => std_logic_vector(to_unsigned(51,8) ,
59896	 => std_logic_vector(to_unsigned(76,8) ,
59897	 => std_logic_vector(to_unsigned(72,8) ,
59898	 => std_logic_vector(to_unsigned(41,8) ,
59899	 => std_logic_vector(to_unsigned(47,8) ,
59900	 => std_logic_vector(to_unsigned(51,8) ,
59901	 => std_logic_vector(to_unsigned(45,8) ,
59902	 => std_logic_vector(to_unsigned(51,8) ,
59903	 => std_logic_vector(to_unsigned(73,8) ,
59904	 => std_logic_vector(to_unsigned(85,8) ,
59905	 => std_logic_vector(to_unsigned(87,8) ,
59906	 => std_logic_vector(to_unsigned(87,8) ,
59907	 => std_logic_vector(to_unsigned(80,8) ,
59908	 => std_logic_vector(to_unsigned(91,8) ,
59909	 => std_logic_vector(to_unsigned(84,8) ,
59910	 => std_logic_vector(to_unsigned(82,8) ,
59911	 => std_logic_vector(to_unsigned(115,8) ,
59912	 => std_logic_vector(to_unsigned(82,8) ,
59913	 => std_logic_vector(to_unsigned(90,8) ,
59914	 => std_logic_vector(to_unsigned(141,8) ,
59915	 => std_logic_vector(to_unsigned(138,8) ,
59916	 => std_logic_vector(to_unsigned(138,8) ,
59917	 => std_logic_vector(to_unsigned(130,8) ,
59918	 => std_logic_vector(to_unsigned(121,8) ,
59919	 => std_logic_vector(to_unsigned(121,8) ,
59920	 => std_logic_vector(to_unsigned(128,8) ,
59921	 => std_logic_vector(to_unsigned(127,8) ,
59922	 => std_logic_vector(to_unsigned(109,8) ,
59923	 => std_logic_vector(to_unsigned(119,8) ,
59924	 => std_logic_vector(to_unsigned(122,8) ,
59925	 => std_logic_vector(to_unsigned(122,8) ,
59926	 => std_logic_vector(to_unsigned(105,8) ,
59927	 => std_logic_vector(to_unsigned(43,8) ,
59928	 => std_logic_vector(to_unsigned(32,8) ,
59929	 => std_logic_vector(to_unsigned(37,8) ,
59930	 => std_logic_vector(to_unsigned(39,8) ,
59931	 => std_logic_vector(to_unsigned(42,8) ,
59932	 => std_logic_vector(to_unsigned(42,8) ,
59933	 => std_logic_vector(to_unsigned(43,8) ,
59934	 => std_logic_vector(to_unsigned(50,8) ,
59935	 => std_logic_vector(to_unsigned(64,8) ,
59936	 => std_logic_vector(to_unsigned(57,8) ,
59937	 => std_logic_vector(to_unsigned(52,8) ,
59938	 => std_logic_vector(to_unsigned(56,8) ,
59939	 => std_logic_vector(to_unsigned(58,8) ,
59940	 => std_logic_vector(to_unsigned(63,8) ,
59941	 => std_logic_vector(to_unsigned(64,8) ,
59942	 => std_logic_vector(to_unsigned(57,8) ,
59943	 => std_logic_vector(to_unsigned(57,8) ,
59944	 => std_logic_vector(to_unsigned(60,8) ,
59945	 => std_logic_vector(to_unsigned(70,8) ,
59946	 => std_logic_vector(to_unsigned(79,8) ,
59947	 => std_logic_vector(to_unsigned(85,8) ,
59948	 => std_logic_vector(to_unsigned(58,8) ,
59949	 => std_logic_vector(to_unsigned(37,8) ,
59950	 => std_logic_vector(to_unsigned(40,8) ,
59951	 => std_logic_vector(to_unsigned(45,8) ,
59952	 => std_logic_vector(to_unsigned(50,8) ,
59953	 => std_logic_vector(to_unsigned(64,8) ,
59954	 => std_logic_vector(to_unsigned(44,8) ,
59955	 => std_logic_vector(to_unsigned(40,8) ,
59956	 => std_logic_vector(to_unsigned(55,8) ,
59957	 => std_logic_vector(to_unsigned(42,8) ,
59958	 => std_logic_vector(to_unsigned(33,8) ,
59959	 => std_logic_vector(to_unsigned(30,8) ,
59960	 => std_logic_vector(to_unsigned(38,8) ,
59961	 => std_logic_vector(to_unsigned(57,8) ,
59962	 => std_logic_vector(to_unsigned(41,8) ,
59963	 => std_logic_vector(to_unsigned(54,8) ,
59964	 => std_logic_vector(to_unsigned(25,8) ,
59965	 => std_logic_vector(to_unsigned(11,8) ,
59966	 => std_logic_vector(to_unsigned(11,8) ,
59967	 => std_logic_vector(to_unsigned(16,8) ,
59968	 => std_logic_vector(to_unsigned(25,8) ,
59969	 => std_logic_vector(to_unsigned(35,8) ,
59970	 => std_logic_vector(to_unsigned(50,8) ,
59971	 => std_logic_vector(to_unsigned(20,8) ,
59972	 => std_logic_vector(to_unsigned(24,8) ,
59973	 => std_logic_vector(to_unsigned(34,8) ,
59974	 => std_logic_vector(to_unsigned(54,8) ,
59975	 => std_logic_vector(to_unsigned(31,8) ,
59976	 => std_logic_vector(to_unsigned(16,8) ,
59977	 => std_logic_vector(to_unsigned(13,8) ,
59978	 => std_logic_vector(to_unsigned(11,8) ,
59979	 => std_logic_vector(to_unsigned(19,8) ,
59980	 => std_logic_vector(to_unsigned(17,8) ,
59981	 => std_logic_vector(to_unsigned(14,8) ,
59982	 => std_logic_vector(to_unsigned(13,8) ,
59983	 => std_logic_vector(to_unsigned(13,8) ,
59984	 => std_logic_vector(to_unsigned(53,8) ,
59985	 => std_logic_vector(to_unsigned(73,8) ,
59986	 => std_logic_vector(to_unsigned(49,8) ,
59987	 => std_logic_vector(to_unsigned(44,8) ,
59988	 => std_logic_vector(to_unsigned(38,8) ,
59989	 => std_logic_vector(to_unsigned(34,8) ,
59990	 => std_logic_vector(to_unsigned(27,8) ,
59991	 => std_logic_vector(to_unsigned(19,8) ,
59992	 => std_logic_vector(to_unsigned(23,8) ,
59993	 => std_logic_vector(to_unsigned(40,8) ,
59994	 => std_logic_vector(to_unsigned(31,8) ,
59995	 => std_logic_vector(to_unsigned(30,8) ,
59996	 => std_logic_vector(to_unsigned(33,8) ,
59997	 => std_logic_vector(to_unsigned(29,8) ,
59998	 => std_logic_vector(to_unsigned(29,8) ,
59999	 => std_logic_vector(to_unsigned(54,8) ,
60000	 => std_logic_vector(to_unsigned(88,8) ,
60001	 => std_logic_vector(to_unsigned(118,8) ,
60002	 => std_logic_vector(to_unsigned(144,8) ,
60003	 => std_logic_vector(to_unsigned(128,8) ,
60004	 => std_logic_vector(to_unsigned(30,8) ,
60005	 => std_logic_vector(to_unsigned(12,8) ,
60006	 => std_logic_vector(to_unsigned(17,8) ,
60007	 => std_logic_vector(to_unsigned(14,8) ,
60008	 => std_logic_vector(to_unsigned(17,8) ,
60009	 => std_logic_vector(to_unsigned(29,8) ,
60010	 => std_logic_vector(to_unsigned(35,8) ,
60011	 => std_logic_vector(to_unsigned(37,8) ,
60012	 => std_logic_vector(to_unsigned(46,8) ,
60013	 => std_logic_vector(to_unsigned(42,8) ,
60014	 => std_logic_vector(to_unsigned(37,8) ,
60015	 => std_logic_vector(to_unsigned(62,8) ,
60016	 => std_logic_vector(to_unsigned(95,8) ,
60017	 => std_logic_vector(to_unsigned(34,8) ,
60018	 => std_logic_vector(to_unsigned(17,8) ,
60019	 => std_logic_vector(to_unsigned(39,8) ,
60020	 => std_logic_vector(to_unsigned(52,8) ,
60021	 => std_logic_vector(to_unsigned(20,8) ,
60022	 => std_logic_vector(to_unsigned(9,8) ,
60023	 => std_logic_vector(to_unsigned(10,8) ,
60024	 => std_logic_vector(to_unsigned(16,8) ,
60025	 => std_logic_vector(to_unsigned(19,8) ,
60026	 => std_logic_vector(to_unsigned(14,8) ,
60027	 => std_logic_vector(to_unsigned(30,8) ,
60028	 => std_logic_vector(to_unsigned(29,8) ,
60029	 => std_logic_vector(to_unsigned(19,8) ,
60030	 => std_logic_vector(to_unsigned(38,8) ,
60031	 => std_logic_vector(to_unsigned(39,8) ,
60032	 => std_logic_vector(to_unsigned(36,8) ,
60033	 => std_logic_vector(to_unsigned(42,8) ,
60034	 => std_logic_vector(to_unsigned(47,8) ,
60035	 => std_logic_vector(to_unsigned(43,8) ,
60036	 => std_logic_vector(to_unsigned(36,8) ,
60037	 => std_logic_vector(to_unsigned(38,8) ,
60038	 => std_logic_vector(to_unsigned(51,8) ,
60039	 => std_logic_vector(to_unsigned(49,8) ,
60040	 => std_logic_vector(to_unsigned(29,8) ,
60041	 => std_logic_vector(to_unsigned(32,8) ,
60042	 => std_logic_vector(to_unsigned(48,8) ,
60043	 => std_logic_vector(to_unsigned(32,8) ,
60044	 => std_logic_vector(to_unsigned(25,8) ,
60045	 => std_logic_vector(to_unsigned(31,8) ,
60046	 => std_logic_vector(to_unsigned(33,8) ,
60047	 => std_logic_vector(to_unsigned(42,8) ,
60048	 => std_logic_vector(to_unsigned(37,8) ,
60049	 => std_logic_vector(to_unsigned(23,8) ,
60050	 => std_logic_vector(to_unsigned(18,8) ,
60051	 => std_logic_vector(to_unsigned(20,8) ,
60052	 => std_logic_vector(to_unsigned(13,8) ,
60053	 => std_logic_vector(to_unsigned(12,8) ,
60054	 => std_logic_vector(to_unsigned(18,8) ,
60055	 => std_logic_vector(to_unsigned(21,8) ,
60056	 => std_logic_vector(to_unsigned(22,8) ,
60057	 => std_logic_vector(to_unsigned(14,8) ,
60058	 => std_logic_vector(to_unsigned(14,8) ,
60059	 => std_logic_vector(to_unsigned(23,8) ,
60060	 => std_logic_vector(to_unsigned(23,8) ,
60061	 => std_logic_vector(to_unsigned(29,8) ,
60062	 => std_logic_vector(to_unsigned(37,8) ,
60063	 => std_logic_vector(to_unsigned(30,8) ,
60064	 => std_logic_vector(to_unsigned(49,8) ,
60065	 => std_logic_vector(to_unsigned(29,8) ,
60066	 => std_logic_vector(to_unsigned(6,8) ,
60067	 => std_logic_vector(to_unsigned(11,8) ,
60068	 => std_logic_vector(to_unsigned(31,8) ,
60069	 => std_logic_vector(to_unsigned(73,8) ,
60070	 => std_logic_vector(to_unsigned(61,8) ,
60071	 => std_logic_vector(to_unsigned(37,8) ,
60072	 => std_logic_vector(to_unsigned(17,8) ,
60073	 => std_logic_vector(to_unsigned(26,8) ,
60074	 => std_logic_vector(to_unsigned(25,8) ,
60075	 => std_logic_vector(to_unsigned(28,8) ,
60076	 => std_logic_vector(to_unsigned(42,8) ,
60077	 => std_logic_vector(to_unsigned(58,8) ,
60078	 => std_logic_vector(to_unsigned(43,8) ,
60079	 => std_logic_vector(to_unsigned(41,8) ,
60080	 => std_logic_vector(to_unsigned(85,8) ,
60081	 => std_logic_vector(to_unsigned(108,8) ,
60082	 => std_logic_vector(to_unsigned(109,8) ,
60083	 => std_logic_vector(to_unsigned(121,8) ,
60084	 => std_logic_vector(to_unsigned(130,8) ,
60085	 => std_logic_vector(to_unsigned(85,8) ,
60086	 => std_logic_vector(to_unsigned(79,8) ,
60087	 => std_logic_vector(to_unsigned(38,8) ,
60088	 => std_logic_vector(to_unsigned(20,8) ,
60089	 => std_logic_vector(to_unsigned(18,8) ,
60090	 => std_logic_vector(to_unsigned(18,8) ,
60091	 => std_logic_vector(to_unsigned(20,8) ,
60092	 => std_logic_vector(to_unsigned(28,8) ,
60093	 => std_logic_vector(to_unsigned(27,8) ,
60094	 => std_logic_vector(to_unsigned(19,8) ,
60095	 => std_logic_vector(to_unsigned(23,8) ,
60096	 => std_logic_vector(to_unsigned(14,8) ,
60097	 => std_logic_vector(to_unsigned(10,8) ,
60098	 => std_logic_vector(to_unsigned(13,8) ,
60099	 => std_logic_vector(to_unsigned(15,8) ,
60100	 => std_logic_vector(to_unsigned(13,8) ,
60101	 => std_logic_vector(to_unsigned(20,8) ,
60102	 => std_logic_vector(to_unsigned(19,8) ,
60103	 => std_logic_vector(to_unsigned(17,8) ,
60104	 => std_logic_vector(to_unsigned(16,8) ,
60105	 => std_logic_vector(to_unsigned(2,8) ,
60106	 => std_logic_vector(to_unsigned(0,8) ,
60107	 => std_logic_vector(to_unsigned(5,8) ,
60108	 => std_logic_vector(to_unsigned(28,8) ,
60109	 => std_logic_vector(to_unsigned(16,8) ,
60110	 => std_logic_vector(to_unsigned(11,8) ,
60111	 => std_logic_vector(to_unsigned(13,8) ,
60112	 => std_logic_vector(to_unsigned(24,8) ,
60113	 => std_logic_vector(to_unsigned(27,8) ,
60114	 => std_logic_vector(to_unsigned(19,8) ,
60115	 => std_logic_vector(to_unsigned(13,8) ,
60116	 => std_logic_vector(to_unsigned(11,8) ,
60117	 => std_logic_vector(to_unsigned(6,8) ,
60118	 => std_logic_vector(to_unsigned(8,8) ,
60119	 => std_logic_vector(to_unsigned(15,8) ,
60120	 => std_logic_vector(to_unsigned(10,8) ,
60121	 => std_logic_vector(to_unsigned(13,8) ,
60122	 => std_logic_vector(to_unsigned(16,8) ,
60123	 => std_logic_vector(to_unsigned(12,8) ,
60124	 => std_logic_vector(to_unsigned(1,8) ,
60125	 => std_logic_vector(to_unsigned(0,8) ,
60126	 => std_logic_vector(to_unsigned(1,8) ,
60127	 => std_logic_vector(to_unsigned(1,8) ,
60128	 => std_logic_vector(to_unsigned(0,8) ,
60129	 => std_logic_vector(to_unsigned(2,8) ,
60130	 => std_logic_vector(to_unsigned(17,8) ,
60131	 => std_logic_vector(to_unsigned(13,8) ,
60132	 => std_logic_vector(to_unsigned(13,8) ,
60133	 => std_logic_vector(to_unsigned(25,8) ,
60134	 => std_logic_vector(to_unsigned(29,8) ,
60135	 => std_logic_vector(to_unsigned(23,8) ,
60136	 => std_logic_vector(to_unsigned(11,8) ,
60137	 => std_logic_vector(to_unsigned(5,8) ,
60138	 => std_logic_vector(to_unsigned(12,8) ,
60139	 => std_logic_vector(to_unsigned(23,8) ,
60140	 => std_logic_vector(to_unsigned(20,8) ,
60141	 => std_logic_vector(to_unsigned(11,8) ,
60142	 => std_logic_vector(to_unsigned(9,8) ,
60143	 => std_logic_vector(to_unsigned(8,8) ,
60144	 => std_logic_vector(to_unsigned(15,8) ,
60145	 => std_logic_vector(to_unsigned(16,8) ,
60146	 => std_logic_vector(to_unsigned(6,8) ,
60147	 => std_logic_vector(to_unsigned(13,8) ,
60148	 => std_logic_vector(to_unsigned(11,8) ,
60149	 => std_logic_vector(to_unsigned(7,8) ,
60150	 => std_logic_vector(to_unsigned(5,8) ,
60151	 => std_logic_vector(to_unsigned(6,8) ,
60152	 => std_logic_vector(to_unsigned(7,8) ,
60153	 => std_logic_vector(to_unsigned(9,8) ,
60154	 => std_logic_vector(to_unsigned(8,8) ,
60155	 => std_logic_vector(to_unsigned(9,8) ,
60156	 => std_logic_vector(to_unsigned(12,8) ,
60157	 => std_logic_vector(to_unsigned(14,8) ,
60158	 => std_logic_vector(to_unsigned(15,8) ,
60159	 => std_logic_vector(to_unsigned(17,8) ,
60160	 => std_logic_vector(to_unsigned(24,8) ,
60161	 => std_logic_vector(to_unsigned(73,8) ,
60162	 => std_logic_vector(to_unsigned(95,8) ,
60163	 => std_logic_vector(to_unsigned(79,8) ,
60164	 => std_logic_vector(to_unsigned(71,8) ,
60165	 => std_logic_vector(to_unsigned(68,8) ,
60166	 => std_logic_vector(to_unsigned(45,8) ,
60167	 => std_logic_vector(to_unsigned(33,8) ,
60168	 => std_logic_vector(to_unsigned(38,8) ,
60169	 => std_logic_vector(to_unsigned(55,8) ,
60170	 => std_logic_vector(to_unsigned(51,8) ,
60171	 => std_logic_vector(to_unsigned(59,8) ,
60172	 => std_logic_vector(to_unsigned(54,8) ,
60173	 => std_logic_vector(to_unsigned(49,8) ,
60174	 => std_logic_vector(to_unsigned(76,8) ,
60175	 => std_logic_vector(to_unsigned(95,8) ,
60176	 => std_logic_vector(to_unsigned(56,8) ,
60177	 => std_logic_vector(to_unsigned(58,8) ,
60178	 => std_logic_vector(to_unsigned(71,8) ,
60179	 => std_logic_vector(to_unsigned(67,8) ,
60180	 => std_logic_vector(to_unsigned(70,8) ,
60181	 => std_logic_vector(to_unsigned(41,8) ,
60182	 => std_logic_vector(to_unsigned(30,8) ,
60183	 => std_logic_vector(to_unsigned(30,8) ,
60184	 => std_logic_vector(to_unsigned(32,8) ,
60185	 => std_logic_vector(to_unsigned(67,8) ,
60186	 => std_logic_vector(to_unsigned(64,8) ,
60187	 => std_logic_vector(to_unsigned(46,8) ,
60188	 => std_logic_vector(to_unsigned(47,8) ,
60189	 => std_logic_vector(to_unsigned(43,8) ,
60190	 => std_logic_vector(to_unsigned(44,8) ,
60191	 => std_logic_vector(to_unsigned(37,8) ,
60192	 => std_logic_vector(to_unsigned(32,8) ,
60193	 => std_logic_vector(to_unsigned(40,8) ,
60194	 => std_logic_vector(to_unsigned(52,8) ,
60195	 => std_logic_vector(to_unsigned(44,8) ,
60196	 => std_logic_vector(to_unsigned(48,8) ,
60197	 => std_logic_vector(to_unsigned(55,8) ,
60198	 => std_logic_vector(to_unsigned(47,8) ,
60199	 => std_logic_vector(to_unsigned(60,8) ,
60200	 => std_logic_vector(to_unsigned(54,8) ,
60201	 => std_logic_vector(to_unsigned(57,8) ,
60202	 => std_logic_vector(to_unsigned(69,8) ,
60203	 => std_logic_vector(to_unsigned(61,8) ,
60204	 => std_logic_vector(to_unsigned(68,8) ,
60205	 => std_logic_vector(to_unsigned(69,8) ,
60206	 => std_logic_vector(to_unsigned(70,8) ,
60207	 => std_logic_vector(to_unsigned(78,8) ,
60208	 => std_logic_vector(to_unsigned(76,8) ,
60209	 => std_logic_vector(to_unsigned(57,8) ,
60210	 => std_logic_vector(to_unsigned(49,8) ,
60211	 => std_logic_vector(to_unsigned(49,8) ,
60212	 => std_logic_vector(to_unsigned(46,8) ,
60213	 => std_logic_vector(to_unsigned(49,8) ,
60214	 => std_logic_vector(to_unsigned(44,8) ,
60215	 => std_logic_vector(to_unsigned(52,8) ,
60216	 => std_logic_vector(to_unsigned(47,8) ,
60217	 => std_logic_vector(to_unsigned(48,8) ,
60218	 => std_logic_vector(to_unsigned(42,8) ,
60219	 => std_logic_vector(to_unsigned(47,8) ,
60220	 => std_logic_vector(to_unsigned(55,8) ,
60221	 => std_logic_vector(to_unsigned(50,8) ,
60222	 => std_logic_vector(to_unsigned(53,8) ,
60223	 => std_logic_vector(to_unsigned(88,8) ,
60224	 => std_logic_vector(to_unsigned(73,8) ,
60225	 => std_logic_vector(to_unsigned(85,8) ,
60226	 => std_logic_vector(to_unsigned(80,8) ,
60227	 => std_logic_vector(to_unsigned(79,8) ,
60228	 => std_logic_vector(to_unsigned(90,8) ,
60229	 => std_logic_vector(to_unsigned(91,8) ,
60230	 => std_logic_vector(to_unsigned(107,8) ,
60231	 => std_logic_vector(to_unsigned(107,8) ,
60232	 => std_logic_vector(to_unsigned(96,8) ,
60233	 => std_logic_vector(to_unsigned(99,8) ,
60234	 => std_logic_vector(to_unsigned(133,8) ,
60235	 => std_logic_vector(to_unsigned(141,8) ,
60236	 => std_logic_vector(to_unsigned(134,8) ,
60237	 => std_logic_vector(to_unsigned(112,8) ,
60238	 => std_logic_vector(to_unsigned(125,8) ,
60239	 => std_logic_vector(to_unsigned(133,8) ,
60240	 => std_logic_vector(to_unsigned(118,8) ,
60241	 => std_logic_vector(to_unsigned(116,8) ,
60242	 => std_logic_vector(to_unsigned(115,8) ,
60243	 => std_logic_vector(to_unsigned(115,8) ,
60244	 => std_logic_vector(to_unsigned(99,8) ,
60245	 => std_logic_vector(to_unsigned(121,8) ,
60246	 => std_logic_vector(to_unsigned(107,8) ,
60247	 => std_logic_vector(to_unsigned(40,8) ,
60248	 => std_logic_vector(to_unsigned(36,8) ,
60249	 => std_logic_vector(to_unsigned(40,8) ,
60250	 => std_logic_vector(to_unsigned(36,8) ,
60251	 => std_logic_vector(to_unsigned(45,8) ,
60252	 => std_logic_vector(to_unsigned(34,8) ,
60253	 => std_logic_vector(to_unsigned(47,8) ,
60254	 => std_logic_vector(to_unsigned(51,8) ,
60255	 => std_logic_vector(to_unsigned(68,8) ,
60256	 => std_logic_vector(to_unsigned(74,8) ,
60257	 => std_logic_vector(to_unsigned(53,8) ,
60258	 => std_logic_vector(to_unsigned(58,8) ,
60259	 => std_logic_vector(to_unsigned(74,8) ,
60260	 => std_logic_vector(to_unsigned(65,8) ,
60261	 => std_logic_vector(to_unsigned(53,8) ,
60262	 => std_logic_vector(to_unsigned(57,8) ,
60263	 => std_logic_vector(to_unsigned(54,8) ,
60264	 => std_logic_vector(to_unsigned(52,8) ,
60265	 => std_logic_vector(to_unsigned(72,8) ,
60266	 => std_logic_vector(to_unsigned(87,8) ,
60267	 => std_logic_vector(to_unsigned(86,8) ,
60268	 => std_logic_vector(to_unsigned(56,8) ,
60269	 => std_logic_vector(to_unsigned(35,8) ,
60270	 => std_logic_vector(to_unsigned(37,8) ,
60271	 => std_logic_vector(to_unsigned(40,8) ,
60272	 => std_logic_vector(to_unsigned(46,8) ,
60273	 => std_logic_vector(to_unsigned(61,8) ,
60274	 => std_logic_vector(to_unsigned(45,8) ,
60275	 => std_logic_vector(to_unsigned(41,8) ,
60276	 => std_logic_vector(to_unsigned(49,8) ,
60277	 => std_logic_vector(to_unsigned(51,8) ,
60278	 => std_logic_vector(to_unsigned(57,8) ,
60279	 => std_logic_vector(to_unsigned(62,8) ,
60280	 => std_logic_vector(to_unsigned(67,8) ,
60281	 => std_logic_vector(to_unsigned(82,8) ,
60282	 => std_logic_vector(to_unsigned(79,8) ,
60283	 => std_logic_vector(to_unsigned(81,8) ,
60284	 => std_logic_vector(to_unsigned(88,8) ,
60285	 => std_logic_vector(to_unsigned(66,8) ,
60286	 => std_logic_vector(to_unsigned(30,8) ,
60287	 => std_logic_vector(to_unsigned(42,8) ,
60288	 => std_logic_vector(to_unsigned(35,8) ,
60289	 => std_logic_vector(to_unsigned(32,8) ,
60290	 => std_logic_vector(to_unsigned(45,8) ,
60291	 => std_logic_vector(to_unsigned(17,8) ,
60292	 => std_logic_vector(to_unsigned(21,8) ,
60293	 => std_logic_vector(to_unsigned(15,8) ,
60294	 => std_logic_vector(to_unsigned(18,8) ,
60295	 => std_logic_vector(to_unsigned(18,8) ,
60296	 => std_logic_vector(to_unsigned(10,8) ,
60297	 => std_logic_vector(to_unsigned(16,8) ,
60298	 => std_logic_vector(to_unsigned(19,8) ,
60299	 => std_logic_vector(to_unsigned(18,8) ,
60300	 => std_logic_vector(to_unsigned(16,8) ,
60301	 => std_logic_vector(to_unsigned(14,8) ,
60302	 => std_logic_vector(to_unsigned(14,8) ,
60303	 => std_logic_vector(to_unsigned(24,8) ,
60304	 => std_logic_vector(to_unsigned(82,8) ,
60305	 => std_logic_vector(to_unsigned(91,8) ,
60306	 => std_logic_vector(to_unsigned(61,8) ,
60307	 => std_logic_vector(to_unsigned(124,8) ,
60308	 => std_logic_vector(to_unsigned(93,8) ,
60309	 => std_logic_vector(to_unsigned(78,8) ,
60310	 => std_logic_vector(to_unsigned(74,8) ,
60311	 => std_logic_vector(to_unsigned(54,8) ,
60312	 => std_logic_vector(to_unsigned(37,8) ,
60313	 => std_logic_vector(to_unsigned(37,8) ,
60314	 => std_logic_vector(to_unsigned(30,8) ,
60315	 => std_logic_vector(to_unsigned(29,8) ,
60316	 => std_logic_vector(to_unsigned(35,8) ,
60317	 => std_logic_vector(to_unsigned(38,8) ,
60318	 => std_logic_vector(to_unsigned(64,8) ,
60319	 => std_logic_vector(to_unsigned(77,8) ,
60320	 => std_logic_vector(to_unsigned(119,8) ,
60321	 => std_logic_vector(to_unsigned(146,8) ,
60322	 => std_logic_vector(to_unsigned(105,8) ,
60323	 => std_logic_vector(to_unsigned(40,8) ,
60324	 => std_logic_vector(to_unsigned(20,8) ,
60325	 => std_logic_vector(to_unsigned(9,8) ,
60326	 => std_logic_vector(to_unsigned(7,8) ,
60327	 => std_logic_vector(to_unsigned(10,8) ,
60328	 => std_logic_vector(to_unsigned(36,8) ,
60329	 => std_logic_vector(to_unsigned(39,8) ,
60330	 => std_logic_vector(to_unsigned(34,8) ,
60331	 => std_logic_vector(to_unsigned(39,8) ,
60332	 => std_logic_vector(to_unsigned(39,8) ,
60333	 => std_logic_vector(to_unsigned(44,8) ,
60334	 => std_logic_vector(to_unsigned(67,8) ,
60335	 => std_logic_vector(to_unsigned(95,8) ,
60336	 => std_logic_vector(to_unsigned(92,8) ,
60337	 => std_logic_vector(to_unsigned(32,8) ,
60338	 => std_logic_vector(to_unsigned(20,8) ,
60339	 => std_logic_vector(to_unsigned(59,8) ,
60340	 => std_logic_vector(to_unsigned(66,8) ,
60341	 => std_logic_vector(to_unsigned(29,8) ,
60342	 => std_logic_vector(to_unsigned(8,8) ,
60343	 => std_logic_vector(to_unsigned(9,8) ,
60344	 => std_logic_vector(to_unsigned(12,8) ,
60345	 => std_logic_vector(to_unsigned(22,8) ,
60346	 => std_logic_vector(to_unsigned(18,8) ,
60347	 => std_logic_vector(to_unsigned(20,8) ,
60348	 => std_logic_vector(to_unsigned(30,8) ,
60349	 => std_logic_vector(to_unsigned(37,8) ,
60350	 => std_logic_vector(to_unsigned(39,8) ,
60351	 => std_logic_vector(to_unsigned(38,8) ,
60352	 => std_logic_vector(to_unsigned(37,8) ,
60353	 => std_logic_vector(to_unsigned(50,8) ,
60354	 => std_logic_vector(to_unsigned(59,8) ,
60355	 => std_logic_vector(to_unsigned(76,8) ,
60356	 => std_logic_vector(to_unsigned(59,8) ,
60357	 => std_logic_vector(to_unsigned(44,8) ,
60358	 => std_logic_vector(to_unsigned(44,8) ,
60359	 => std_logic_vector(to_unsigned(32,8) ,
60360	 => std_logic_vector(to_unsigned(22,8) ,
60361	 => std_logic_vector(to_unsigned(38,8) ,
60362	 => std_logic_vector(to_unsigned(47,8) ,
60363	 => std_logic_vector(to_unsigned(39,8) ,
60364	 => std_logic_vector(to_unsigned(29,8) ,
60365	 => std_logic_vector(to_unsigned(32,8) ,
60366	 => std_logic_vector(to_unsigned(33,8) ,
60367	 => std_logic_vector(to_unsigned(37,8) ,
60368	 => std_logic_vector(to_unsigned(35,8) ,
60369	 => std_logic_vector(to_unsigned(24,8) ,
60370	 => std_logic_vector(to_unsigned(18,8) ,
60371	 => std_logic_vector(to_unsigned(17,8) ,
60372	 => std_logic_vector(to_unsigned(17,8) ,
60373	 => std_logic_vector(to_unsigned(22,8) ,
60374	 => std_logic_vector(to_unsigned(24,8) ,
60375	 => std_logic_vector(to_unsigned(31,8) ,
60376	 => std_logic_vector(to_unsigned(48,8) ,
60377	 => std_logic_vector(to_unsigned(45,8) ,
60378	 => std_logic_vector(to_unsigned(26,8) ,
60379	 => std_logic_vector(to_unsigned(17,8) ,
60380	 => std_logic_vector(to_unsigned(22,8) ,
60381	 => std_logic_vector(to_unsigned(21,8) ,
60382	 => std_logic_vector(to_unsigned(25,8) ,
60383	 => std_logic_vector(to_unsigned(45,8) ,
60384	 => std_logic_vector(to_unsigned(57,8) ,
60385	 => std_logic_vector(to_unsigned(16,8) ,
60386	 => std_logic_vector(to_unsigned(19,8) ,
60387	 => std_logic_vector(to_unsigned(32,8) ,
60388	 => std_logic_vector(to_unsigned(44,8) ,
60389	 => std_logic_vector(to_unsigned(53,8) ,
60390	 => std_logic_vector(to_unsigned(47,8) ,
60391	 => std_logic_vector(to_unsigned(29,8) ,
60392	 => std_logic_vector(to_unsigned(26,8) ,
60393	 => std_logic_vector(to_unsigned(51,8) ,
60394	 => std_logic_vector(to_unsigned(41,8) ,
60395	 => std_logic_vector(to_unsigned(35,8) ,
60396	 => std_logic_vector(to_unsigned(30,8) ,
60397	 => std_logic_vector(to_unsigned(32,8) ,
60398	 => std_logic_vector(to_unsigned(34,8) ,
60399	 => std_logic_vector(to_unsigned(33,8) ,
60400	 => std_logic_vector(to_unsigned(51,8) ,
60401	 => std_logic_vector(to_unsigned(71,8) ,
60402	 => std_logic_vector(to_unsigned(73,8) ,
60403	 => std_logic_vector(to_unsigned(80,8) ,
60404	 => std_logic_vector(to_unsigned(90,8) ,
60405	 => std_logic_vector(to_unsigned(45,8) ,
60406	 => std_logic_vector(to_unsigned(32,8) ,
60407	 => std_logic_vector(to_unsigned(64,8) ,
60408	 => std_logic_vector(to_unsigned(96,8) ,
60409	 => std_logic_vector(to_unsigned(52,8) ,
60410	 => std_logic_vector(to_unsigned(22,8) ,
60411	 => std_logic_vector(to_unsigned(13,8) ,
60412	 => std_logic_vector(to_unsigned(15,8) ,
60413	 => std_logic_vector(to_unsigned(17,8) ,
60414	 => std_logic_vector(to_unsigned(11,8) ,
60415	 => std_logic_vector(to_unsigned(15,8) ,
60416	 => std_logic_vector(to_unsigned(12,8) ,
60417	 => std_logic_vector(to_unsigned(8,8) ,
60418	 => std_logic_vector(to_unsigned(12,8) ,
60419	 => std_logic_vector(to_unsigned(19,8) ,
60420	 => std_logic_vector(to_unsigned(22,8) ,
60421	 => std_logic_vector(to_unsigned(13,8) ,
60422	 => std_logic_vector(to_unsigned(20,8) ,
60423	 => std_logic_vector(to_unsigned(25,8) ,
60424	 => std_logic_vector(to_unsigned(27,8) ,
60425	 => std_logic_vector(to_unsigned(10,8) ,
60426	 => std_logic_vector(to_unsigned(0,8) ,
60427	 => std_logic_vector(to_unsigned(1,8) ,
60428	 => std_logic_vector(to_unsigned(10,8) ,
60429	 => std_logic_vector(to_unsigned(20,8) ,
60430	 => std_logic_vector(to_unsigned(17,8) ,
60431	 => std_logic_vector(to_unsigned(21,8) ,
60432	 => std_logic_vector(to_unsigned(29,8) ,
60433	 => std_logic_vector(to_unsigned(26,8) ,
60434	 => std_logic_vector(to_unsigned(23,8) ,
60435	 => std_logic_vector(to_unsigned(16,8) ,
60436	 => std_logic_vector(to_unsigned(11,8) ,
60437	 => std_logic_vector(to_unsigned(8,8) ,
60438	 => std_logic_vector(to_unsigned(10,8) ,
60439	 => std_logic_vector(to_unsigned(16,8) ,
60440	 => std_logic_vector(to_unsigned(16,8) ,
60441	 => std_logic_vector(to_unsigned(23,8) ,
60442	 => std_logic_vector(to_unsigned(16,8) ,
60443	 => std_logic_vector(to_unsigned(11,8) ,
60444	 => std_logic_vector(to_unsigned(2,8) ,
60445	 => std_logic_vector(to_unsigned(0,8) ,
60446	 => std_logic_vector(to_unsigned(2,8) ,
60447	 => std_logic_vector(to_unsigned(3,8) ,
60448	 => std_logic_vector(to_unsigned(0,8) ,
60449	 => std_logic_vector(to_unsigned(0,8) ,
60450	 => std_logic_vector(to_unsigned(14,8) ,
60451	 => std_logic_vector(to_unsigned(24,8) ,
60452	 => std_logic_vector(to_unsigned(20,8) ,
60453	 => std_logic_vector(to_unsigned(33,8) ,
60454	 => std_logic_vector(to_unsigned(27,8) ,
60455	 => std_logic_vector(to_unsigned(24,8) ,
60456	 => std_logic_vector(to_unsigned(13,8) ,
60457	 => std_logic_vector(to_unsigned(4,8) ,
60458	 => std_logic_vector(to_unsigned(10,8) ,
60459	 => std_logic_vector(to_unsigned(26,8) ,
60460	 => std_logic_vector(to_unsigned(35,8) ,
60461	 => std_logic_vector(to_unsigned(35,8) ,
60462	 => std_logic_vector(to_unsigned(10,8) ,
60463	 => std_logic_vector(to_unsigned(9,8) ,
60464	 => std_logic_vector(to_unsigned(9,8) ,
60465	 => std_logic_vector(to_unsigned(7,8) ,
60466	 => std_logic_vector(to_unsigned(11,8) ,
60467	 => std_logic_vector(to_unsigned(12,8) ,
60468	 => std_logic_vector(to_unsigned(11,8) ,
60469	 => std_logic_vector(to_unsigned(9,8) ,
60470	 => std_logic_vector(to_unsigned(5,8) ,
60471	 => std_logic_vector(to_unsigned(5,8) ,
60472	 => std_logic_vector(to_unsigned(6,8) ,
60473	 => std_logic_vector(to_unsigned(8,8) ,
60474	 => std_logic_vector(to_unsigned(8,8) ,
60475	 => std_logic_vector(to_unsigned(8,8) ,
60476	 => std_logic_vector(to_unsigned(10,8) ,
60477	 => std_logic_vector(to_unsigned(9,8) ,
60478	 => std_logic_vector(to_unsigned(14,8) ,
60479	 => std_logic_vector(to_unsigned(13,8) ,
60480	 => std_logic_vector(to_unsigned(19,8) ,
60481	 => std_logic_vector(to_unsigned(74,8) ,
60482	 => std_logic_vector(to_unsigned(91,8) ,
60483	 => std_logic_vector(to_unsigned(79,8) ,
60484	 => std_logic_vector(to_unsigned(65,8) ,
60485	 => std_logic_vector(to_unsigned(67,8) ,
60486	 => std_logic_vector(to_unsigned(41,8) ,
60487	 => std_logic_vector(to_unsigned(34,8) ,
60488	 => std_logic_vector(to_unsigned(41,8) ,
60489	 => std_logic_vector(to_unsigned(54,8) ,
60490	 => std_logic_vector(to_unsigned(51,8) ,
60491	 => std_logic_vector(to_unsigned(53,8) ,
60492	 => std_logic_vector(to_unsigned(51,8) ,
60493	 => std_logic_vector(to_unsigned(47,8) ,
60494	 => std_logic_vector(to_unsigned(66,8) ,
60495	 => std_logic_vector(to_unsigned(85,8) ,
60496	 => std_logic_vector(to_unsigned(65,8) ,
60497	 => std_logic_vector(to_unsigned(65,8) ,
60498	 => std_logic_vector(to_unsigned(69,8) ,
60499	 => std_logic_vector(to_unsigned(57,8) ,
60500	 => std_logic_vector(to_unsigned(53,8) ,
60501	 => std_logic_vector(to_unsigned(56,8) ,
60502	 => std_logic_vector(to_unsigned(44,8) ,
60503	 => std_logic_vector(to_unsigned(38,8) ,
60504	 => std_logic_vector(to_unsigned(25,8) ,
60505	 => std_logic_vector(to_unsigned(52,8) ,
60506	 => std_logic_vector(to_unsigned(64,8) ,
60507	 => std_logic_vector(to_unsigned(46,8) ,
60508	 => std_logic_vector(to_unsigned(44,8) ,
60509	 => std_logic_vector(to_unsigned(41,8) ,
60510	 => std_logic_vector(to_unsigned(45,8) ,
60511	 => std_logic_vector(to_unsigned(41,8) ,
60512	 => std_logic_vector(to_unsigned(35,8) ,
60513	 => std_logic_vector(to_unsigned(43,8) ,
60514	 => std_logic_vector(to_unsigned(43,8) ,
60515	 => std_logic_vector(to_unsigned(41,8) ,
60516	 => std_logic_vector(to_unsigned(45,8) ,
60517	 => std_logic_vector(to_unsigned(48,8) ,
60518	 => std_logic_vector(to_unsigned(46,8) ,
60519	 => std_logic_vector(to_unsigned(54,8) ,
60520	 => std_logic_vector(to_unsigned(52,8) ,
60521	 => std_logic_vector(to_unsigned(57,8) ,
60522	 => std_logic_vector(to_unsigned(68,8) ,
60523	 => std_logic_vector(to_unsigned(69,8) ,
60524	 => std_logic_vector(to_unsigned(64,8) ,
60525	 => std_logic_vector(to_unsigned(64,8) ,
60526	 => std_logic_vector(to_unsigned(68,8) ,
60527	 => std_logic_vector(to_unsigned(78,8) ,
60528	 => std_logic_vector(to_unsigned(59,8) ,
60529	 => std_logic_vector(to_unsigned(46,8) ,
60530	 => std_logic_vector(to_unsigned(52,8) ,
60531	 => std_logic_vector(to_unsigned(51,8) ,
60532	 => std_logic_vector(to_unsigned(42,8) ,
60533	 => std_logic_vector(to_unsigned(43,8) ,
60534	 => std_logic_vector(to_unsigned(45,8) ,
60535	 => std_logic_vector(to_unsigned(45,8) ,
60536	 => std_logic_vector(to_unsigned(46,8) ,
60537	 => std_logic_vector(to_unsigned(68,8) ,
60538	 => std_logic_vector(to_unsigned(68,8) ,
60539	 => std_logic_vector(to_unsigned(60,8) ,
60540	 => std_logic_vector(to_unsigned(51,8) ,
60541	 => std_logic_vector(to_unsigned(47,8) ,
60542	 => std_logic_vector(to_unsigned(51,8) ,
60543	 => std_logic_vector(to_unsigned(90,8) ,
60544	 => std_logic_vector(to_unsigned(80,8) ,
60545	 => std_logic_vector(to_unsigned(93,8) ,
60546	 => std_logic_vector(to_unsigned(84,8) ,
60547	 => std_logic_vector(to_unsigned(71,8) ,
60548	 => std_logic_vector(to_unsigned(104,8) ,
60549	 => std_logic_vector(to_unsigned(70,8) ,
60550	 => std_logic_vector(to_unsigned(81,8) ,
60551	 => std_logic_vector(to_unsigned(115,8) ,
60552	 => std_logic_vector(to_unsigned(88,8) ,
60553	 => std_logic_vector(to_unsigned(104,8) ,
60554	 => std_logic_vector(to_unsigned(142,8) ,
60555	 => std_logic_vector(to_unsigned(146,8) ,
60556	 => std_logic_vector(to_unsigned(139,8) ,
60557	 => std_logic_vector(to_unsigned(133,8) ,
60558	 => std_logic_vector(to_unsigned(133,8) ,
60559	 => std_logic_vector(to_unsigned(121,8) ,
60560	 => std_logic_vector(to_unsigned(109,8) ,
60561	 => std_logic_vector(to_unsigned(118,8) ,
60562	 => std_logic_vector(to_unsigned(115,8) ,
60563	 => std_logic_vector(to_unsigned(108,8) ,
60564	 => std_logic_vector(to_unsigned(100,8) ,
60565	 => std_logic_vector(to_unsigned(118,8) ,
60566	 => std_logic_vector(to_unsigned(108,8) ,
60567	 => std_logic_vector(to_unsigned(44,8) ,
60568	 => std_logic_vector(to_unsigned(36,8) ,
60569	 => std_logic_vector(to_unsigned(39,8) ,
60570	 => std_logic_vector(to_unsigned(33,8) ,
60571	 => std_logic_vector(to_unsigned(38,8) ,
60572	 => std_logic_vector(to_unsigned(29,8) ,
60573	 => std_logic_vector(to_unsigned(44,8) ,
60574	 => std_logic_vector(to_unsigned(42,8) ,
60575	 => std_logic_vector(to_unsigned(52,8) ,
60576	 => std_logic_vector(to_unsigned(62,8) ,
60577	 => std_logic_vector(to_unsigned(66,8) ,
60578	 => std_logic_vector(to_unsigned(61,8) ,
60579	 => std_logic_vector(to_unsigned(66,8) ,
60580	 => std_logic_vector(to_unsigned(72,8) ,
60581	 => std_logic_vector(to_unsigned(67,8) ,
60582	 => std_logic_vector(to_unsigned(61,8) ,
60583	 => std_logic_vector(to_unsigned(60,8) ,
60584	 => std_logic_vector(to_unsigned(58,8) ,
60585	 => std_logic_vector(to_unsigned(62,8) ,
60586	 => std_logic_vector(to_unsigned(65,8) ,
60587	 => std_logic_vector(to_unsigned(85,8) ,
60588	 => std_logic_vector(to_unsigned(62,8) ,
60589	 => std_logic_vector(to_unsigned(41,8) ,
60590	 => std_logic_vector(to_unsigned(38,8) ,
60591	 => std_logic_vector(to_unsigned(37,8) ,
60592	 => std_logic_vector(to_unsigned(48,8) ,
60593	 => std_logic_vector(to_unsigned(67,8) ,
60594	 => std_logic_vector(to_unsigned(42,8) ,
60595	 => std_logic_vector(to_unsigned(41,8) ,
60596	 => std_logic_vector(to_unsigned(64,8) ,
60597	 => std_logic_vector(to_unsigned(86,8) ,
60598	 => std_logic_vector(to_unsigned(68,8) ,
60599	 => std_logic_vector(to_unsigned(50,8) ,
60600	 => std_logic_vector(to_unsigned(45,8) ,
60601	 => std_logic_vector(to_unsigned(64,8) ,
60602	 => std_logic_vector(to_unsigned(70,8) ,
60603	 => std_logic_vector(to_unsigned(74,8) ,
60604	 => std_logic_vector(to_unsigned(76,8) ,
60605	 => std_logic_vector(to_unsigned(82,8) ,
60606	 => std_logic_vector(to_unsigned(67,8) ,
60607	 => std_logic_vector(to_unsigned(49,8) ,
60608	 => std_logic_vector(to_unsigned(46,8) ,
60609	 => std_logic_vector(to_unsigned(41,8) ,
60610	 => std_logic_vector(to_unsigned(36,8) ,
60611	 => std_logic_vector(to_unsigned(18,8) ,
60612	 => std_logic_vector(to_unsigned(24,8) ,
60613	 => std_logic_vector(to_unsigned(17,8) ,
60614	 => std_logic_vector(to_unsigned(23,8) ,
60615	 => std_logic_vector(to_unsigned(30,8) ,
60616	 => std_logic_vector(to_unsigned(16,8) ,
60617	 => std_logic_vector(to_unsigned(17,8) ,
60618	 => std_logic_vector(to_unsigned(18,8) ,
60619	 => std_logic_vector(to_unsigned(16,8) ,
60620	 => std_logic_vector(to_unsigned(17,8) ,
60621	 => std_logic_vector(to_unsigned(24,8) ,
60622	 => std_logic_vector(to_unsigned(28,8) ,
60623	 => std_logic_vector(to_unsigned(38,8) ,
60624	 => std_logic_vector(to_unsigned(56,8) ,
60625	 => std_logic_vector(to_unsigned(49,8) ,
60626	 => std_logic_vector(to_unsigned(44,8) ,
60627	 => std_logic_vector(to_unsigned(109,8) ,
60628	 => std_logic_vector(to_unsigned(99,8) ,
60629	 => std_logic_vector(to_unsigned(56,8) ,
60630	 => std_logic_vector(to_unsigned(95,8) ,
60631	 => std_logic_vector(to_unsigned(105,8) ,
60632	 => std_logic_vector(to_unsigned(87,8) ,
60633	 => std_logic_vector(to_unsigned(82,8) ,
60634	 => std_logic_vector(to_unsigned(67,8) ,
60635	 => std_logic_vector(to_unsigned(55,8) ,
60636	 => std_logic_vector(to_unsigned(47,8) ,
60637	 => std_logic_vector(to_unsigned(91,8) ,
60638	 => std_logic_vector(to_unsigned(119,8) ,
60639	 => std_logic_vector(to_unsigned(56,8) ,
60640	 => std_logic_vector(to_unsigned(57,8) ,
60641	 => std_logic_vector(to_unsigned(82,8) ,
60642	 => std_logic_vector(to_unsigned(52,8) ,
60643	 => std_logic_vector(to_unsigned(7,8) ,
60644	 => std_logic_vector(to_unsigned(31,8) ,
60645	 => std_logic_vector(to_unsigned(25,8) ,
60646	 => std_logic_vector(to_unsigned(22,8) ,
60647	 => std_logic_vector(to_unsigned(33,8) ,
60648	 => std_logic_vector(to_unsigned(48,8) ,
60649	 => std_logic_vector(to_unsigned(41,8) ,
60650	 => std_logic_vector(to_unsigned(32,8) ,
60651	 => std_logic_vector(to_unsigned(37,8) ,
60652	 => std_logic_vector(to_unsigned(39,8) ,
60653	 => std_logic_vector(to_unsigned(49,8) ,
60654	 => std_logic_vector(to_unsigned(90,8) ,
60655	 => std_logic_vector(to_unsigned(76,8) ,
60656	 => std_logic_vector(to_unsigned(51,8) ,
60657	 => std_logic_vector(to_unsigned(58,8) ,
60658	 => std_logic_vector(to_unsigned(62,8) ,
60659	 => std_logic_vector(to_unsigned(61,8) ,
60660	 => std_logic_vector(to_unsigned(48,8) ,
60661	 => std_logic_vector(to_unsigned(17,8) ,
60662	 => std_logic_vector(to_unsigned(8,8) ,
60663	 => std_logic_vector(to_unsigned(11,8) ,
60664	 => std_logic_vector(to_unsigned(12,8) ,
60665	 => std_logic_vector(to_unsigned(12,8) ,
60666	 => std_logic_vector(to_unsigned(11,8) ,
60667	 => std_logic_vector(to_unsigned(17,8) ,
60668	 => std_logic_vector(to_unsigned(41,8) ,
60669	 => std_logic_vector(to_unsigned(42,8) ,
60670	 => std_logic_vector(to_unsigned(27,8) ,
60671	 => std_logic_vector(to_unsigned(42,8) ,
60672	 => std_logic_vector(to_unsigned(53,8) ,
60673	 => std_logic_vector(to_unsigned(32,8) ,
60674	 => std_logic_vector(to_unsigned(22,8) ,
60675	 => std_logic_vector(to_unsigned(35,8) ,
60676	 => std_logic_vector(to_unsigned(51,8) ,
60677	 => std_logic_vector(to_unsigned(45,8) ,
60678	 => std_logic_vector(to_unsigned(45,8) ,
60679	 => std_logic_vector(to_unsigned(33,8) ,
60680	 => std_logic_vector(to_unsigned(27,8) ,
60681	 => std_logic_vector(to_unsigned(32,8) ,
60682	 => std_logic_vector(to_unsigned(29,8) ,
60683	 => std_logic_vector(to_unsigned(29,8) ,
60684	 => std_logic_vector(to_unsigned(34,8) ,
60685	 => std_logic_vector(to_unsigned(34,8) ,
60686	 => std_logic_vector(to_unsigned(57,8) ,
60687	 => std_logic_vector(to_unsigned(80,8) ,
60688	 => std_logic_vector(to_unsigned(68,8) ,
60689	 => std_logic_vector(to_unsigned(27,8) ,
60690	 => std_logic_vector(to_unsigned(23,8) ,
60691	 => std_logic_vector(to_unsigned(8,8) ,
60692	 => std_logic_vector(to_unsigned(14,8) ,
60693	 => std_logic_vector(to_unsigned(34,8) ,
60694	 => std_logic_vector(to_unsigned(23,8) ,
60695	 => std_logic_vector(to_unsigned(43,8) ,
60696	 => std_logic_vector(to_unsigned(81,8) ,
60697	 => std_logic_vector(to_unsigned(87,8) ,
60698	 => std_logic_vector(to_unsigned(55,8) ,
60699	 => std_logic_vector(to_unsigned(20,8) ,
60700	 => std_logic_vector(to_unsigned(28,8) ,
60701	 => std_logic_vector(to_unsigned(32,8) ,
60702	 => std_logic_vector(to_unsigned(31,8) ,
60703	 => std_logic_vector(to_unsigned(24,8) ,
60704	 => std_logic_vector(to_unsigned(34,8) ,
60705	 => std_logic_vector(to_unsigned(28,8) ,
60706	 => std_logic_vector(to_unsigned(24,8) ,
60707	 => std_logic_vector(to_unsigned(29,8) ,
60708	 => std_logic_vector(to_unsigned(32,8) ,
60709	 => std_logic_vector(to_unsigned(59,8) ,
60710	 => std_logic_vector(to_unsigned(50,8) ,
60711	 => std_logic_vector(to_unsigned(15,8) ,
60712	 => std_logic_vector(to_unsigned(23,8) ,
60713	 => std_logic_vector(to_unsigned(57,8) ,
60714	 => std_logic_vector(to_unsigned(59,8) ,
60715	 => std_logic_vector(to_unsigned(61,8) ,
60716	 => std_logic_vector(to_unsigned(62,8) ,
60717	 => std_logic_vector(to_unsigned(65,8) ,
60718	 => std_logic_vector(to_unsigned(63,8) ,
60719	 => std_logic_vector(to_unsigned(52,8) ,
60720	 => std_logic_vector(to_unsigned(39,8) ,
60721	 => std_logic_vector(to_unsigned(41,8) ,
60722	 => std_logic_vector(to_unsigned(41,8) ,
60723	 => std_logic_vector(to_unsigned(25,8) ,
60724	 => std_logic_vector(to_unsigned(32,8) ,
60725	 => std_logic_vector(to_unsigned(30,8) ,
60726	 => std_logic_vector(to_unsigned(20,8) ,
60727	 => std_logic_vector(to_unsigned(41,8) ,
60728	 => std_logic_vector(to_unsigned(65,8) ,
60729	 => std_logic_vector(to_unsigned(34,8) ,
60730	 => std_logic_vector(to_unsigned(10,8) ,
60731	 => std_logic_vector(to_unsigned(10,8) ,
60732	 => std_logic_vector(to_unsigned(11,8) ,
60733	 => std_logic_vector(to_unsigned(12,8) ,
60734	 => std_logic_vector(to_unsigned(11,8) ,
60735	 => std_logic_vector(to_unsigned(10,8) ,
60736	 => std_logic_vector(to_unsigned(10,8) ,
60737	 => std_logic_vector(to_unsigned(9,8) ,
60738	 => std_logic_vector(to_unsigned(9,8) ,
60739	 => std_logic_vector(to_unsigned(11,8) ,
60740	 => std_logic_vector(to_unsigned(11,8) ,
60741	 => std_logic_vector(to_unsigned(10,8) ,
60742	 => std_logic_vector(to_unsigned(13,8) ,
60743	 => std_logic_vector(to_unsigned(17,8) ,
60744	 => std_logic_vector(to_unsigned(22,8) ,
60745	 => std_logic_vector(to_unsigned(17,8) ,
60746	 => std_logic_vector(to_unsigned(1,8) ,
60747	 => std_logic_vector(to_unsigned(0,8) ,
60748	 => std_logic_vector(to_unsigned(4,8) ,
60749	 => std_logic_vector(to_unsigned(32,8) ,
60750	 => std_logic_vector(to_unsigned(35,8) ,
60751	 => std_logic_vector(to_unsigned(35,8) ,
60752	 => std_logic_vector(to_unsigned(37,8) ,
60753	 => std_logic_vector(to_unsigned(25,8) ,
60754	 => std_logic_vector(to_unsigned(18,8) ,
60755	 => std_logic_vector(to_unsigned(18,8) ,
60756	 => std_logic_vector(to_unsigned(8,8) ,
60757	 => std_logic_vector(to_unsigned(10,8) ,
60758	 => std_logic_vector(to_unsigned(8,8) ,
60759	 => std_logic_vector(to_unsigned(9,8) ,
60760	 => std_logic_vector(to_unsigned(12,8) ,
60761	 => std_logic_vector(to_unsigned(13,8) ,
60762	 => std_logic_vector(to_unsigned(13,8) ,
60763	 => std_logic_vector(to_unsigned(14,8) ,
60764	 => std_logic_vector(to_unsigned(3,8) ,
60765	 => std_logic_vector(to_unsigned(0,8) ,
60766	 => std_logic_vector(to_unsigned(2,8) ,
60767	 => std_logic_vector(to_unsigned(7,8) ,
60768	 => std_logic_vector(to_unsigned(1,8) ,
60769	 => std_logic_vector(to_unsigned(0,8) ,
60770	 => std_logic_vector(to_unsigned(16,8) ,
60771	 => std_logic_vector(to_unsigned(29,8) ,
60772	 => std_logic_vector(to_unsigned(22,8) ,
60773	 => std_logic_vector(to_unsigned(32,8) ,
60774	 => std_logic_vector(to_unsigned(25,8) ,
60775	 => std_logic_vector(to_unsigned(14,8) ,
60776	 => std_logic_vector(to_unsigned(10,8) ,
60777	 => std_logic_vector(to_unsigned(10,8) ,
60778	 => std_logic_vector(to_unsigned(12,8) ,
60779	 => std_logic_vector(to_unsigned(11,8) ,
60780	 => std_logic_vector(to_unsigned(10,8) ,
60781	 => std_logic_vector(to_unsigned(29,8) ,
60782	 => std_logic_vector(to_unsigned(20,8) ,
60783	 => std_logic_vector(to_unsigned(13,8) ,
60784	 => std_logic_vector(to_unsigned(18,8) ,
60785	 => std_logic_vector(to_unsigned(22,8) ,
60786	 => std_logic_vector(to_unsigned(18,8) ,
60787	 => std_logic_vector(to_unsigned(8,8) ,
60788	 => std_logic_vector(to_unsigned(6,8) ,
60789	 => std_logic_vector(to_unsigned(6,8) ,
60790	 => std_logic_vector(to_unsigned(3,8) ,
60791	 => std_logic_vector(to_unsigned(4,8) ,
60792	 => std_logic_vector(to_unsigned(6,8) ,
60793	 => std_logic_vector(to_unsigned(7,8) ,
60794	 => std_logic_vector(to_unsigned(8,8) ,
60795	 => std_logic_vector(to_unsigned(10,8) ,
60796	 => std_logic_vector(to_unsigned(13,8) ,
60797	 => std_logic_vector(to_unsigned(12,8) ,
60798	 => std_logic_vector(to_unsigned(12,8) ,
60799	 => std_logic_vector(to_unsigned(14,8) ,
60800	 => std_logic_vector(to_unsigned(18,8) ,
60801	 => std_logic_vector(to_unsigned(71,8) ,
60802	 => std_logic_vector(to_unsigned(93,8) ,
60803	 => std_logic_vector(to_unsigned(78,8) ,
60804	 => std_logic_vector(to_unsigned(57,8) ,
60805	 => std_logic_vector(to_unsigned(67,8) ,
60806	 => std_logic_vector(to_unsigned(47,8) ,
60807	 => std_logic_vector(to_unsigned(35,8) ,
60808	 => std_logic_vector(to_unsigned(39,8) ,
60809	 => std_logic_vector(to_unsigned(56,8) ,
60810	 => std_logic_vector(to_unsigned(52,8) ,
60811	 => std_logic_vector(to_unsigned(48,8) ,
60812	 => std_logic_vector(to_unsigned(46,8) ,
60813	 => std_logic_vector(to_unsigned(47,8) ,
60814	 => std_logic_vector(to_unsigned(48,8) ,
60815	 => std_logic_vector(to_unsigned(45,8) ,
60816	 => std_logic_vector(to_unsigned(43,8) ,
60817	 => std_logic_vector(to_unsigned(41,8) ,
60818	 => std_logic_vector(to_unsigned(37,8) ,
60819	 => std_logic_vector(to_unsigned(51,8) ,
60820	 => std_logic_vector(to_unsigned(51,8) ,
60821	 => std_logic_vector(to_unsigned(44,8) ,
60822	 => std_logic_vector(to_unsigned(41,8) ,
60823	 => std_logic_vector(to_unsigned(30,8) ,
60824	 => std_logic_vector(to_unsigned(22,8) ,
60825	 => std_logic_vector(to_unsigned(45,8) ,
60826	 => std_logic_vector(to_unsigned(52,8) ,
60827	 => std_logic_vector(to_unsigned(45,8) ,
60828	 => std_logic_vector(to_unsigned(38,8) ,
60829	 => std_logic_vector(to_unsigned(33,8) ,
60830	 => std_logic_vector(to_unsigned(42,8) ,
60831	 => std_logic_vector(to_unsigned(39,8) ,
60832	 => std_logic_vector(to_unsigned(29,8) ,
60833	 => std_logic_vector(to_unsigned(38,8) ,
60834	 => std_logic_vector(to_unsigned(53,8) ,
60835	 => std_logic_vector(to_unsigned(53,8) ,
60836	 => std_logic_vector(to_unsigned(52,8) ,
60837	 => std_logic_vector(to_unsigned(49,8) ,
60838	 => std_logic_vector(to_unsigned(42,8) ,
60839	 => std_logic_vector(to_unsigned(48,8) ,
60840	 => std_logic_vector(to_unsigned(42,8) ,
60841	 => std_logic_vector(to_unsigned(45,8) ,
60842	 => std_logic_vector(to_unsigned(52,8) ,
60843	 => std_logic_vector(to_unsigned(60,8) ,
60844	 => std_logic_vector(to_unsigned(58,8) ,
60845	 => std_logic_vector(to_unsigned(55,8) ,
60846	 => std_logic_vector(to_unsigned(62,8) ,
60847	 => std_logic_vector(to_unsigned(65,8) ,
60848	 => std_logic_vector(to_unsigned(53,8) ,
60849	 => std_logic_vector(to_unsigned(51,8) ,
60850	 => std_logic_vector(to_unsigned(54,8) ,
60851	 => std_logic_vector(to_unsigned(45,8) ,
60852	 => std_logic_vector(to_unsigned(39,8) ,
60853	 => std_logic_vector(to_unsigned(38,8) ,
60854	 => std_logic_vector(to_unsigned(46,8) ,
60855	 => std_logic_vector(to_unsigned(55,8) ,
60856	 => std_logic_vector(to_unsigned(74,8) ,
60857	 => std_logic_vector(to_unsigned(95,8) ,
60858	 => std_logic_vector(to_unsigned(85,8) ,
60859	 => std_logic_vector(to_unsigned(68,8) ,
60860	 => std_logic_vector(to_unsigned(60,8) ,
60861	 => std_logic_vector(to_unsigned(48,8) ,
60862	 => std_logic_vector(to_unsigned(51,8) ,
60863	 => std_logic_vector(to_unsigned(90,8) ,
60864	 => std_logic_vector(to_unsigned(103,8) ,
60865	 => std_logic_vector(to_unsigned(85,8) ,
60866	 => std_logic_vector(to_unsigned(91,8) ,
60867	 => std_logic_vector(to_unsigned(93,8) ,
60868	 => std_logic_vector(to_unsigned(103,8) ,
60869	 => std_logic_vector(to_unsigned(82,8) ,
60870	 => std_logic_vector(to_unsigned(88,8) ,
60871	 => std_logic_vector(to_unsigned(114,8) ,
60872	 => std_logic_vector(to_unsigned(71,8) ,
60873	 => std_logic_vector(to_unsigned(90,8) ,
60874	 => std_logic_vector(to_unsigned(146,8) ,
60875	 => std_logic_vector(to_unsigned(138,8) ,
60876	 => std_logic_vector(to_unsigned(128,8) ,
60877	 => std_logic_vector(to_unsigned(127,8) ,
60878	 => std_logic_vector(to_unsigned(125,8) ,
60879	 => std_logic_vector(to_unsigned(122,8) ,
60880	 => std_logic_vector(to_unsigned(112,8) ,
60881	 => std_logic_vector(to_unsigned(116,8) ,
60882	 => std_logic_vector(to_unsigned(105,8) ,
60883	 => std_logic_vector(to_unsigned(109,8) ,
60884	 => std_logic_vector(to_unsigned(119,8) ,
60885	 => std_logic_vector(to_unsigned(122,8) ,
60886	 => std_logic_vector(to_unsigned(115,8) ,
60887	 => std_logic_vector(to_unsigned(41,8) ,
60888	 => std_logic_vector(to_unsigned(29,8) ,
60889	 => std_logic_vector(to_unsigned(37,8) ,
60890	 => std_logic_vector(to_unsigned(41,8) ,
60891	 => std_logic_vector(to_unsigned(38,8) ,
60892	 => std_logic_vector(to_unsigned(35,8) ,
60893	 => std_logic_vector(to_unsigned(40,8) ,
60894	 => std_logic_vector(to_unsigned(38,8) ,
60895	 => std_logic_vector(to_unsigned(53,8) ,
60896	 => std_logic_vector(to_unsigned(49,8) ,
60897	 => std_logic_vector(to_unsigned(51,8) ,
60898	 => std_logic_vector(to_unsigned(65,8) ,
60899	 => std_logic_vector(to_unsigned(53,8) ,
60900	 => std_logic_vector(to_unsigned(69,8) ,
60901	 => std_logic_vector(to_unsigned(96,8) ,
60902	 => std_logic_vector(to_unsigned(67,8) ,
60903	 => std_logic_vector(to_unsigned(48,8) ,
60904	 => std_logic_vector(to_unsigned(62,8) ,
60905	 => std_logic_vector(to_unsigned(50,8) ,
60906	 => std_logic_vector(to_unsigned(47,8) ,
60907	 => std_logic_vector(to_unsigned(62,8) ,
60908	 => std_logic_vector(to_unsigned(54,8) ,
60909	 => std_logic_vector(to_unsigned(45,8) ,
60910	 => std_logic_vector(to_unsigned(39,8) ,
60911	 => std_logic_vector(to_unsigned(41,8) ,
60912	 => std_logic_vector(to_unsigned(51,8) ,
60913	 => std_logic_vector(to_unsigned(59,8) ,
60914	 => std_logic_vector(to_unsigned(52,8) ,
60915	 => std_logic_vector(to_unsigned(81,8) ,
60916	 => std_logic_vector(to_unsigned(76,8) ,
60917	 => std_logic_vector(to_unsigned(67,8) ,
60918	 => std_logic_vector(to_unsigned(51,8) ,
60919	 => std_logic_vector(to_unsigned(34,8) ,
60920	 => std_logic_vector(to_unsigned(37,8) ,
60921	 => std_logic_vector(to_unsigned(57,8) ,
60922	 => std_logic_vector(to_unsigned(65,8) ,
60923	 => std_logic_vector(to_unsigned(41,8) ,
60924	 => std_logic_vector(to_unsigned(53,8) ,
60925	 => std_logic_vector(to_unsigned(73,8) ,
60926	 => std_logic_vector(to_unsigned(80,8) ,
60927	 => std_logic_vector(to_unsigned(31,8) ,
60928	 => std_logic_vector(to_unsigned(34,8) ,
60929	 => std_logic_vector(to_unsigned(36,8) ,
60930	 => std_logic_vector(to_unsigned(29,8) ,
60931	 => std_logic_vector(to_unsigned(27,8) ,
60932	 => std_logic_vector(to_unsigned(36,8) ,
60933	 => std_logic_vector(to_unsigned(23,8) ,
60934	 => std_logic_vector(to_unsigned(24,8) ,
60935	 => std_logic_vector(to_unsigned(31,8) ,
60936	 => std_logic_vector(to_unsigned(22,8) ,
60937	 => std_logic_vector(to_unsigned(16,8) ,
60938	 => std_logic_vector(to_unsigned(14,8) ,
60939	 => std_logic_vector(to_unsigned(17,8) ,
60940	 => std_logic_vector(to_unsigned(17,8) ,
60941	 => std_logic_vector(to_unsigned(19,8) ,
60942	 => std_logic_vector(to_unsigned(27,8) ,
60943	 => std_logic_vector(to_unsigned(23,8) ,
60944	 => std_logic_vector(to_unsigned(14,8) ,
60945	 => std_logic_vector(to_unsigned(14,8) ,
60946	 => std_logic_vector(to_unsigned(19,8) ,
60947	 => std_logic_vector(to_unsigned(23,8) ,
60948	 => std_logic_vector(to_unsigned(24,8) ,
60949	 => std_logic_vector(to_unsigned(25,8) ,
60950	 => std_logic_vector(to_unsigned(51,8) ,
60951	 => std_logic_vector(to_unsigned(80,8) ,
60952	 => std_logic_vector(to_unsigned(54,8) ,
60953	 => std_logic_vector(to_unsigned(154,8) ,
60954	 => std_logic_vector(to_unsigned(136,8) ,
60955	 => std_logic_vector(to_unsigned(73,8) ,
60956	 => std_logic_vector(to_unsigned(112,8) ,
60957	 => std_logic_vector(to_unsigned(130,8) ,
60958	 => std_logic_vector(to_unsigned(73,8) ,
60959	 => std_logic_vector(to_unsigned(37,8) ,
60960	 => std_logic_vector(to_unsigned(19,8) ,
60961	 => std_logic_vector(to_unsigned(16,8) ,
60962	 => std_logic_vector(to_unsigned(18,8) ,
60963	 => std_logic_vector(to_unsigned(12,8) ,
60964	 => std_logic_vector(to_unsigned(17,8) ,
60965	 => std_logic_vector(to_unsigned(19,8) ,
60966	 => std_logic_vector(to_unsigned(24,8) ,
60967	 => std_logic_vector(to_unsigned(30,8) ,
60968	 => std_logic_vector(to_unsigned(22,8) ,
60969	 => std_logic_vector(to_unsigned(23,8) ,
60970	 => std_logic_vector(to_unsigned(35,8) ,
60971	 => std_logic_vector(to_unsigned(32,8) ,
60972	 => std_logic_vector(to_unsigned(66,8) ,
60973	 => std_logic_vector(to_unsigned(95,8) ,
60974	 => std_logic_vector(to_unsigned(39,8) ,
60975	 => std_logic_vector(to_unsigned(22,8) ,
60976	 => std_logic_vector(to_unsigned(29,8) ,
60977	 => std_logic_vector(to_unsigned(60,8) ,
60978	 => std_logic_vector(to_unsigned(61,8) ,
60979	 => std_logic_vector(to_unsigned(54,8) ,
60980	 => std_logic_vector(to_unsigned(49,8) ,
60981	 => std_logic_vector(to_unsigned(13,8) ,
60982	 => std_logic_vector(to_unsigned(8,8) ,
60983	 => std_logic_vector(to_unsigned(12,8) ,
60984	 => std_logic_vector(to_unsigned(16,8) ,
60985	 => std_logic_vector(to_unsigned(17,8) ,
60986	 => std_logic_vector(to_unsigned(14,8) ,
60987	 => std_logic_vector(to_unsigned(30,8) ,
60988	 => std_logic_vector(to_unsigned(38,8) ,
60989	 => std_logic_vector(to_unsigned(26,8) ,
60990	 => std_logic_vector(to_unsigned(33,8) ,
60991	 => std_logic_vector(to_unsigned(42,8) ,
60992	 => std_logic_vector(to_unsigned(45,8) ,
60993	 => std_logic_vector(to_unsigned(43,8) ,
60994	 => std_logic_vector(to_unsigned(37,8) ,
60995	 => std_logic_vector(to_unsigned(34,8) ,
60996	 => std_logic_vector(to_unsigned(53,8) ,
60997	 => std_logic_vector(to_unsigned(52,8) ,
60998	 => std_logic_vector(to_unsigned(45,8) ,
60999	 => std_logic_vector(to_unsigned(42,8) ,
61000	 => std_logic_vector(to_unsigned(39,8) ,
61001	 => std_logic_vector(to_unsigned(41,8) ,
61002	 => std_logic_vector(to_unsigned(48,8) ,
61003	 => std_logic_vector(to_unsigned(39,8) ,
61004	 => std_logic_vector(to_unsigned(35,8) ,
61005	 => std_logic_vector(to_unsigned(39,8) ,
61006	 => std_logic_vector(to_unsigned(51,8) ,
61007	 => std_logic_vector(to_unsigned(69,8) ,
61008	 => std_logic_vector(to_unsigned(65,8) ,
61009	 => std_logic_vector(to_unsigned(29,8) ,
61010	 => std_logic_vector(to_unsigned(23,8) ,
61011	 => std_logic_vector(to_unsigned(17,8) ,
61012	 => std_logic_vector(to_unsigned(21,8) ,
61013	 => std_logic_vector(to_unsigned(29,8) ,
61014	 => std_logic_vector(to_unsigned(27,8) ,
61015	 => std_logic_vector(to_unsigned(43,8) ,
61016	 => std_logic_vector(to_unsigned(67,8) ,
61017	 => std_logic_vector(to_unsigned(72,8) ,
61018	 => std_logic_vector(to_unsigned(56,8) ,
61019	 => std_logic_vector(to_unsigned(30,8) ,
61020	 => std_logic_vector(to_unsigned(34,8) ,
61021	 => std_logic_vector(to_unsigned(57,8) ,
61022	 => std_logic_vector(to_unsigned(34,8) ,
61023	 => std_logic_vector(to_unsigned(11,8) ,
61024	 => std_logic_vector(to_unsigned(19,8) ,
61025	 => std_logic_vector(to_unsigned(31,8) ,
61026	 => std_logic_vector(to_unsigned(36,8) ,
61027	 => std_logic_vector(to_unsigned(37,8) ,
61028	 => std_logic_vector(to_unsigned(37,8) ,
61029	 => std_logic_vector(to_unsigned(43,8) ,
61030	 => std_logic_vector(to_unsigned(30,8) ,
61031	 => std_logic_vector(to_unsigned(10,8) ,
61032	 => std_logic_vector(to_unsigned(17,8) ,
61033	 => std_logic_vector(to_unsigned(27,8) ,
61034	 => std_logic_vector(to_unsigned(21,8) ,
61035	 => std_logic_vector(to_unsigned(32,8) ,
61036	 => std_logic_vector(to_unsigned(37,8) ,
61037	 => std_logic_vector(to_unsigned(44,8) ,
61038	 => std_logic_vector(to_unsigned(56,8) ,
61039	 => std_logic_vector(to_unsigned(62,8) ,
61040	 => std_logic_vector(to_unsigned(60,8) ,
61041	 => std_logic_vector(to_unsigned(70,8) ,
61042	 => std_logic_vector(to_unsigned(71,8) ,
61043	 => std_logic_vector(to_unsigned(57,8) ,
61044	 => std_logic_vector(to_unsigned(55,8) ,
61045	 => std_logic_vector(to_unsigned(46,8) ,
61046	 => std_logic_vector(to_unsigned(44,8) ,
61047	 => std_logic_vector(to_unsigned(34,8) ,
61048	 => std_logic_vector(to_unsigned(23,8) ,
61049	 => std_logic_vector(to_unsigned(17,8) ,
61050	 => std_logic_vector(to_unsigned(10,8) ,
61051	 => std_logic_vector(to_unsigned(9,8) ,
61052	 => std_logic_vector(to_unsigned(11,8) ,
61053	 => std_logic_vector(to_unsigned(16,8) ,
61054	 => std_logic_vector(to_unsigned(13,8) ,
61055	 => std_logic_vector(to_unsigned(13,8) ,
61056	 => std_logic_vector(to_unsigned(12,8) ,
61057	 => std_logic_vector(to_unsigned(11,8) ,
61058	 => std_logic_vector(to_unsigned(15,8) ,
61059	 => std_logic_vector(to_unsigned(12,8) ,
61060	 => std_logic_vector(to_unsigned(16,8) ,
61061	 => std_logic_vector(to_unsigned(12,8) ,
61062	 => std_logic_vector(to_unsigned(10,8) ,
61063	 => std_logic_vector(to_unsigned(10,8) ,
61064	 => std_logic_vector(to_unsigned(11,8) ,
61065	 => std_logic_vector(to_unsigned(11,8) ,
61066	 => std_logic_vector(to_unsigned(3,8) ,
61067	 => std_logic_vector(to_unsigned(0,8) ,
61068	 => std_logic_vector(to_unsigned(1,8) ,
61069	 => std_logic_vector(to_unsigned(13,8) ,
61070	 => std_logic_vector(to_unsigned(18,8) ,
61071	 => std_logic_vector(to_unsigned(18,8) ,
61072	 => std_logic_vector(to_unsigned(20,8) ,
61073	 => std_logic_vector(to_unsigned(19,8) ,
61074	 => std_logic_vector(to_unsigned(23,8) ,
61075	 => std_logic_vector(to_unsigned(14,8) ,
61076	 => std_logic_vector(to_unsigned(5,8) ,
61077	 => std_logic_vector(to_unsigned(8,8) ,
61078	 => std_logic_vector(to_unsigned(8,8) ,
61079	 => std_logic_vector(to_unsigned(6,8) ,
61080	 => std_logic_vector(to_unsigned(6,8) ,
61081	 => std_logic_vector(to_unsigned(6,8) ,
61082	 => std_logic_vector(to_unsigned(5,8) ,
61083	 => std_logic_vector(to_unsigned(12,8) ,
61084	 => std_logic_vector(to_unsigned(5,8) ,
61085	 => std_logic_vector(to_unsigned(0,8) ,
61086	 => std_logic_vector(to_unsigned(1,8) ,
61087	 => std_logic_vector(to_unsigned(13,8) ,
61088	 => std_logic_vector(to_unsigned(3,8) ,
61089	 => std_logic_vector(to_unsigned(0,8) ,
61090	 => std_logic_vector(to_unsigned(2,8) ,
61091	 => std_logic_vector(to_unsigned(17,8) ,
61092	 => std_logic_vector(to_unsigned(25,8) ,
61093	 => std_logic_vector(to_unsigned(23,8) ,
61094	 => std_logic_vector(to_unsigned(16,8) ,
61095	 => std_logic_vector(to_unsigned(6,8) ,
61096	 => std_logic_vector(to_unsigned(8,8) ,
61097	 => std_logic_vector(to_unsigned(10,8) ,
61098	 => std_logic_vector(to_unsigned(11,8) ,
61099	 => std_logic_vector(to_unsigned(7,8) ,
61100	 => std_logic_vector(to_unsigned(10,8) ,
61101	 => std_logic_vector(to_unsigned(14,8) ,
61102	 => std_logic_vector(to_unsigned(20,8) ,
61103	 => std_logic_vector(to_unsigned(27,8) ,
61104	 => std_logic_vector(to_unsigned(14,8) ,
61105	 => std_logic_vector(to_unsigned(12,8) ,
61106	 => std_logic_vector(to_unsigned(13,8) ,
61107	 => std_logic_vector(to_unsigned(10,8) ,
61108	 => std_logic_vector(to_unsigned(8,8) ,
61109	 => std_logic_vector(to_unsigned(8,8) ,
61110	 => std_logic_vector(to_unsigned(4,8) ,
61111	 => std_logic_vector(to_unsigned(3,8) ,
61112	 => std_logic_vector(to_unsigned(5,8) ,
61113	 => std_logic_vector(to_unsigned(7,8) ,
61114	 => std_logic_vector(to_unsigned(8,8) ,
61115	 => std_logic_vector(to_unsigned(9,8) ,
61116	 => std_logic_vector(to_unsigned(10,8) ,
61117	 => std_logic_vector(to_unsigned(12,8) ,
61118	 => std_logic_vector(to_unsigned(11,8) ,
61119	 => std_logic_vector(to_unsigned(13,8) ,
61120	 => std_logic_vector(to_unsigned(23,8) ,
61121	 => std_logic_vector(to_unsigned(65,8) ,
61122	 => std_logic_vector(to_unsigned(92,8) ,
61123	 => std_logic_vector(to_unsigned(79,8) ,
61124	 => std_logic_vector(to_unsigned(59,8) ,
61125	 => std_logic_vector(to_unsigned(73,8) ,
61126	 => std_logic_vector(to_unsigned(51,8) ,
61127	 => std_logic_vector(to_unsigned(32,8) ,
61128	 => std_logic_vector(to_unsigned(35,8) ,
61129	 => std_logic_vector(to_unsigned(46,8) ,
61130	 => std_logic_vector(to_unsigned(51,8) ,
61131	 => std_logic_vector(to_unsigned(51,8) ,
61132	 => std_logic_vector(to_unsigned(45,8) ,
61133	 => std_logic_vector(to_unsigned(41,8) ,
61134	 => std_logic_vector(to_unsigned(32,8) ,
61135	 => std_logic_vector(to_unsigned(30,8) ,
61136	 => std_logic_vector(to_unsigned(32,8) ,
61137	 => std_logic_vector(to_unsigned(24,8) ,
61138	 => std_logic_vector(to_unsigned(24,8) ,
61139	 => std_logic_vector(to_unsigned(34,8) ,
61140	 => std_logic_vector(to_unsigned(40,8) ,
61141	 => std_logic_vector(to_unsigned(33,8) ,
61142	 => std_logic_vector(to_unsigned(31,8) ,
61143	 => std_logic_vector(to_unsigned(32,8) ,
61144	 => std_logic_vector(to_unsigned(21,8) ,
61145	 => std_logic_vector(to_unsigned(32,8) ,
61146	 => std_logic_vector(to_unsigned(51,8) ,
61147	 => std_logic_vector(to_unsigned(37,8) ,
61148	 => std_logic_vector(to_unsigned(43,8) ,
61149	 => std_logic_vector(to_unsigned(40,8) ,
61150	 => std_logic_vector(to_unsigned(43,8) ,
61151	 => std_logic_vector(to_unsigned(34,8) ,
61152	 => std_logic_vector(to_unsigned(26,8) ,
61153	 => std_logic_vector(to_unsigned(35,8) ,
61154	 => std_logic_vector(to_unsigned(65,8) ,
61155	 => std_logic_vector(to_unsigned(57,8) ,
61156	 => std_logic_vector(to_unsigned(71,8) ,
61157	 => std_logic_vector(to_unsigned(79,8) ,
61158	 => std_logic_vector(to_unsigned(36,8) ,
61159	 => std_logic_vector(to_unsigned(51,8) ,
61160	 => std_logic_vector(to_unsigned(59,8) ,
61161	 => std_logic_vector(to_unsigned(37,8) ,
61162	 => std_logic_vector(to_unsigned(44,8) ,
61163	 => std_logic_vector(to_unsigned(51,8) ,
61164	 => std_logic_vector(to_unsigned(55,8) ,
61165	 => std_logic_vector(to_unsigned(61,8) ,
61166	 => std_logic_vector(to_unsigned(58,8) ,
61167	 => std_logic_vector(to_unsigned(59,8) ,
61168	 => std_logic_vector(to_unsigned(58,8) ,
61169	 => std_logic_vector(to_unsigned(51,8) ,
61170	 => std_logic_vector(to_unsigned(49,8) ,
61171	 => std_logic_vector(to_unsigned(41,8) ,
61172	 => std_logic_vector(to_unsigned(35,8) ,
61173	 => std_logic_vector(to_unsigned(47,8) ,
61174	 => std_logic_vector(to_unsigned(53,8) ,
61175	 => std_logic_vector(to_unsigned(51,8) ,
61176	 => std_logic_vector(to_unsigned(59,8) ,
61177	 => std_logic_vector(to_unsigned(69,8) ,
61178	 => std_logic_vector(to_unsigned(69,8) ,
61179	 => std_logic_vector(to_unsigned(52,8) ,
61180	 => std_logic_vector(to_unsigned(53,8) ,
61181	 => std_logic_vector(to_unsigned(53,8) ,
61182	 => std_logic_vector(to_unsigned(61,8) ,
61183	 => std_logic_vector(to_unsigned(104,8) ,
61184	 => std_logic_vector(to_unsigned(122,8) ,
61185	 => std_logic_vector(to_unsigned(112,8) ,
61186	 => std_logic_vector(to_unsigned(85,8) ,
61187	 => std_logic_vector(to_unsigned(67,8) ,
61188	 => std_logic_vector(to_unsigned(92,8) ,
61189	 => std_logic_vector(to_unsigned(96,8) ,
61190	 => std_logic_vector(to_unsigned(97,8) ,
61191	 => std_logic_vector(to_unsigned(101,8) ,
61192	 => std_logic_vector(to_unsigned(101,8) ,
61193	 => std_logic_vector(to_unsigned(105,8) ,
61194	 => std_logic_vector(to_unsigned(139,8) ,
61195	 => std_logic_vector(to_unsigned(128,8) ,
61196	 => std_logic_vector(to_unsigned(116,8) ,
61197	 => std_logic_vector(to_unsigned(124,8) ,
61198	 => std_logic_vector(to_unsigned(131,8) ,
61199	 => std_logic_vector(to_unsigned(122,8) ,
61200	 => std_logic_vector(to_unsigned(107,8) ,
61201	 => std_logic_vector(to_unsigned(116,8) ,
61202	 => std_logic_vector(to_unsigned(119,8) ,
61203	 => std_logic_vector(to_unsigned(115,8) ,
61204	 => std_logic_vector(to_unsigned(103,8) ,
61205	 => std_logic_vector(to_unsigned(119,8) ,
61206	 => std_logic_vector(to_unsigned(121,8) ,
61207	 => std_logic_vector(to_unsigned(47,8) ,
61208	 => std_logic_vector(to_unsigned(24,8) ,
61209	 => std_logic_vector(to_unsigned(30,8) ,
61210	 => std_logic_vector(to_unsigned(30,8) ,
61211	 => std_logic_vector(to_unsigned(36,8) ,
61212	 => std_logic_vector(to_unsigned(41,8) ,
61213	 => std_logic_vector(to_unsigned(41,8) ,
61214	 => std_logic_vector(to_unsigned(49,8) ,
61215	 => std_logic_vector(to_unsigned(51,8) ,
61216	 => std_logic_vector(to_unsigned(46,8) ,
61217	 => std_logic_vector(to_unsigned(51,8) ,
61218	 => std_logic_vector(to_unsigned(65,8) ,
61219	 => std_logic_vector(to_unsigned(61,8) ,
61220	 => std_logic_vector(to_unsigned(78,8) ,
61221	 => std_logic_vector(to_unsigned(108,8) ,
61222	 => std_logic_vector(to_unsigned(79,8) ,
61223	 => std_logic_vector(to_unsigned(56,8) ,
61224	 => std_logic_vector(to_unsigned(53,8) ,
61225	 => std_logic_vector(to_unsigned(50,8) ,
61226	 => std_logic_vector(to_unsigned(51,8) ,
61227	 => std_logic_vector(to_unsigned(52,8) ,
61228	 => std_logic_vector(to_unsigned(54,8) ,
61229	 => std_logic_vector(to_unsigned(53,8) ,
61230	 => std_logic_vector(to_unsigned(45,8) ,
61231	 => std_logic_vector(to_unsigned(52,8) ,
61232	 => std_logic_vector(to_unsigned(45,8) ,
61233	 => std_logic_vector(to_unsigned(51,8) ,
61234	 => std_logic_vector(to_unsigned(92,8) ,
61235	 => std_logic_vector(to_unsigned(97,8) ,
61236	 => std_logic_vector(to_unsigned(71,8) ,
61237	 => std_logic_vector(to_unsigned(50,8) ,
61238	 => std_logic_vector(to_unsigned(33,8) ,
61239	 => std_logic_vector(to_unsigned(45,8) ,
61240	 => std_logic_vector(to_unsigned(60,8) ,
61241	 => std_logic_vector(to_unsigned(51,8) ,
61242	 => std_logic_vector(to_unsigned(40,8) ,
61243	 => std_logic_vector(to_unsigned(35,8) ,
61244	 => std_logic_vector(to_unsigned(57,8) ,
61245	 => std_logic_vector(to_unsigned(74,8) ,
61246	 => std_logic_vector(to_unsigned(45,8) ,
61247	 => std_logic_vector(to_unsigned(38,8) ,
61248	 => std_logic_vector(to_unsigned(55,8) ,
61249	 => std_logic_vector(to_unsigned(59,8) ,
61250	 => std_logic_vector(to_unsigned(55,8) ,
61251	 => std_logic_vector(to_unsigned(27,8) ,
61252	 => std_logic_vector(to_unsigned(32,8) ,
61253	 => std_logic_vector(to_unsigned(26,8) ,
61254	 => std_logic_vector(to_unsigned(20,8) ,
61255	 => std_logic_vector(to_unsigned(27,8) ,
61256	 => std_logic_vector(to_unsigned(30,8) ,
61257	 => std_logic_vector(to_unsigned(28,8) ,
61258	 => std_logic_vector(to_unsigned(16,8) ,
61259	 => std_logic_vector(to_unsigned(22,8) ,
61260	 => std_logic_vector(to_unsigned(32,8) ,
61261	 => std_logic_vector(to_unsigned(30,8) ,
61262	 => std_logic_vector(to_unsigned(27,8) ,
61263	 => std_logic_vector(to_unsigned(30,8) ,
61264	 => std_logic_vector(to_unsigned(30,8) ,
61265	 => std_logic_vector(to_unsigned(22,8) ,
61266	 => std_logic_vector(to_unsigned(22,8) ,
61267	 => std_logic_vector(to_unsigned(17,8) ,
61268	 => std_logic_vector(to_unsigned(15,8) ,
61269	 => std_logic_vector(to_unsigned(20,8) ,
61270	 => std_logic_vector(to_unsigned(30,8) ,
61271	 => std_logic_vector(to_unsigned(64,8) ,
61272	 => std_logic_vector(to_unsigned(72,8) ,
61273	 => std_logic_vector(to_unsigned(154,8) ,
61274	 => std_logic_vector(to_unsigned(122,8) ,
61275	 => std_logic_vector(to_unsigned(43,8) ,
61276	 => std_logic_vector(to_unsigned(121,8) ,
61277	 => std_logic_vector(to_unsigned(90,8) ,
61278	 => std_logic_vector(to_unsigned(25,8) ,
61279	 => std_logic_vector(to_unsigned(31,8) ,
61280	 => std_logic_vector(to_unsigned(49,8) ,
61281	 => std_logic_vector(to_unsigned(58,8) ,
61282	 => std_logic_vector(to_unsigned(51,8) ,
61283	 => std_logic_vector(to_unsigned(45,8) ,
61284	 => std_logic_vector(to_unsigned(10,8) ,
61285	 => std_logic_vector(to_unsigned(11,8) ,
61286	 => std_logic_vector(to_unsigned(10,8) ,
61287	 => std_logic_vector(to_unsigned(22,8) ,
61288	 => std_logic_vector(to_unsigned(39,8) ,
61289	 => std_logic_vector(to_unsigned(29,8) ,
61290	 => std_logic_vector(to_unsigned(20,8) ,
61291	 => std_logic_vector(to_unsigned(32,8) ,
61292	 => std_logic_vector(to_unsigned(68,8) ,
61293	 => std_logic_vector(to_unsigned(109,8) ,
61294	 => std_logic_vector(to_unsigned(17,8) ,
61295	 => std_logic_vector(to_unsigned(19,8) ,
61296	 => std_logic_vector(to_unsigned(57,8) ,
61297	 => std_logic_vector(to_unsigned(59,8) ,
61298	 => std_logic_vector(to_unsigned(51,8) ,
61299	 => std_logic_vector(to_unsigned(61,8) ,
61300	 => std_logic_vector(to_unsigned(85,8) ,
61301	 => std_logic_vector(to_unsigned(13,8) ,
61302	 => std_logic_vector(to_unsigned(6,8) ,
61303	 => std_logic_vector(to_unsigned(12,8) ,
61304	 => std_logic_vector(to_unsigned(12,8) ,
61305	 => std_logic_vector(to_unsigned(10,8) ,
61306	 => std_logic_vector(to_unsigned(21,8) ,
61307	 => std_logic_vector(to_unsigned(47,8) ,
61308	 => std_logic_vector(to_unsigned(10,8) ,
61309	 => std_logic_vector(to_unsigned(4,8) ,
61310	 => std_logic_vector(to_unsigned(26,8) ,
61311	 => std_logic_vector(to_unsigned(44,8) ,
61312	 => std_logic_vector(to_unsigned(29,8) ,
61313	 => std_logic_vector(to_unsigned(35,8) ,
61314	 => std_logic_vector(to_unsigned(41,8) ,
61315	 => std_logic_vector(to_unsigned(47,8) ,
61316	 => std_logic_vector(to_unsigned(44,8) ,
61317	 => std_logic_vector(to_unsigned(45,8) ,
61318	 => std_logic_vector(to_unsigned(56,8) ,
61319	 => std_logic_vector(to_unsigned(42,8) ,
61320	 => std_logic_vector(to_unsigned(32,8) ,
61321	 => std_logic_vector(to_unsigned(52,8) ,
61322	 => std_logic_vector(to_unsigned(63,8) ,
61323	 => std_logic_vector(to_unsigned(53,8) ,
61324	 => std_logic_vector(to_unsigned(33,8) ,
61325	 => std_logic_vector(to_unsigned(40,8) ,
61326	 => std_logic_vector(to_unsigned(45,8) ,
61327	 => std_logic_vector(to_unsigned(42,8) ,
61328	 => std_logic_vector(to_unsigned(36,8) ,
61329	 => std_logic_vector(to_unsigned(32,8) ,
61330	 => std_logic_vector(to_unsigned(23,8) ,
61331	 => std_logic_vector(to_unsigned(24,8) ,
61332	 => std_logic_vector(to_unsigned(30,8) ,
61333	 => std_logic_vector(to_unsigned(30,8) ,
61334	 => std_logic_vector(to_unsigned(33,8) ,
61335	 => std_logic_vector(to_unsigned(41,8) ,
61336	 => std_logic_vector(to_unsigned(53,8) ,
61337	 => std_logic_vector(to_unsigned(55,8) ,
61338	 => std_logic_vector(to_unsigned(44,8) ,
61339	 => std_logic_vector(to_unsigned(37,8) ,
61340	 => std_logic_vector(to_unsigned(37,8) ,
61341	 => std_logic_vector(to_unsigned(39,8) ,
61342	 => std_logic_vector(to_unsigned(36,8) ,
61343	 => std_logic_vector(to_unsigned(37,8) ,
61344	 => std_logic_vector(to_unsigned(35,8) ,
61345	 => std_logic_vector(to_unsigned(36,8) ,
61346	 => std_logic_vector(to_unsigned(41,8) ,
61347	 => std_logic_vector(to_unsigned(47,8) ,
61348	 => std_logic_vector(to_unsigned(53,8) ,
61349	 => std_logic_vector(to_unsigned(32,8) ,
61350	 => std_logic_vector(to_unsigned(29,8) ,
61351	 => std_logic_vector(to_unsigned(24,8) ,
61352	 => std_logic_vector(to_unsigned(27,8) ,
61353	 => std_logic_vector(to_unsigned(20,8) ,
61354	 => std_logic_vector(to_unsigned(17,8) ,
61355	 => std_logic_vector(to_unsigned(17,8) ,
61356	 => std_logic_vector(to_unsigned(15,8) ,
61357	 => std_logic_vector(to_unsigned(12,8) ,
61358	 => std_logic_vector(to_unsigned(25,8) ,
61359	 => std_logic_vector(to_unsigned(29,8) ,
61360	 => std_logic_vector(to_unsigned(20,8) ,
61361	 => std_logic_vector(to_unsigned(47,8) ,
61362	 => std_logic_vector(to_unsigned(50,8) ,
61363	 => std_logic_vector(to_unsigned(58,8) ,
61364	 => std_logic_vector(to_unsigned(69,8) ,
61365	 => std_logic_vector(to_unsigned(70,8) ,
61366	 => std_logic_vector(to_unsigned(73,8) ,
61367	 => std_logic_vector(to_unsigned(68,8) ,
61368	 => std_logic_vector(to_unsigned(62,8) ,
61369	 => std_logic_vector(to_unsigned(53,8) ,
61370	 => std_logic_vector(to_unsigned(30,8) ,
61371	 => std_logic_vector(to_unsigned(10,8) ,
61372	 => std_logic_vector(to_unsigned(12,8) ,
61373	 => std_logic_vector(to_unsigned(16,8) ,
61374	 => std_logic_vector(to_unsigned(13,8) ,
61375	 => std_logic_vector(to_unsigned(12,8) ,
61376	 => std_logic_vector(to_unsigned(12,8) ,
61377	 => std_logic_vector(to_unsigned(10,8) ,
61378	 => std_logic_vector(to_unsigned(14,8) ,
61379	 => std_logic_vector(to_unsigned(5,8) ,
61380	 => std_logic_vector(to_unsigned(10,8) ,
61381	 => std_logic_vector(to_unsigned(10,8) ,
61382	 => std_logic_vector(to_unsigned(11,8) ,
61383	 => std_logic_vector(to_unsigned(15,8) ,
61384	 => std_logic_vector(to_unsigned(12,8) ,
61385	 => std_logic_vector(to_unsigned(14,8) ,
61386	 => std_logic_vector(to_unsigned(8,8) ,
61387	 => std_logic_vector(to_unsigned(0,8) ,
61388	 => std_logic_vector(to_unsigned(0,8) ,
61389	 => std_logic_vector(to_unsigned(4,8) ,
61390	 => std_logic_vector(to_unsigned(10,8) ,
61391	 => std_logic_vector(to_unsigned(9,8) ,
61392	 => std_logic_vector(to_unsigned(8,8) ,
61393	 => std_logic_vector(to_unsigned(14,8) ,
61394	 => std_logic_vector(to_unsigned(24,8) ,
61395	 => std_logic_vector(to_unsigned(7,8) ,
61396	 => std_logic_vector(to_unsigned(8,8) ,
61397	 => std_logic_vector(to_unsigned(9,8) ,
61398	 => std_logic_vector(to_unsigned(9,8) ,
61399	 => std_logic_vector(to_unsigned(8,8) ,
61400	 => std_logic_vector(to_unsigned(8,8) ,
61401	 => std_logic_vector(to_unsigned(8,8) ,
61402	 => std_logic_vector(to_unsigned(4,8) ,
61403	 => std_logic_vector(to_unsigned(27,8) ,
61404	 => std_logic_vector(to_unsigned(16,8) ,
61405	 => std_logic_vector(to_unsigned(0,8) ,
61406	 => std_logic_vector(to_unsigned(1,8) ,
61407	 => std_logic_vector(to_unsigned(51,8) ,
61408	 => std_logic_vector(to_unsigned(22,8) ,
61409	 => std_logic_vector(to_unsigned(0,8) ,
61410	 => std_logic_vector(to_unsigned(0,8) ,
61411	 => std_logic_vector(to_unsigned(13,8) ,
61412	 => std_logic_vector(to_unsigned(38,8) ,
61413	 => std_logic_vector(to_unsigned(28,8) ,
61414	 => std_logic_vector(to_unsigned(14,8) ,
61415	 => std_logic_vector(to_unsigned(6,8) ,
61416	 => std_logic_vector(to_unsigned(6,8) ,
61417	 => std_logic_vector(to_unsigned(9,8) ,
61418	 => std_logic_vector(to_unsigned(9,8) ,
61419	 => std_logic_vector(to_unsigned(6,8) ,
61420	 => std_logic_vector(to_unsigned(18,8) ,
61421	 => std_logic_vector(to_unsigned(15,8) ,
61422	 => std_logic_vector(to_unsigned(15,8) ,
61423	 => std_logic_vector(to_unsigned(21,8) ,
61424	 => std_logic_vector(to_unsigned(9,8) ,
61425	 => std_logic_vector(to_unsigned(8,8) ,
61426	 => std_logic_vector(to_unsigned(9,8) ,
61427	 => std_logic_vector(to_unsigned(14,8) ,
61428	 => std_logic_vector(to_unsigned(13,8) ,
61429	 => std_logic_vector(to_unsigned(16,8) ,
61430	 => std_logic_vector(to_unsigned(13,8) ,
61431	 => std_logic_vector(to_unsigned(9,8) ,
61432	 => std_logic_vector(to_unsigned(7,8) ,
61433	 => std_logic_vector(to_unsigned(9,8) ,
61434	 => std_logic_vector(to_unsigned(12,8) ,
61435	 => std_logic_vector(to_unsigned(9,8) ,
61436	 => std_logic_vector(to_unsigned(9,8) ,
61437	 => std_logic_vector(to_unsigned(8,8) ,
61438	 => std_logic_vector(to_unsigned(7,8) ,
61439	 => std_logic_vector(to_unsigned(8,8) ,
61440	 => std_logic_vector(to_unsigned(16,8) ,
61441	 => std_logic_vector(to_unsigned(57,8) ,
61442	 => std_logic_vector(to_unsigned(88,8) ,
61443	 => std_logic_vector(to_unsigned(81,8) ,
61444	 => std_logic_vector(to_unsigned(61,8) ,
61445	 => std_logic_vector(to_unsigned(73,8) ,
61446	 => std_logic_vector(to_unsigned(44,8) ,
61447	 => std_logic_vector(to_unsigned(31,8) ,
61448	 => std_logic_vector(to_unsigned(52,8) ,
61449	 => std_logic_vector(to_unsigned(58,8) ,
61450	 => std_logic_vector(to_unsigned(49,8) ,
61451	 => std_logic_vector(to_unsigned(43,8) ,
61452	 => std_logic_vector(to_unsigned(31,8) ,
61453	 => std_logic_vector(to_unsigned(27,8) ,
61454	 => std_logic_vector(to_unsigned(25,8) ,
61455	 => std_logic_vector(to_unsigned(27,8) ,
61456	 => std_logic_vector(to_unsigned(20,8) ,
61457	 => std_logic_vector(to_unsigned(24,8) ,
61458	 => std_logic_vector(to_unsigned(29,8) ,
61459	 => std_logic_vector(to_unsigned(40,8) ,
61460	 => std_logic_vector(to_unsigned(43,8) ,
61461	 => std_logic_vector(to_unsigned(40,8) ,
61462	 => std_logic_vector(to_unsigned(40,8) ,
61463	 => std_logic_vector(to_unsigned(35,8) ,
61464	 => std_logic_vector(to_unsigned(22,8) ,
61465	 => std_logic_vector(to_unsigned(32,8) ,
61466	 => std_logic_vector(to_unsigned(49,8) ,
61467	 => std_logic_vector(to_unsigned(32,8) ,
61468	 => std_logic_vector(to_unsigned(35,8) ,
61469	 => std_logic_vector(to_unsigned(25,8) ,
61470	 => std_logic_vector(to_unsigned(38,8) ,
61471	 => std_logic_vector(to_unsigned(35,8) ,
61472	 => std_logic_vector(to_unsigned(27,8) ,
61473	 => std_logic_vector(to_unsigned(39,8) ,
61474	 => std_logic_vector(to_unsigned(48,8) ,
61475	 => std_logic_vector(to_unsigned(44,8) ,
61476	 => std_logic_vector(to_unsigned(60,8) ,
61477	 => std_logic_vector(to_unsigned(71,8) ,
61478	 => std_logic_vector(to_unsigned(41,8) ,
61479	 => std_logic_vector(to_unsigned(53,8) ,
61480	 => std_logic_vector(to_unsigned(74,8) ,
61481	 => std_logic_vector(to_unsigned(35,8) ,
61482	 => std_logic_vector(to_unsigned(49,8) ,
61483	 => std_logic_vector(to_unsigned(78,8) ,
61484	 => std_logic_vector(to_unsigned(76,8) ,
61485	 => std_logic_vector(to_unsigned(69,8) ,
61486	 => std_logic_vector(to_unsigned(64,8) ,
61487	 => std_logic_vector(to_unsigned(64,8) ,
61488	 => std_logic_vector(to_unsigned(53,8) ,
61489	 => std_logic_vector(to_unsigned(46,8) ,
61490	 => std_logic_vector(to_unsigned(41,8) ,
61491	 => std_logic_vector(to_unsigned(37,8) ,
61492	 => std_logic_vector(to_unsigned(32,8) ,
61493	 => std_logic_vector(to_unsigned(51,8) ,
61494	 => std_logic_vector(to_unsigned(50,8) ,
61495	 => std_logic_vector(to_unsigned(58,8) ,
61496	 => std_logic_vector(to_unsigned(68,8) ,
61497	 => std_logic_vector(to_unsigned(53,8) ,
61498	 => std_logic_vector(to_unsigned(51,8) ,
61499	 => std_logic_vector(to_unsigned(51,8) ,
61500	 => std_logic_vector(to_unsigned(45,8) ,
61501	 => std_logic_vector(to_unsigned(45,8) ,
61502	 => std_logic_vector(to_unsigned(50,8) ,
61503	 => std_logic_vector(to_unsigned(85,8) ,
61504	 => std_logic_vector(to_unsigned(104,8) ,
61505	 => std_logic_vector(to_unsigned(101,8) ,
61506	 => std_logic_vector(to_unsigned(74,8) ,
61507	 => std_logic_vector(to_unsigned(64,8) ,
61508	 => std_logic_vector(to_unsigned(93,8) ,
61509	 => std_logic_vector(to_unsigned(91,8) ,
61510	 => std_logic_vector(to_unsigned(100,8) ,
61511	 => std_logic_vector(to_unsigned(99,8) ,
61512	 => std_logic_vector(to_unsigned(73,8) ,
61513	 => std_logic_vector(to_unsigned(95,8) ,
61514	 => std_logic_vector(to_unsigned(134,8) ,
61515	 => std_logic_vector(to_unsigned(136,8) ,
61516	 => std_logic_vector(to_unsigned(118,8) ,
61517	 => std_logic_vector(to_unsigned(116,8) ,
61518	 => std_logic_vector(to_unsigned(127,8) ,
61519	 => std_logic_vector(to_unsigned(127,8) ,
61520	 => std_logic_vector(to_unsigned(128,8) ,
61521	 => std_logic_vector(to_unsigned(131,8) ,
61522	 => std_logic_vector(to_unsigned(118,8) ,
61523	 => std_logic_vector(to_unsigned(119,8) ,
61524	 => std_logic_vector(to_unsigned(116,8) ,
61525	 => std_logic_vector(to_unsigned(116,8) ,
61526	 => std_logic_vector(to_unsigned(116,8) ,
61527	 => std_logic_vector(to_unsigned(93,8) ,
61528	 => std_logic_vector(to_unsigned(64,8) ,
61529	 => std_logic_vector(to_unsigned(58,8) ,
61530	 => std_logic_vector(to_unsigned(45,8) ,
61531	 => std_logic_vector(to_unsigned(39,8) ,
61532	 => std_logic_vector(to_unsigned(34,8) ,
61533	 => std_logic_vector(to_unsigned(33,8) ,
61534	 => std_logic_vector(to_unsigned(36,8) ,
61535	 => std_logic_vector(to_unsigned(41,8) ,
61536	 => std_logic_vector(to_unsigned(45,8) ,
61537	 => std_logic_vector(to_unsigned(47,8) ,
61538	 => std_logic_vector(to_unsigned(58,8) ,
61539	 => std_logic_vector(to_unsigned(68,8) ,
61540	 => std_logic_vector(to_unsigned(77,8) ,
61541	 => std_logic_vector(to_unsigned(93,8) ,
61542	 => std_logic_vector(to_unsigned(90,8) ,
61543	 => std_logic_vector(to_unsigned(93,8) ,
61544	 => std_logic_vector(to_unsigned(80,8) ,
61545	 => std_logic_vector(to_unsigned(37,8) ,
61546	 => std_logic_vector(to_unsigned(17,8) ,
61547	 => std_logic_vector(to_unsigned(23,8) ,
61548	 => std_logic_vector(to_unsigned(30,8) ,
61549	 => std_logic_vector(to_unsigned(25,8) ,
61550	 => std_logic_vector(to_unsigned(40,8) ,
61551	 => std_logic_vector(to_unsigned(79,8) ,
61552	 => std_logic_vector(to_unsigned(76,8) ,
61553	 => std_logic_vector(to_unsigned(73,8) ,
61554	 => std_logic_vector(to_unsigned(77,8) ,
61555	 => std_logic_vector(to_unsigned(54,8) ,
61556	 => std_logic_vector(to_unsigned(84,8) ,
61557	 => std_logic_vector(to_unsigned(82,8) ,
61558	 => std_logic_vector(to_unsigned(50,8) ,
61559	 => std_logic_vector(to_unsigned(73,8) ,
61560	 => std_logic_vector(to_unsigned(76,8) ,
61561	 => std_logic_vector(to_unsigned(51,8) ,
61562	 => std_logic_vector(to_unsigned(44,8) ,
61563	 => std_logic_vector(to_unsigned(76,8) ,
61564	 => std_logic_vector(to_unsigned(66,8) ,
61565	 => std_logic_vector(to_unsigned(45,8) ,
61566	 => std_logic_vector(to_unsigned(35,8) ,
61567	 => std_logic_vector(to_unsigned(35,8) ,
61568	 => std_logic_vector(to_unsigned(37,8) ,
61569	 => std_logic_vector(to_unsigned(37,8) ,
61570	 => std_logic_vector(to_unsigned(53,8) ,
61571	 => std_logic_vector(to_unsigned(26,8) ,
61572	 => std_logic_vector(to_unsigned(23,8) ,
61573	 => std_logic_vector(to_unsigned(32,8) ,
61574	 => std_logic_vector(to_unsigned(41,8) ,
61575	 => std_logic_vector(to_unsigned(36,8) ,
61576	 => std_logic_vector(to_unsigned(27,8) ,
61577	 => std_logic_vector(to_unsigned(22,8) ,
61578	 => std_logic_vector(to_unsigned(21,8) ,
61579	 => std_logic_vector(to_unsigned(35,8) ,
61580	 => std_logic_vector(to_unsigned(40,8) ,
61581	 => std_logic_vector(to_unsigned(37,8) ,
61582	 => std_logic_vector(to_unsigned(26,8) ,
61583	 => std_logic_vector(to_unsigned(57,8) ,
61584	 => std_logic_vector(to_unsigned(60,8) ,
61585	 => std_logic_vector(to_unsigned(15,8) ,
61586	 => std_logic_vector(to_unsigned(41,8) ,
61587	 => std_logic_vector(to_unsigned(19,8) ,
61588	 => std_logic_vector(to_unsigned(38,8) ,
61589	 => std_logic_vector(to_unsigned(67,8) ,
61590	 => std_logic_vector(to_unsigned(54,8) ,
61591	 => std_logic_vector(to_unsigned(56,8) ,
61592	 => std_logic_vector(to_unsigned(60,8) ,
61593	 => std_logic_vector(to_unsigned(59,8) ,
61594	 => std_logic_vector(to_unsigned(57,8) ,
61595	 => std_logic_vector(to_unsigned(56,8) ,
61596	 => std_logic_vector(to_unsigned(70,8) ,
61597	 => std_logic_vector(to_unsigned(50,8) ,
61598	 => std_logic_vector(to_unsigned(37,8) ,
61599	 => std_logic_vector(to_unsigned(32,8) ,
61600	 => std_logic_vector(to_unsigned(32,8) ,
61601	 => std_logic_vector(to_unsigned(54,8) ,
61602	 => std_logic_vector(to_unsigned(60,8) ,
61603	 => std_logic_vector(to_unsigned(29,8) ,
61604	 => std_logic_vector(to_unsigned(5,8) ,
61605	 => std_logic_vector(to_unsigned(11,8) ,
61606	 => std_logic_vector(to_unsigned(7,8) ,
61607	 => std_logic_vector(to_unsigned(24,8) ,
61608	 => std_logic_vector(to_unsigned(64,8) ,
61609	 => std_logic_vector(to_unsigned(30,8) ,
61610	 => std_logic_vector(to_unsigned(4,8) ,
61611	 => std_logic_vector(to_unsigned(37,8) ,
61612	 => std_logic_vector(to_unsigned(52,8) ,
61613	 => std_logic_vector(to_unsigned(45,8) ,
61614	 => std_logic_vector(to_unsigned(26,8) ,
61615	 => std_logic_vector(to_unsigned(43,8) ,
61616	 => std_logic_vector(to_unsigned(57,8) ,
61617	 => std_logic_vector(to_unsigned(49,8) ,
61618	 => std_logic_vector(to_unsigned(57,8) ,
61619	 => std_logic_vector(to_unsigned(108,8) ,
61620	 => std_logic_vector(to_unsigned(66,8) ,
61621	 => std_logic_vector(to_unsigned(10,8) ,
61622	 => std_logic_vector(to_unsigned(8,8) ,
61623	 => std_logic_vector(to_unsigned(11,8) ,
61624	 => std_logic_vector(to_unsigned(12,8) ,
61625	 => std_logic_vector(to_unsigned(8,8) ,
61626	 => std_logic_vector(to_unsigned(19,8) ,
61627	 => std_logic_vector(to_unsigned(52,8) ,
61628	 => std_logic_vector(to_unsigned(12,8) ,
61629	 => std_logic_vector(to_unsigned(13,8) ,
61630	 => std_logic_vector(to_unsigned(39,8) ,
61631	 => std_logic_vector(to_unsigned(48,8) ,
61632	 => std_logic_vector(to_unsigned(41,8) ,
61633	 => std_logic_vector(to_unsigned(29,8) ,
61634	 => std_logic_vector(to_unsigned(22,8) ,
61635	 => std_logic_vector(to_unsigned(25,8) ,
61636	 => std_logic_vector(to_unsigned(35,8) ,
61637	 => std_logic_vector(to_unsigned(38,8) ,
61638	 => std_logic_vector(to_unsigned(49,8) ,
61639	 => std_logic_vector(to_unsigned(41,8) ,
61640	 => std_logic_vector(to_unsigned(28,8) ,
61641	 => std_logic_vector(to_unsigned(48,8) ,
61642	 => std_logic_vector(to_unsigned(66,8) ,
61643	 => std_logic_vector(to_unsigned(51,8) ,
61644	 => std_logic_vector(to_unsigned(35,8) ,
61645	 => std_logic_vector(to_unsigned(39,8) ,
61646	 => std_logic_vector(to_unsigned(64,8) ,
61647	 => std_logic_vector(to_unsigned(68,8) ,
61648	 => std_logic_vector(to_unsigned(57,8) ,
61649	 => std_logic_vector(to_unsigned(32,8) ,
61650	 => std_logic_vector(to_unsigned(24,8) ,
61651	 => std_logic_vector(to_unsigned(27,8) ,
61652	 => std_logic_vector(to_unsigned(37,8) ,
61653	 => std_logic_vector(to_unsigned(35,8) ,
61654	 => std_logic_vector(to_unsigned(34,8) ,
61655	 => std_logic_vector(to_unsigned(51,8) ,
61656	 => std_logic_vector(to_unsigned(81,8) ,
61657	 => std_logic_vector(to_unsigned(78,8) ,
61658	 => std_logic_vector(to_unsigned(54,8) ,
61659	 => std_logic_vector(to_unsigned(33,8) ,
61660	 => std_logic_vector(to_unsigned(41,8) ,
61661	 => std_logic_vector(to_unsigned(29,8) ,
61662	 => std_logic_vector(to_unsigned(17,8) ,
61663	 => std_logic_vector(to_unsigned(19,8) ,
61664	 => std_logic_vector(to_unsigned(31,8) ,
61665	 => std_logic_vector(to_unsigned(32,8) ,
61666	 => std_logic_vector(to_unsigned(35,8) ,
61667	 => std_logic_vector(to_unsigned(49,8) ,
61668	 => std_logic_vector(to_unsigned(37,8) ,
61669	 => std_logic_vector(to_unsigned(37,8) ,
61670	 => std_logic_vector(to_unsigned(43,8) ,
61671	 => std_logic_vector(to_unsigned(39,8) ,
61672	 => std_logic_vector(to_unsigned(35,8) ,
61673	 => std_logic_vector(to_unsigned(36,8) ,
61674	 => std_logic_vector(to_unsigned(32,8) ,
61675	 => std_logic_vector(to_unsigned(31,8) ,
61676	 => std_logic_vector(to_unsigned(29,8) ,
61677	 => std_logic_vector(to_unsigned(23,8) ,
61678	 => std_logic_vector(to_unsigned(23,8) ,
61679	 => std_logic_vector(to_unsigned(25,8) ,
61680	 => std_logic_vector(to_unsigned(17,8) ,
61681	 => std_logic_vector(to_unsigned(24,8) ,
61682	 => std_logic_vector(to_unsigned(17,8) ,
61683	 => std_logic_vector(to_unsigned(27,8) ,
61684	 => std_logic_vector(to_unsigned(35,8) ,
61685	 => std_logic_vector(to_unsigned(31,8) ,
61686	 => std_logic_vector(to_unsigned(45,8) ,
61687	 => std_logic_vector(to_unsigned(50,8) ,
61688	 => std_logic_vector(to_unsigned(42,8) ,
61689	 => std_logic_vector(to_unsigned(49,8) ,
61690	 => std_logic_vector(to_unsigned(41,8) ,
61691	 => std_logic_vector(to_unsigned(8,8) ,
61692	 => std_logic_vector(to_unsigned(9,8) ,
61693	 => std_logic_vector(to_unsigned(10,8) ,
61694	 => std_logic_vector(to_unsigned(9,8) ,
61695	 => std_logic_vector(to_unsigned(9,8) ,
61696	 => std_logic_vector(to_unsigned(9,8) ,
61697	 => std_logic_vector(to_unsigned(12,8) ,
61698	 => std_logic_vector(to_unsigned(14,8) ,
61699	 => std_logic_vector(to_unsigned(10,8) ,
61700	 => std_logic_vector(to_unsigned(9,8) ,
61701	 => std_logic_vector(to_unsigned(8,8) ,
61702	 => std_logic_vector(to_unsigned(11,8) ,
61703	 => std_logic_vector(to_unsigned(13,8) ,
61704	 => std_logic_vector(to_unsigned(9,8) ,
61705	 => std_logic_vector(to_unsigned(8,8) ,
61706	 => std_logic_vector(to_unsigned(9,8) ,
61707	 => std_logic_vector(to_unsigned(1,8) ,
61708	 => std_logic_vector(to_unsigned(0,8) ,
61709	 => std_logic_vector(to_unsigned(2,8) ,
61710	 => std_logic_vector(to_unsigned(12,8) ,
61711	 => std_logic_vector(to_unsigned(14,8) ,
61712	 => std_logic_vector(to_unsigned(12,8) ,
61713	 => std_logic_vector(to_unsigned(15,8) ,
61714	 => std_logic_vector(to_unsigned(13,8) ,
61715	 => std_logic_vector(to_unsigned(8,8) ,
61716	 => std_logic_vector(to_unsigned(10,8) ,
61717	 => std_logic_vector(to_unsigned(10,8) ,
61718	 => std_logic_vector(to_unsigned(9,8) ,
61719	 => std_logic_vector(to_unsigned(9,8) ,
61720	 => std_logic_vector(to_unsigned(7,8) ,
61721	 => std_logic_vector(to_unsigned(10,8) ,
61722	 => std_logic_vector(to_unsigned(5,8) ,
61723	 => std_logic_vector(to_unsigned(32,8) ,
61724	 => std_logic_vector(to_unsigned(16,8) ,
61725	 => std_logic_vector(to_unsigned(0,8) ,
61726	 => std_logic_vector(to_unsigned(1,8) ,
61727	 => std_logic_vector(to_unsigned(71,8) ,
61728	 => std_logic_vector(to_unsigned(71,8) ,
61729	 => std_logic_vector(to_unsigned(2,8) ,
61730	 => std_logic_vector(to_unsigned(0,8) ,
61731	 => std_logic_vector(to_unsigned(5,8) ,
61732	 => std_logic_vector(to_unsigned(68,8) ,
61733	 => std_logic_vector(to_unsigned(61,8) ,
61734	 => std_logic_vector(to_unsigned(15,8) ,
61735	 => std_logic_vector(to_unsigned(9,8) ,
61736	 => std_logic_vector(to_unsigned(11,8) ,
61737	 => std_logic_vector(to_unsigned(10,8) ,
61738	 => std_logic_vector(to_unsigned(9,8) ,
61739	 => std_logic_vector(to_unsigned(10,8) ,
61740	 => std_logic_vector(to_unsigned(9,8) ,
61741	 => std_logic_vector(to_unsigned(9,8) ,
61742	 => std_logic_vector(to_unsigned(15,8) ,
61743	 => std_logic_vector(to_unsigned(7,8) ,
61744	 => std_logic_vector(to_unsigned(9,8) ,
61745	 => std_logic_vector(to_unsigned(11,8) ,
61746	 => std_logic_vector(to_unsigned(9,8) ,
61747	 => std_logic_vector(to_unsigned(9,8) ,
61748	 => std_logic_vector(to_unsigned(9,8) ,
61749	 => std_logic_vector(to_unsigned(13,8) ,
61750	 => std_logic_vector(to_unsigned(21,8) ,
61751	 => std_logic_vector(to_unsigned(17,8) ,
61752	 => std_logic_vector(to_unsigned(17,8) ,
61753	 => std_logic_vector(to_unsigned(13,8) ,
61754	 => std_logic_vector(to_unsigned(13,8) ,
61755	 => std_logic_vector(to_unsigned(16,8) ,
61756	 => std_logic_vector(to_unsigned(9,8) ,
61757	 => std_logic_vector(to_unsigned(5,8) ,
61758	 => std_logic_vector(to_unsigned(7,8) ,
61759	 => std_logic_vector(to_unsigned(9,8) ,
61760	 => std_logic_vector(to_unsigned(11,8) ,
61761	 => std_logic_vector(to_unsigned(57,8) ,
61762	 => std_logic_vector(to_unsigned(84,8) ,
61763	 => std_logic_vector(to_unsigned(88,8) ,
61764	 => std_logic_vector(to_unsigned(61,8) ,
61765	 => std_logic_vector(to_unsigned(64,8) ,
61766	 => std_logic_vector(to_unsigned(46,8) ,
61767	 => std_logic_vector(to_unsigned(30,8) ,
61768	 => std_logic_vector(to_unsigned(39,8) ,
61769	 => std_logic_vector(to_unsigned(51,8) ,
61770	 => std_logic_vector(to_unsigned(38,8) ,
61771	 => std_logic_vector(to_unsigned(37,8) ,
61772	 => std_logic_vector(to_unsigned(30,8) ,
61773	 => std_logic_vector(to_unsigned(20,8) ,
61774	 => std_logic_vector(to_unsigned(22,8) ,
61775	 => std_logic_vector(to_unsigned(24,8) ,
61776	 => std_logic_vector(to_unsigned(24,8) ,
61777	 => std_logic_vector(to_unsigned(22,8) ,
61778	 => std_logic_vector(to_unsigned(24,8) ,
61779	 => std_logic_vector(to_unsigned(32,8) ,
61780	 => std_logic_vector(to_unsigned(37,8) ,
61781	 => std_logic_vector(to_unsigned(47,8) ,
61782	 => std_logic_vector(to_unsigned(47,8) ,
61783	 => std_logic_vector(to_unsigned(25,8) ,
61784	 => std_logic_vector(to_unsigned(20,8) ,
61785	 => std_logic_vector(to_unsigned(28,8) ,
61786	 => std_logic_vector(to_unsigned(27,8) ,
61787	 => std_logic_vector(to_unsigned(21,8) ,
61788	 => std_logic_vector(to_unsigned(31,8) ,
61789	 => std_logic_vector(to_unsigned(32,8) ,
61790	 => std_logic_vector(to_unsigned(37,8) ,
61791	 => std_logic_vector(to_unsigned(35,8) ,
61792	 => std_logic_vector(to_unsigned(30,8) ,
61793	 => std_logic_vector(to_unsigned(35,8) ,
61794	 => std_logic_vector(to_unsigned(33,8) ,
61795	 => std_logic_vector(to_unsigned(40,8) ,
61796	 => std_logic_vector(to_unsigned(30,8) ,
61797	 => std_logic_vector(to_unsigned(23,8) ,
61798	 => std_logic_vector(to_unsigned(35,8) ,
61799	 => std_logic_vector(to_unsigned(46,8) ,
61800	 => std_logic_vector(to_unsigned(51,8) ,
61801	 => std_logic_vector(to_unsigned(42,8) ,
61802	 => std_logic_vector(to_unsigned(46,8) ,
61803	 => std_logic_vector(to_unsigned(62,8) ,
61804	 => std_logic_vector(to_unsigned(81,8) ,
61805	 => std_logic_vector(to_unsigned(74,8) ,
61806	 => std_logic_vector(to_unsigned(45,8) ,
61807	 => std_logic_vector(to_unsigned(56,8) ,
61808	 => std_logic_vector(to_unsigned(54,8) ,
61809	 => std_logic_vector(to_unsigned(44,8) ,
61810	 => std_logic_vector(to_unsigned(41,8) ,
61811	 => std_logic_vector(to_unsigned(37,8) ,
61812	 => std_logic_vector(to_unsigned(32,8) ,
61813	 => std_logic_vector(to_unsigned(52,8) ,
61814	 => std_logic_vector(to_unsigned(61,8) ,
61815	 => std_logic_vector(to_unsigned(77,8) ,
61816	 => std_logic_vector(to_unsigned(68,8) ,
61817	 => std_logic_vector(to_unsigned(54,8) ,
61818	 => std_logic_vector(to_unsigned(48,8) ,
61819	 => std_logic_vector(to_unsigned(57,8) ,
61820	 => std_logic_vector(to_unsigned(55,8) ,
61821	 => std_logic_vector(to_unsigned(41,8) ,
61822	 => std_logic_vector(to_unsigned(56,8) ,
61823	 => std_logic_vector(to_unsigned(85,8) ,
61824	 => std_logic_vector(to_unsigned(73,8) ,
61825	 => std_logic_vector(to_unsigned(85,8) ,
61826	 => std_logic_vector(to_unsigned(84,8) ,
61827	 => std_logic_vector(to_unsigned(82,8) ,
61828	 => std_logic_vector(to_unsigned(91,8) ,
61829	 => std_logic_vector(to_unsigned(97,8) ,
61830	 => std_logic_vector(to_unsigned(103,8) ,
61831	 => std_logic_vector(to_unsigned(108,8) ,
61832	 => std_logic_vector(to_unsigned(81,8) ,
61833	 => std_logic_vector(to_unsigned(95,8) ,
61834	 => std_logic_vector(to_unsigned(139,8) ,
61835	 => std_logic_vector(to_unsigned(131,8) ,
61836	 => std_logic_vector(to_unsigned(122,8) ,
61837	 => std_logic_vector(to_unsigned(107,8) ,
61838	 => std_logic_vector(to_unsigned(124,8) ,
61839	 => std_logic_vector(to_unsigned(139,8) ,
61840	 => std_logic_vector(to_unsigned(121,8) ,
61841	 => std_logic_vector(to_unsigned(119,8) ,
61842	 => std_logic_vector(to_unsigned(122,8) ,
61843	 => std_logic_vector(to_unsigned(114,8) ,
61844	 => std_logic_vector(to_unsigned(111,8) ,
61845	 => std_logic_vector(to_unsigned(118,8) ,
61846	 => std_logic_vector(to_unsigned(67,8) ,
61847	 => std_logic_vector(to_unsigned(41,8) ,
61848	 => std_logic_vector(to_unsigned(101,8) ,
61849	 => std_logic_vector(to_unsigned(154,8) ,
61850	 => std_logic_vector(to_unsigned(146,8) ,
61851	 => std_logic_vector(to_unsigned(125,8) ,
61852	 => std_logic_vector(to_unsigned(99,8) ,
61853	 => std_logic_vector(to_unsigned(77,8) ,
61854	 => std_logic_vector(to_unsigned(63,8) ,
61855	 => std_logic_vector(to_unsigned(59,8) ,
61856	 => std_logic_vector(to_unsigned(51,8) ,
61857	 => std_logic_vector(to_unsigned(50,8) ,
61858	 => std_logic_vector(to_unsigned(58,8) ,
61859	 => std_logic_vector(to_unsigned(51,8) ,
61860	 => std_logic_vector(to_unsigned(59,8) ,
61861	 => std_logic_vector(to_unsigned(51,8) ,
61862	 => std_logic_vector(to_unsigned(55,8) ,
61863	 => std_logic_vector(to_unsigned(66,8) ,
61864	 => std_logic_vector(to_unsigned(49,8) ,
61865	 => std_logic_vector(to_unsigned(17,8) ,
61866	 => std_logic_vector(to_unsigned(12,8) ,
61867	 => std_logic_vector(to_unsigned(27,8) ,
61868	 => std_logic_vector(to_unsigned(29,8) ,
61869	 => std_logic_vector(to_unsigned(22,8) ,
61870	 => std_logic_vector(to_unsigned(49,8) ,
61871	 => std_logic_vector(to_unsigned(105,8) ,
61872	 => std_logic_vector(to_unsigned(90,8) ,
61873	 => std_logic_vector(to_unsigned(65,8) ,
61874	 => std_logic_vector(to_unsigned(45,8) ,
61875	 => std_logic_vector(to_unsigned(36,8) ,
61876	 => std_logic_vector(to_unsigned(80,8) ,
61877	 => std_logic_vector(to_unsigned(104,8) ,
61878	 => std_logic_vector(to_unsigned(70,8) ,
61879	 => std_logic_vector(to_unsigned(81,8) ,
61880	 => std_logic_vector(to_unsigned(84,8) ,
61881	 => std_logic_vector(to_unsigned(76,8) ,
61882	 => std_logic_vector(to_unsigned(77,8) ,
61883	 => std_logic_vector(to_unsigned(88,8) ,
61884	 => std_logic_vector(to_unsigned(71,8) ,
61885	 => std_logic_vector(to_unsigned(39,8) ,
61886	 => std_logic_vector(to_unsigned(52,8) ,
61887	 => std_logic_vector(to_unsigned(62,8) ,
61888	 => std_logic_vector(to_unsigned(38,8) ,
61889	 => std_logic_vector(to_unsigned(24,8) ,
61890	 => std_logic_vector(to_unsigned(30,8) ,
61891	 => std_logic_vector(to_unsigned(27,8) ,
61892	 => std_logic_vector(to_unsigned(24,8) ,
61893	 => std_logic_vector(to_unsigned(35,8) ,
61894	 => std_logic_vector(to_unsigned(35,8) ,
61895	 => std_logic_vector(to_unsigned(24,8) ,
61896	 => std_logic_vector(to_unsigned(23,8) ,
61897	 => std_logic_vector(to_unsigned(25,8) ,
61898	 => std_logic_vector(to_unsigned(32,8) ,
61899	 => std_logic_vector(to_unsigned(29,8) ,
61900	 => std_logic_vector(to_unsigned(25,8) ,
61901	 => std_logic_vector(to_unsigned(25,8) ,
61902	 => std_logic_vector(to_unsigned(22,8) ,
61903	 => std_logic_vector(to_unsigned(62,8) ,
61904	 => std_logic_vector(to_unsigned(63,8) ,
61905	 => std_logic_vector(to_unsigned(30,8) ,
61906	 => std_logic_vector(to_unsigned(49,8) ,
61907	 => std_logic_vector(to_unsigned(11,8) ,
61908	 => std_logic_vector(to_unsigned(33,8) ,
61909	 => std_logic_vector(to_unsigned(103,8) ,
61910	 => std_logic_vector(to_unsigned(93,8) ,
61911	 => std_logic_vector(to_unsigned(88,8) ,
61912	 => std_logic_vector(to_unsigned(76,8) ,
61913	 => std_logic_vector(to_unsigned(64,8) ,
61914	 => std_logic_vector(to_unsigned(55,8) ,
61915	 => std_logic_vector(to_unsigned(51,8) ,
61916	 => std_logic_vector(to_unsigned(45,8) ,
61917	 => std_logic_vector(to_unsigned(51,8) ,
61918	 => std_logic_vector(to_unsigned(35,8) ,
61919	 => std_logic_vector(to_unsigned(18,8) ,
61920	 => std_logic_vector(to_unsigned(13,8) ,
61921	 => std_logic_vector(to_unsigned(17,8) ,
61922	 => std_logic_vector(to_unsigned(13,8) ,
61923	 => std_logic_vector(to_unsigned(6,8) ,
61924	 => std_logic_vector(to_unsigned(10,8) ,
61925	 => std_logic_vector(to_unsigned(16,8) ,
61926	 => std_logic_vector(to_unsigned(19,8) ,
61927	 => std_logic_vector(to_unsigned(34,8) ,
61928	 => std_logic_vector(to_unsigned(43,8) ,
61929	 => std_logic_vector(to_unsigned(22,8) ,
61930	 => std_logic_vector(to_unsigned(7,8) ,
61931	 => std_logic_vector(to_unsigned(30,8) ,
61932	 => std_logic_vector(to_unsigned(37,8) ,
61933	 => std_logic_vector(to_unsigned(34,8) ,
61934	 => std_logic_vector(to_unsigned(46,8) ,
61935	 => std_logic_vector(to_unsigned(51,8) ,
61936	 => std_logic_vector(to_unsigned(45,8) ,
61937	 => std_logic_vector(to_unsigned(50,8) ,
61938	 => std_logic_vector(to_unsigned(101,8) ,
61939	 => std_logic_vector(to_unsigned(61,8) ,
61940	 => std_logic_vector(to_unsigned(22,8) ,
61941	 => std_logic_vector(to_unsigned(15,8) ,
61942	 => std_logic_vector(to_unsigned(8,8) ,
61943	 => std_logic_vector(to_unsigned(9,8) ,
61944	 => std_logic_vector(to_unsigned(15,8) ,
61945	 => std_logic_vector(to_unsigned(16,8) ,
61946	 => std_logic_vector(to_unsigned(20,8) ,
61947	 => std_logic_vector(to_unsigned(45,8) ,
61948	 => std_logic_vector(to_unsigned(52,8) ,
61949	 => std_logic_vector(to_unsigned(50,8) ,
61950	 => std_logic_vector(to_unsigned(74,8) ,
61951	 => std_logic_vector(to_unsigned(50,8) ,
61952	 => std_logic_vector(to_unsigned(36,8) ,
61953	 => std_logic_vector(to_unsigned(22,8) ,
61954	 => std_logic_vector(to_unsigned(13,8) ,
61955	 => std_logic_vector(to_unsigned(15,8) ,
61956	 => std_logic_vector(to_unsigned(65,8) ,
61957	 => std_logic_vector(to_unsigned(55,8) ,
61958	 => std_logic_vector(to_unsigned(40,8) ,
61959	 => std_logic_vector(to_unsigned(38,8) ,
61960	 => std_logic_vector(to_unsigned(17,8) ,
61961	 => std_logic_vector(to_unsigned(37,8) ,
61962	 => std_logic_vector(to_unsigned(37,8) ,
61963	 => std_logic_vector(to_unsigned(29,8) ,
61964	 => std_logic_vector(to_unsigned(28,8) ,
61965	 => std_logic_vector(to_unsigned(44,8) ,
61966	 => std_logic_vector(to_unsigned(60,8) ,
61967	 => std_logic_vector(to_unsigned(66,8) ,
61968	 => std_logic_vector(to_unsigned(58,8) ,
61969	 => std_logic_vector(to_unsigned(33,8) ,
61970	 => std_logic_vector(to_unsigned(29,8) ,
61971	 => std_logic_vector(to_unsigned(22,8) ,
61972	 => std_logic_vector(to_unsigned(29,8) ,
61973	 => std_logic_vector(to_unsigned(35,8) ,
61974	 => std_logic_vector(to_unsigned(37,8) ,
61975	 => std_logic_vector(to_unsigned(51,8) ,
61976	 => std_logic_vector(to_unsigned(77,8) ,
61977	 => std_logic_vector(to_unsigned(107,8) ,
61978	 => std_logic_vector(to_unsigned(71,8) ,
61979	 => std_logic_vector(to_unsigned(30,8) ,
61980	 => std_logic_vector(to_unsigned(41,8) ,
61981	 => std_logic_vector(to_unsigned(32,8) ,
61982	 => std_logic_vector(to_unsigned(12,8) ,
61983	 => std_logic_vector(to_unsigned(7,8) ,
61984	 => std_logic_vector(to_unsigned(17,8) ,
61985	 => std_logic_vector(to_unsigned(41,8) ,
61986	 => std_logic_vector(to_unsigned(54,8) ,
61987	 => std_logic_vector(to_unsigned(56,8) ,
61988	 => std_logic_vector(to_unsigned(30,8) ,
61989	 => std_logic_vector(to_unsigned(24,8) ,
61990	 => std_logic_vector(to_unsigned(32,8) ,
61991	 => std_logic_vector(to_unsigned(37,8) ,
61992	 => std_logic_vector(to_unsigned(35,8) ,
61993	 => std_logic_vector(to_unsigned(35,8) ,
61994	 => std_logic_vector(to_unsigned(35,8) ,
61995	 => std_logic_vector(to_unsigned(40,8) ,
61996	 => std_logic_vector(to_unsigned(30,8) ,
61997	 => std_logic_vector(to_unsigned(30,8) ,
61998	 => std_logic_vector(to_unsigned(41,8) ,
61999	 => std_logic_vector(to_unsigned(40,8) ,
62000	 => std_logic_vector(to_unsigned(36,8) ,
62001	 => std_logic_vector(to_unsigned(35,8) ,
62002	 => std_logic_vector(to_unsigned(30,8) ,
62003	 => std_logic_vector(to_unsigned(27,8) ,
62004	 => std_logic_vector(to_unsigned(29,8) ,
62005	 => std_logic_vector(to_unsigned(13,8) ,
62006	 => std_logic_vector(to_unsigned(21,8) ,
62007	 => std_logic_vector(to_unsigned(40,8) ,
62008	 => std_logic_vector(to_unsigned(32,8) ,
62009	 => std_logic_vector(to_unsigned(30,8) ,
62010	 => std_logic_vector(to_unsigned(29,8) ,
62011	 => std_logic_vector(to_unsigned(10,8) ,
62012	 => std_logic_vector(to_unsigned(11,8) ,
62013	 => std_logic_vector(to_unsigned(11,8) ,
62014	 => std_logic_vector(to_unsigned(9,8) ,
62015	 => std_logic_vector(to_unsigned(8,8) ,
62016	 => std_logic_vector(to_unsigned(8,8) ,
62017	 => std_logic_vector(to_unsigned(9,8) ,
62018	 => std_logic_vector(to_unsigned(12,8) ,
62019	 => std_logic_vector(to_unsigned(12,8) ,
62020	 => std_logic_vector(to_unsigned(13,8) ,
62021	 => std_logic_vector(to_unsigned(13,8) ,
62022	 => std_logic_vector(to_unsigned(13,8) ,
62023	 => std_logic_vector(to_unsigned(18,8) ,
62024	 => std_logic_vector(to_unsigned(13,8) ,
62025	 => std_logic_vector(to_unsigned(12,8) ,
62026	 => std_logic_vector(to_unsigned(18,8) ,
62027	 => std_logic_vector(to_unsigned(4,8) ,
62028	 => std_logic_vector(to_unsigned(0,8) ,
62029	 => std_logic_vector(to_unsigned(1,8) ,
62030	 => std_logic_vector(to_unsigned(11,8) ,
62031	 => std_logic_vector(to_unsigned(18,8) ,
62032	 => std_logic_vector(to_unsigned(9,8) ,
62033	 => std_logic_vector(to_unsigned(9,8) ,
62034	 => std_logic_vector(to_unsigned(9,8) ,
62035	 => std_logic_vector(to_unsigned(8,8) ,
62036	 => std_logic_vector(to_unsigned(9,8) ,
62037	 => std_logic_vector(to_unsigned(9,8) ,
62038	 => std_logic_vector(to_unsigned(8,8) ,
62039	 => std_logic_vector(to_unsigned(7,8) ,
62040	 => std_logic_vector(to_unsigned(4,8) ,
62041	 => std_logic_vector(to_unsigned(3,8) ,
62042	 => std_logic_vector(to_unsigned(3,8) ,
62043	 => std_logic_vector(to_unsigned(25,8) ,
62044	 => std_logic_vector(to_unsigned(10,8) ,
62045	 => std_logic_vector(to_unsigned(0,8) ,
62046	 => std_logic_vector(to_unsigned(1,8) ,
62047	 => std_logic_vector(to_unsigned(20,8) ,
62048	 => std_logic_vector(to_unsigned(25,8) ,
62049	 => std_logic_vector(to_unsigned(6,8) ,
62050	 => std_logic_vector(to_unsigned(0,8) ,
62051	 => std_logic_vector(to_unsigned(1,8) ,
62052	 => std_logic_vector(to_unsigned(41,8) ,
62053	 => std_logic_vector(to_unsigned(66,8) ,
62054	 => std_logic_vector(to_unsigned(10,8) ,
62055	 => std_logic_vector(to_unsigned(10,8) ,
62056	 => std_logic_vector(to_unsigned(12,8) ,
62057	 => std_logic_vector(to_unsigned(12,8) ,
62058	 => std_logic_vector(to_unsigned(11,8) ,
62059	 => std_logic_vector(to_unsigned(24,8) ,
62060	 => std_logic_vector(to_unsigned(15,8) ,
62061	 => std_logic_vector(to_unsigned(16,8) ,
62062	 => std_logic_vector(to_unsigned(22,8) ,
62063	 => std_logic_vector(to_unsigned(15,8) ,
62064	 => std_logic_vector(to_unsigned(12,8) ,
62065	 => std_logic_vector(to_unsigned(9,8) ,
62066	 => std_logic_vector(to_unsigned(6,8) ,
62067	 => std_logic_vector(to_unsigned(4,8) ,
62068	 => std_logic_vector(to_unsigned(4,8) ,
62069	 => std_logic_vector(to_unsigned(10,8) ,
62070	 => std_logic_vector(to_unsigned(10,8) ,
62071	 => std_logic_vector(to_unsigned(11,8) ,
62072	 => std_logic_vector(to_unsigned(13,8) ,
62073	 => std_logic_vector(to_unsigned(12,8) ,
62074	 => std_logic_vector(to_unsigned(11,8) ,
62075	 => std_logic_vector(to_unsigned(13,8) ,
62076	 => std_logic_vector(to_unsigned(6,8) ,
62077	 => std_logic_vector(to_unsigned(6,8) ,
62078	 => std_logic_vector(to_unsigned(14,8) ,
62079	 => std_logic_vector(to_unsigned(15,8) ,
62080	 => std_logic_vector(to_unsigned(11,8) ,
62081	 => std_logic_vector(to_unsigned(64,8) ,
62082	 => std_logic_vector(to_unsigned(88,8) ,
62083	 => std_logic_vector(to_unsigned(92,8) ,
62084	 => std_logic_vector(to_unsigned(58,8) ,
62085	 => std_logic_vector(to_unsigned(65,8) ,
62086	 => std_logic_vector(to_unsigned(52,8) ,
62087	 => std_logic_vector(to_unsigned(40,8) ,
62088	 => std_logic_vector(to_unsigned(37,8) ,
62089	 => std_logic_vector(to_unsigned(40,8) ,
62090	 => std_logic_vector(to_unsigned(51,8) ,
62091	 => std_logic_vector(to_unsigned(52,8) ,
62092	 => std_logic_vector(to_unsigned(35,8) ,
62093	 => std_logic_vector(to_unsigned(22,8) ,
62094	 => std_logic_vector(to_unsigned(25,8) ,
62095	 => std_logic_vector(to_unsigned(23,8) ,
62096	 => std_logic_vector(to_unsigned(25,8) ,
62097	 => std_logic_vector(to_unsigned(23,8) ,
62098	 => std_logic_vector(to_unsigned(20,8) ,
62099	 => std_logic_vector(to_unsigned(14,8) ,
62100	 => std_logic_vector(to_unsigned(20,8) ,
62101	 => std_logic_vector(to_unsigned(56,8) ,
62102	 => std_logic_vector(to_unsigned(51,8) ,
62103	 => std_logic_vector(to_unsigned(21,8) ,
62104	 => std_logic_vector(to_unsigned(17,8) ,
62105	 => std_logic_vector(to_unsigned(15,8) ,
62106	 => std_logic_vector(to_unsigned(16,8) ,
62107	 => std_logic_vector(to_unsigned(16,8) ,
62108	 => std_logic_vector(to_unsigned(29,8) ,
62109	 => std_logic_vector(to_unsigned(50,8) ,
62110	 => std_logic_vector(to_unsigned(44,8) ,
62111	 => std_logic_vector(to_unsigned(32,8) ,
62112	 => std_logic_vector(to_unsigned(32,8) ,
62113	 => std_logic_vector(to_unsigned(36,8) ,
62114	 => std_logic_vector(to_unsigned(40,8) ,
62115	 => std_logic_vector(to_unsigned(37,8) ,
62116	 => std_logic_vector(to_unsigned(29,8) ,
62117	 => std_logic_vector(to_unsigned(29,8) ,
62118	 => std_logic_vector(to_unsigned(33,8) ,
62119	 => std_logic_vector(to_unsigned(34,8) ,
62120	 => std_logic_vector(to_unsigned(29,8) ,
62121	 => std_logic_vector(to_unsigned(34,8) ,
62122	 => std_logic_vector(to_unsigned(34,8) ,
62123	 => std_logic_vector(to_unsigned(39,8) ,
62124	 => std_logic_vector(to_unsigned(56,8) ,
62125	 => std_logic_vector(to_unsigned(60,8) ,
62126	 => std_logic_vector(to_unsigned(56,8) ,
62127	 => std_logic_vector(to_unsigned(59,8) ,
62128	 => std_logic_vector(to_unsigned(53,8) ,
62129	 => std_logic_vector(to_unsigned(48,8) ,
62130	 => std_logic_vector(to_unsigned(48,8) ,
62131	 => std_logic_vector(to_unsigned(39,8) ,
62132	 => std_logic_vector(to_unsigned(32,8) ,
62133	 => std_logic_vector(to_unsigned(46,8) ,
62134	 => std_logic_vector(to_unsigned(58,8) ,
62135	 => std_logic_vector(to_unsigned(72,8) ,
62136	 => std_logic_vector(to_unsigned(69,8) ,
62137	 => std_logic_vector(to_unsigned(54,8) ,
62138	 => std_logic_vector(to_unsigned(55,8) ,
62139	 => std_logic_vector(to_unsigned(58,8) ,
62140	 => std_logic_vector(to_unsigned(54,8) ,
62141	 => std_logic_vector(to_unsigned(51,8) ,
62142	 => std_logic_vector(to_unsigned(68,8) ,
62143	 => std_logic_vector(to_unsigned(90,8) ,
62144	 => std_logic_vector(to_unsigned(57,8) ,
62145	 => std_logic_vector(to_unsigned(80,8) ,
62146	 => std_logic_vector(to_unsigned(88,8) ,
62147	 => std_logic_vector(to_unsigned(67,8) ,
62148	 => std_logic_vector(to_unsigned(91,8) ,
62149	 => std_logic_vector(to_unsigned(76,8) ,
62150	 => std_logic_vector(to_unsigned(88,8) ,
62151	 => std_logic_vector(to_unsigned(103,8) ,
62152	 => std_logic_vector(to_unsigned(101,8) ,
62153	 => std_logic_vector(to_unsigned(111,8) ,
62154	 => std_logic_vector(to_unsigned(136,8) ,
62155	 => std_logic_vector(to_unsigned(119,8) ,
62156	 => std_logic_vector(to_unsigned(108,8) ,
62157	 => std_logic_vector(to_unsigned(136,8) ,
62158	 => std_logic_vector(to_unsigned(138,8) ,
62159	 => std_logic_vector(to_unsigned(127,8) ,
62160	 => std_logic_vector(to_unsigned(121,8) ,
62161	 => std_logic_vector(to_unsigned(119,8) ,
62162	 => std_logic_vector(to_unsigned(99,8) ,
62163	 => std_logic_vector(to_unsigned(73,8) ,
62164	 => std_logic_vector(to_unsigned(74,8) ,
62165	 => std_logic_vector(to_unsigned(88,8) ,
62166	 => std_logic_vector(to_unsigned(59,8) ,
62167	 => std_logic_vector(to_unsigned(41,8) ,
62168	 => std_logic_vector(to_unsigned(74,8) ,
62169	 => std_logic_vector(to_unsigned(105,8) ,
62170	 => std_logic_vector(to_unsigned(111,8) ,
62171	 => std_logic_vector(to_unsigned(134,8) ,
62172	 => std_logic_vector(to_unsigned(151,8) ,
62173	 => std_logic_vector(to_unsigned(144,8) ,
62174	 => std_logic_vector(to_unsigned(127,8) ,
62175	 => std_logic_vector(to_unsigned(125,8) ,
62176	 => std_logic_vector(to_unsigned(86,8) ,
62177	 => std_logic_vector(to_unsigned(74,8) ,
62178	 => std_logic_vector(to_unsigned(66,8) ,
62179	 => std_logic_vector(to_unsigned(54,8) ,
62180	 => std_logic_vector(to_unsigned(49,8) ,
62181	 => std_logic_vector(to_unsigned(38,8) ,
62182	 => std_logic_vector(to_unsigned(36,8) ,
62183	 => std_logic_vector(to_unsigned(41,8) ,
62184	 => std_logic_vector(to_unsigned(35,8) ,
62185	 => std_logic_vector(to_unsigned(42,8) ,
62186	 => std_logic_vector(to_unsigned(71,8) ,
62187	 => std_logic_vector(to_unsigned(68,8) ,
62188	 => std_logic_vector(to_unsigned(67,8) ,
62189	 => std_logic_vector(to_unsigned(71,8) ,
62190	 => std_logic_vector(to_unsigned(77,8) ,
62191	 => std_logic_vector(to_unsigned(70,8) ,
62192	 => std_logic_vector(to_unsigned(52,8) ,
62193	 => std_logic_vector(to_unsigned(68,8) ,
62194	 => std_logic_vector(to_unsigned(57,8) ,
62195	 => std_logic_vector(to_unsigned(45,8) ,
62196	 => std_logic_vector(to_unsigned(87,8) ,
62197	 => std_logic_vector(to_unsigned(81,8) ,
62198	 => std_logic_vector(to_unsigned(63,8) ,
62199	 => std_logic_vector(to_unsigned(87,8) ,
62200	 => std_logic_vector(to_unsigned(77,8) ,
62201	 => std_logic_vector(to_unsigned(87,8) ,
62202	 => std_logic_vector(to_unsigned(64,8) ,
62203	 => std_logic_vector(to_unsigned(53,8) ,
62204	 => std_logic_vector(to_unsigned(60,8) ,
62205	 => std_logic_vector(to_unsigned(49,8) ,
62206	 => std_logic_vector(to_unsigned(63,8) ,
62207	 => std_logic_vector(to_unsigned(81,8) ,
62208	 => std_logic_vector(to_unsigned(52,8) ,
62209	 => std_logic_vector(to_unsigned(45,8) ,
62210	 => std_logic_vector(to_unsigned(33,8) ,
62211	 => std_logic_vector(to_unsigned(19,8) ,
62212	 => std_logic_vector(to_unsigned(30,8) ,
62213	 => std_logic_vector(to_unsigned(37,8) ,
62214	 => std_logic_vector(to_unsigned(30,8) ,
62215	 => std_logic_vector(to_unsigned(28,8) ,
62216	 => std_logic_vector(to_unsigned(25,8) ,
62217	 => std_logic_vector(to_unsigned(30,8) ,
62218	 => std_logic_vector(to_unsigned(24,8) ,
62219	 => std_logic_vector(to_unsigned(18,8) ,
62220	 => std_logic_vector(to_unsigned(23,8) ,
62221	 => std_logic_vector(to_unsigned(17,8) ,
62222	 => std_logic_vector(to_unsigned(10,8) ,
62223	 => std_logic_vector(to_unsigned(42,8) ,
62224	 => std_logic_vector(to_unsigned(61,8) ,
62225	 => std_logic_vector(to_unsigned(41,8) ,
62226	 => std_logic_vector(to_unsigned(54,8) ,
62227	 => std_logic_vector(to_unsigned(32,8) ,
62228	 => std_logic_vector(to_unsigned(55,8) ,
62229	 => std_logic_vector(to_unsigned(93,8) ,
62230	 => std_logic_vector(to_unsigned(77,8) ,
62231	 => std_logic_vector(to_unsigned(84,8) ,
62232	 => std_logic_vector(to_unsigned(97,8) ,
62233	 => std_logic_vector(to_unsigned(90,8) ,
62234	 => std_logic_vector(to_unsigned(85,8) ,
62235	 => std_logic_vector(to_unsigned(85,8) ,
62236	 => std_logic_vector(to_unsigned(65,8) ,
62237	 => std_logic_vector(to_unsigned(38,8) ,
62238	 => std_logic_vector(to_unsigned(29,8) ,
62239	 => std_logic_vector(to_unsigned(23,8) ,
62240	 => std_logic_vector(to_unsigned(24,8) ,
62241	 => std_logic_vector(to_unsigned(13,8) ,
62242	 => std_logic_vector(to_unsigned(5,8) ,
62243	 => std_logic_vector(to_unsigned(17,8) ,
62244	 => std_logic_vector(to_unsigned(27,8) ,
62245	 => std_logic_vector(to_unsigned(30,8) ,
62246	 => std_logic_vector(to_unsigned(32,8) ,
62247	 => std_logic_vector(to_unsigned(41,8) ,
62248	 => std_logic_vector(to_unsigned(27,8) ,
62249	 => std_logic_vector(to_unsigned(14,8) ,
62250	 => std_logic_vector(to_unsigned(18,8) ,
62251	 => std_logic_vector(to_unsigned(27,8) ,
62252	 => std_logic_vector(to_unsigned(35,8) ,
62253	 => std_logic_vector(to_unsigned(45,8) ,
62254	 => std_logic_vector(to_unsigned(47,8) ,
62255	 => std_logic_vector(to_unsigned(43,8) ,
62256	 => std_logic_vector(to_unsigned(48,8) ,
62257	 => std_logic_vector(to_unsigned(104,8) ,
62258	 => std_logic_vector(to_unsigned(61,8) ,
62259	 => std_logic_vector(to_unsigned(17,8) ,
62260	 => std_logic_vector(to_unsigned(34,8) ,
62261	 => std_logic_vector(to_unsigned(22,8) ,
62262	 => std_logic_vector(to_unsigned(9,8) ,
62263	 => std_logic_vector(to_unsigned(12,8) ,
62264	 => std_logic_vector(to_unsigned(14,8) ,
62265	 => std_logic_vector(to_unsigned(17,8) ,
62266	 => std_logic_vector(to_unsigned(19,8) ,
62267	 => std_logic_vector(to_unsigned(43,8) ,
62268	 => std_logic_vector(to_unsigned(53,8) ,
62269	 => std_logic_vector(to_unsigned(41,8) ,
62270	 => std_logic_vector(to_unsigned(51,8) ,
62271	 => std_logic_vector(to_unsigned(45,8) ,
62272	 => std_logic_vector(to_unsigned(29,8) ,
62273	 => std_logic_vector(to_unsigned(25,8) ,
62274	 => std_logic_vector(to_unsigned(20,8) ,
62275	 => std_logic_vector(to_unsigned(19,8) ,
62276	 => std_logic_vector(to_unsigned(76,8) ,
62277	 => std_logic_vector(to_unsigned(66,8) ,
62278	 => std_logic_vector(to_unsigned(45,8) ,
62279	 => std_logic_vector(to_unsigned(40,8) ,
62280	 => std_logic_vector(to_unsigned(30,8) ,
62281	 => std_logic_vector(to_unsigned(60,8) ,
62282	 => std_logic_vector(to_unsigned(35,8) ,
62283	 => std_logic_vector(to_unsigned(21,8) ,
62284	 => std_logic_vector(to_unsigned(30,8) ,
62285	 => std_logic_vector(to_unsigned(42,8) ,
62286	 => std_logic_vector(to_unsigned(41,8) ,
62287	 => std_logic_vector(to_unsigned(44,8) ,
62288	 => std_logic_vector(to_unsigned(42,8) ,
62289	 => std_logic_vector(to_unsigned(41,8) ,
62290	 => std_logic_vector(to_unsigned(23,8) ,
62291	 => std_logic_vector(to_unsigned(11,8) ,
62292	 => std_logic_vector(to_unsigned(19,8) ,
62293	 => std_logic_vector(to_unsigned(39,8) ,
62294	 => std_logic_vector(to_unsigned(46,8) ,
62295	 => std_logic_vector(to_unsigned(47,8) ,
62296	 => std_logic_vector(to_unsigned(51,8) ,
62297	 => std_logic_vector(to_unsigned(60,8) ,
62298	 => std_logic_vector(to_unsigned(50,8) ,
62299	 => std_logic_vector(to_unsigned(37,8) ,
62300	 => std_logic_vector(to_unsigned(36,8) ,
62301	 => std_logic_vector(to_unsigned(34,8) ,
62302	 => std_logic_vector(to_unsigned(24,8) ,
62303	 => std_logic_vector(to_unsigned(22,8) ,
62304	 => std_logic_vector(to_unsigned(27,8) ,
62305	 => std_logic_vector(to_unsigned(50,8) ,
62306	 => std_logic_vector(to_unsigned(68,8) ,
62307	 => std_logic_vector(to_unsigned(47,8) ,
62308	 => std_logic_vector(to_unsigned(36,8) ,
62309	 => std_logic_vector(to_unsigned(32,8) ,
62310	 => std_logic_vector(to_unsigned(30,8) ,
62311	 => std_logic_vector(to_unsigned(29,8) ,
62312	 => std_logic_vector(to_unsigned(28,8) ,
62313	 => std_logic_vector(to_unsigned(26,8) ,
62314	 => std_logic_vector(to_unsigned(30,8) ,
62315	 => std_logic_vector(to_unsigned(32,8) ,
62316	 => std_logic_vector(to_unsigned(17,8) ,
62317	 => std_logic_vector(to_unsigned(23,8) ,
62318	 => std_logic_vector(to_unsigned(27,8) ,
62319	 => std_logic_vector(to_unsigned(28,8) ,
62320	 => std_logic_vector(to_unsigned(41,8) ,
62321	 => std_logic_vector(to_unsigned(44,8) ,
62322	 => std_logic_vector(to_unsigned(39,8) ,
62323	 => std_logic_vector(to_unsigned(32,8) ,
62324	 => std_logic_vector(to_unsigned(28,8) ,
62325	 => std_logic_vector(to_unsigned(22,8) ,
62326	 => std_logic_vector(to_unsigned(29,8) ,
62327	 => std_logic_vector(to_unsigned(35,8) ,
62328	 => std_logic_vector(to_unsigned(34,8) ,
62329	 => std_logic_vector(to_unsigned(32,8) ,
62330	 => std_logic_vector(to_unsigned(30,8) ,
62331	 => std_logic_vector(to_unsigned(27,8) ,
62332	 => std_logic_vector(to_unsigned(19,8) ,
62333	 => std_logic_vector(to_unsigned(13,8) ,
62334	 => std_logic_vector(to_unsigned(12,8) ,
62335	 => std_logic_vector(to_unsigned(8,8) ,
62336	 => std_logic_vector(to_unsigned(9,8) ,
62337	 => std_logic_vector(to_unsigned(10,8) ,
62338	 => std_logic_vector(to_unsigned(11,8) ,
62339	 => std_logic_vector(to_unsigned(8,8) ,
62340	 => std_logic_vector(to_unsigned(11,8) ,
62341	 => std_logic_vector(to_unsigned(12,8) ,
62342	 => std_logic_vector(to_unsigned(11,8) ,
62343	 => std_logic_vector(to_unsigned(13,8) ,
62344	 => std_logic_vector(to_unsigned(12,8) ,
62345	 => std_logic_vector(to_unsigned(12,8) ,
62346	 => std_logic_vector(to_unsigned(15,8) ,
62347	 => std_logic_vector(to_unsigned(9,8) ,
62348	 => std_logic_vector(to_unsigned(1,8) ,
62349	 => std_logic_vector(to_unsigned(0,8) ,
62350	 => std_logic_vector(to_unsigned(4,8) ,
62351	 => std_logic_vector(to_unsigned(14,8) ,
62352	 => std_logic_vector(to_unsigned(10,8) ,
62353	 => std_logic_vector(to_unsigned(9,8) ,
62354	 => std_logic_vector(to_unsigned(8,8) ,
62355	 => std_logic_vector(to_unsigned(12,8) ,
62356	 => std_logic_vector(to_unsigned(10,8) ,
62357	 => std_logic_vector(to_unsigned(6,8) ,
62358	 => std_logic_vector(to_unsigned(6,8) ,
62359	 => std_logic_vector(to_unsigned(6,8) ,
62360	 => std_logic_vector(to_unsigned(6,8) ,
62361	 => std_logic_vector(to_unsigned(5,8) ,
62362	 => std_logic_vector(to_unsigned(3,8) ,
62363	 => std_logic_vector(to_unsigned(32,8) ,
62364	 => std_logic_vector(to_unsigned(18,8) ,
62365	 => std_logic_vector(to_unsigned(0,8) ,
62366	 => std_logic_vector(to_unsigned(1,8) ,
62367	 => std_logic_vector(to_unsigned(9,8) ,
62368	 => std_logic_vector(to_unsigned(17,8) ,
62369	 => std_logic_vector(to_unsigned(22,8) ,
62370	 => std_logic_vector(to_unsigned(2,8) ,
62371	 => std_logic_vector(to_unsigned(0,8) ,
62372	 => std_logic_vector(to_unsigned(8,8) ,
62373	 => std_logic_vector(to_unsigned(45,8) ,
62374	 => std_logic_vector(to_unsigned(14,8) ,
62375	 => std_logic_vector(to_unsigned(12,8) ,
62376	 => std_logic_vector(to_unsigned(12,8) ,
62377	 => std_logic_vector(to_unsigned(12,8) ,
62378	 => std_logic_vector(to_unsigned(12,8) ,
62379	 => std_logic_vector(to_unsigned(27,8) ,
62380	 => std_logic_vector(to_unsigned(25,8) ,
62381	 => std_logic_vector(to_unsigned(33,8) ,
62382	 => std_logic_vector(to_unsigned(35,8) ,
62383	 => std_logic_vector(to_unsigned(35,8) ,
62384	 => std_logic_vector(to_unsigned(18,8) ,
62385	 => std_logic_vector(to_unsigned(13,8) ,
62386	 => std_logic_vector(to_unsigned(16,8) ,
62387	 => std_logic_vector(to_unsigned(8,8) ,
62388	 => std_logic_vector(to_unsigned(8,8) ,
62389	 => std_logic_vector(to_unsigned(16,8) ,
62390	 => std_logic_vector(to_unsigned(17,8) ,
62391	 => std_logic_vector(to_unsigned(16,8) ,
62392	 => std_logic_vector(to_unsigned(11,8) ,
62393	 => std_logic_vector(to_unsigned(12,8) ,
62394	 => std_logic_vector(to_unsigned(18,8) ,
62395	 => std_logic_vector(to_unsigned(16,8) ,
62396	 => std_logic_vector(to_unsigned(12,8) ,
62397	 => std_logic_vector(to_unsigned(15,8) ,
62398	 => std_logic_vector(to_unsigned(14,8) ,
62399	 => std_logic_vector(to_unsigned(9,8) ,
62400	 => std_logic_vector(to_unsigned(9,8) ,
62401	 => std_logic_vector(to_unsigned(51,8) ,
62402	 => std_logic_vector(to_unsigned(77,8) ,
62403	 => std_logic_vector(to_unsigned(88,8) ,
62404	 => std_logic_vector(to_unsigned(54,8) ,
62405	 => std_logic_vector(to_unsigned(62,8) ,
62406	 => std_logic_vector(to_unsigned(55,8) ,
62407	 => std_logic_vector(to_unsigned(48,8) ,
62408	 => std_logic_vector(to_unsigned(57,8) ,
62409	 => std_logic_vector(to_unsigned(60,8) ,
62410	 => std_logic_vector(to_unsigned(56,8) ,
62411	 => std_logic_vector(to_unsigned(52,8) ,
62412	 => std_logic_vector(to_unsigned(41,8) ,
62413	 => std_logic_vector(to_unsigned(27,8) ,
62414	 => std_logic_vector(to_unsigned(29,8) ,
62415	 => std_logic_vector(to_unsigned(27,8) ,
62416	 => std_logic_vector(to_unsigned(35,8) ,
62417	 => std_logic_vector(to_unsigned(40,8) ,
62418	 => std_logic_vector(to_unsigned(29,8) ,
62419	 => std_logic_vector(to_unsigned(31,8) ,
62420	 => std_logic_vector(to_unsigned(46,8) ,
62421	 => std_logic_vector(to_unsigned(60,8) ,
62422	 => std_logic_vector(to_unsigned(49,8) ,
62423	 => std_logic_vector(to_unsigned(22,8) ,
62424	 => std_logic_vector(to_unsigned(15,8) ,
62425	 => std_logic_vector(to_unsigned(16,8) ,
62426	 => std_logic_vector(to_unsigned(24,8) ,
62427	 => std_logic_vector(to_unsigned(24,8) ,
62428	 => std_logic_vector(to_unsigned(27,8) ,
62429	 => std_logic_vector(to_unsigned(51,8) ,
62430	 => std_logic_vector(to_unsigned(46,8) ,
62431	 => std_logic_vector(to_unsigned(27,8) ,
62432	 => std_logic_vector(to_unsigned(30,8) ,
62433	 => std_logic_vector(to_unsigned(36,8) ,
62434	 => std_logic_vector(to_unsigned(40,8) ,
62435	 => std_logic_vector(to_unsigned(32,8) ,
62436	 => std_logic_vector(to_unsigned(32,8) ,
62437	 => std_logic_vector(to_unsigned(37,8) ,
62438	 => std_logic_vector(to_unsigned(30,8) ,
62439	 => std_logic_vector(to_unsigned(35,8) ,
62440	 => std_logic_vector(to_unsigned(36,8) ,
62441	 => std_logic_vector(to_unsigned(32,8) ,
62442	 => std_logic_vector(to_unsigned(35,8) ,
62443	 => std_logic_vector(to_unsigned(42,8) ,
62444	 => std_logic_vector(to_unsigned(49,8) ,
62445	 => std_logic_vector(to_unsigned(51,8) ,
62446	 => std_logic_vector(to_unsigned(64,8) ,
62447	 => std_logic_vector(to_unsigned(61,8) ,
62448	 => std_logic_vector(to_unsigned(59,8) ,
62449	 => std_logic_vector(to_unsigned(54,8) ,
62450	 => std_logic_vector(to_unsigned(47,8) ,
62451	 => std_logic_vector(to_unsigned(36,8) ,
62452	 => std_logic_vector(to_unsigned(29,8) ,
62453	 => std_logic_vector(to_unsigned(43,8) ,
62454	 => std_logic_vector(to_unsigned(56,8) ,
62455	 => std_logic_vector(to_unsigned(80,8) ,
62456	 => std_logic_vector(to_unsigned(91,8) ,
62457	 => std_logic_vector(to_unsigned(55,8) ,
62458	 => std_logic_vector(to_unsigned(54,8) ,
62459	 => std_logic_vector(to_unsigned(67,8) ,
62460	 => std_logic_vector(to_unsigned(70,8) ,
62461	 => std_logic_vector(to_unsigned(58,8) ,
62462	 => std_logic_vector(to_unsigned(58,8) ,
62463	 => std_logic_vector(to_unsigned(86,8) ,
62464	 => std_logic_vector(to_unsigned(85,8) ,
62465	 => std_logic_vector(to_unsigned(87,8) ,
62466	 => std_logic_vector(to_unsigned(84,8) ,
62467	 => std_logic_vector(to_unsigned(82,8) ,
62468	 => std_logic_vector(to_unsigned(93,8) ,
62469	 => std_logic_vector(to_unsigned(73,8) ,
62470	 => std_logic_vector(to_unsigned(88,8) ,
62471	 => std_logic_vector(to_unsigned(93,8) ,
62472	 => std_logic_vector(to_unsigned(72,8) ,
62473	 => std_logic_vector(to_unsigned(95,8) ,
62474	 => std_logic_vector(to_unsigned(124,8) ,
62475	 => std_logic_vector(to_unsigned(121,8) ,
62476	 => std_logic_vector(to_unsigned(125,8) ,
62477	 => std_logic_vector(to_unsigned(125,8) ,
62478	 => std_logic_vector(to_unsigned(124,8) ,
62479	 => std_logic_vector(to_unsigned(130,8) ,
62480	 => std_logic_vector(to_unsigned(127,8) ,
62481	 => std_logic_vector(to_unsigned(107,8) ,
62482	 => std_logic_vector(to_unsigned(58,8) ,
62483	 => std_logic_vector(to_unsigned(54,8) ,
62484	 => std_logic_vector(to_unsigned(81,8) ,
62485	 => std_logic_vector(to_unsigned(92,8) ,
62486	 => std_logic_vector(to_unsigned(88,8) ,
62487	 => std_logic_vector(to_unsigned(90,8) ,
62488	 => std_logic_vector(to_unsigned(95,8) ,
62489	 => std_logic_vector(to_unsigned(79,8) ,
62490	 => std_logic_vector(to_unsigned(67,8) ,
62491	 => std_logic_vector(to_unsigned(66,8) ,
62492	 => std_logic_vector(to_unsigned(71,8) ,
62493	 => std_logic_vector(to_unsigned(87,8) ,
62494	 => std_logic_vector(to_unsigned(82,8) ,
62495	 => std_logic_vector(to_unsigned(79,8) ,
62496	 => std_logic_vector(to_unsigned(58,8) ,
62497	 => std_logic_vector(to_unsigned(64,8) ,
62498	 => std_logic_vector(to_unsigned(63,8) ,
62499	 => std_logic_vector(to_unsigned(59,8) ,
62500	 => std_logic_vector(to_unsigned(49,8) ,
62501	 => std_logic_vector(to_unsigned(38,8) ,
62502	 => std_logic_vector(to_unsigned(39,8) ,
62503	 => std_logic_vector(to_unsigned(45,8) ,
62504	 => std_logic_vector(to_unsigned(46,8) ,
62505	 => std_logic_vector(to_unsigned(68,8) ,
62506	 => std_logic_vector(to_unsigned(56,8) ,
62507	 => std_logic_vector(to_unsigned(35,8) ,
62508	 => std_logic_vector(to_unsigned(52,8) ,
62509	 => std_logic_vector(to_unsigned(51,8) ,
62510	 => std_logic_vector(to_unsigned(49,8) ,
62511	 => std_logic_vector(to_unsigned(51,8) ,
62512	 => std_logic_vector(to_unsigned(44,8) ,
62513	 => std_logic_vector(to_unsigned(48,8) ,
62514	 => std_logic_vector(to_unsigned(56,8) ,
62515	 => std_logic_vector(to_unsigned(60,8) ,
62516	 => std_logic_vector(to_unsigned(80,8) ,
62517	 => std_logic_vector(to_unsigned(79,8) ,
62518	 => std_logic_vector(to_unsigned(71,8) ,
62519	 => std_logic_vector(to_unsigned(87,8) ,
62520	 => std_logic_vector(to_unsigned(63,8) ,
62521	 => std_logic_vector(to_unsigned(108,8) ,
62522	 => std_logic_vector(to_unsigned(77,8) ,
62523	 => std_logic_vector(to_unsigned(30,8) ,
62524	 => std_logic_vector(to_unsigned(30,8) ,
62525	 => std_logic_vector(to_unsigned(43,8) ,
62526	 => std_logic_vector(to_unsigned(60,8) ,
62527	 => std_logic_vector(to_unsigned(73,8) ,
62528	 => std_logic_vector(to_unsigned(52,8) ,
62529	 => std_logic_vector(to_unsigned(39,8) ,
62530	 => std_logic_vector(to_unsigned(23,8) ,
62531	 => std_logic_vector(to_unsigned(13,8) ,
62532	 => std_logic_vector(to_unsigned(16,8) ,
62533	 => std_logic_vector(to_unsigned(32,8) ,
62534	 => std_logic_vector(to_unsigned(52,8) ,
62535	 => std_logic_vector(to_unsigned(45,8) ,
62536	 => std_logic_vector(to_unsigned(37,8) ,
62537	 => std_logic_vector(to_unsigned(47,8) ,
62538	 => std_logic_vector(to_unsigned(38,8) ,
62539	 => std_logic_vector(to_unsigned(32,8) ,
62540	 => std_logic_vector(to_unsigned(32,8) ,
62541	 => std_logic_vector(to_unsigned(14,8) ,
62542	 => std_logic_vector(to_unsigned(5,8) ,
62543	 => std_logic_vector(to_unsigned(25,8) ,
62544	 => std_logic_vector(to_unsigned(45,8) ,
62545	 => std_logic_vector(to_unsigned(37,8) ,
62546	 => std_logic_vector(to_unsigned(50,8) ,
62547	 => std_logic_vector(to_unsigned(28,8) ,
62548	 => std_logic_vector(to_unsigned(53,8) ,
62549	 => std_logic_vector(to_unsigned(96,8) ,
62550	 => std_logic_vector(to_unsigned(65,8) ,
62551	 => std_logic_vector(to_unsigned(61,8) ,
62552	 => std_logic_vector(to_unsigned(87,8) ,
62553	 => std_logic_vector(to_unsigned(59,8) ,
62554	 => std_logic_vector(to_unsigned(66,8) ,
62555	 => std_logic_vector(to_unsigned(87,8) ,
62556	 => std_logic_vector(to_unsigned(60,8) ,
62557	 => std_logic_vector(to_unsigned(27,8) ,
62558	 => std_logic_vector(to_unsigned(24,8) ,
62559	 => std_logic_vector(to_unsigned(22,8) ,
62560	 => std_logic_vector(to_unsigned(22,8) ,
62561	 => std_logic_vector(to_unsigned(13,8) ,
62562	 => std_logic_vector(to_unsigned(9,8) ,
62563	 => std_logic_vector(to_unsigned(25,8) ,
62564	 => std_logic_vector(to_unsigned(35,8) ,
62565	 => std_logic_vector(to_unsigned(14,8) ,
62566	 => std_logic_vector(to_unsigned(10,8) ,
62567	 => std_logic_vector(to_unsigned(34,8) ,
62568	 => std_logic_vector(to_unsigned(30,8) ,
62569	 => std_logic_vector(to_unsigned(8,8) ,
62570	 => std_logic_vector(to_unsigned(15,8) ,
62571	 => std_logic_vector(to_unsigned(42,8) ,
62572	 => std_logic_vector(to_unsigned(50,8) ,
62573	 => std_logic_vector(to_unsigned(45,8) ,
62574	 => std_logic_vector(to_unsigned(43,8) ,
62575	 => std_logic_vector(to_unsigned(50,8) ,
62576	 => std_logic_vector(to_unsigned(96,8) ,
62577	 => std_logic_vector(to_unsigned(50,8) ,
62578	 => std_logic_vector(to_unsigned(17,8) ,
62579	 => std_logic_vector(to_unsigned(41,8) ,
62580	 => std_logic_vector(to_unsigned(32,8) ,
62581	 => std_logic_vector(to_unsigned(8,8) ,
62582	 => std_logic_vector(to_unsigned(9,8) ,
62583	 => std_logic_vector(to_unsigned(13,8) ,
62584	 => std_logic_vector(to_unsigned(12,8) ,
62585	 => std_logic_vector(to_unsigned(17,8) ,
62586	 => std_logic_vector(to_unsigned(28,8) ,
62587	 => std_logic_vector(to_unsigned(59,8) ,
62588	 => std_logic_vector(to_unsigned(46,8) ,
62589	 => std_logic_vector(to_unsigned(36,8) ,
62590	 => std_logic_vector(to_unsigned(36,8) ,
62591	 => std_logic_vector(to_unsigned(43,8) ,
62592	 => std_logic_vector(to_unsigned(41,8) ,
62593	 => std_logic_vector(to_unsigned(47,8) ,
62594	 => std_logic_vector(to_unsigned(50,8) ,
62595	 => std_logic_vector(to_unsigned(50,8) ,
62596	 => std_logic_vector(to_unsigned(65,8) ,
62597	 => std_logic_vector(to_unsigned(51,8) ,
62598	 => std_logic_vector(to_unsigned(45,8) ,
62599	 => std_logic_vector(to_unsigned(52,8) ,
62600	 => std_logic_vector(to_unsigned(53,8) ,
62601	 => std_logic_vector(to_unsigned(57,8) ,
62602	 => std_logic_vector(to_unsigned(35,8) ,
62603	 => std_logic_vector(to_unsigned(25,8) ,
62604	 => std_logic_vector(to_unsigned(45,8) ,
62605	 => std_logic_vector(to_unsigned(53,8) ,
62606	 => std_logic_vector(to_unsigned(48,8) ,
62607	 => std_logic_vector(to_unsigned(37,8) ,
62608	 => std_logic_vector(to_unsigned(45,8) ,
62609	 => std_logic_vector(to_unsigned(65,8) ,
62610	 => std_logic_vector(to_unsigned(14,8) ,
62611	 => std_logic_vector(to_unsigned(7,8) ,
62612	 => std_logic_vector(to_unsigned(15,8) ,
62613	 => std_logic_vector(to_unsigned(47,8) ,
62614	 => std_logic_vector(to_unsigned(76,8) ,
62615	 => std_logic_vector(to_unsigned(72,8) ,
62616	 => std_logic_vector(to_unsigned(64,8) ,
62617	 => std_logic_vector(to_unsigned(51,8) ,
62618	 => std_logic_vector(to_unsigned(53,8) ,
62619	 => std_logic_vector(to_unsigned(46,8) ,
62620	 => std_logic_vector(to_unsigned(32,8) ,
62621	 => std_logic_vector(to_unsigned(29,8) ,
62622	 => std_logic_vector(to_unsigned(32,8) ,
62623	 => std_logic_vector(to_unsigned(29,8) ,
62624	 => std_logic_vector(to_unsigned(32,8) ,
62625	 => std_logic_vector(to_unsigned(36,8) ,
62626	 => std_logic_vector(to_unsigned(39,8) ,
62627	 => std_logic_vector(to_unsigned(41,8) ,
62628	 => std_logic_vector(to_unsigned(44,8) ,
62629	 => std_logic_vector(to_unsigned(35,8) ,
62630	 => std_logic_vector(to_unsigned(37,8) ,
62631	 => std_logic_vector(to_unsigned(31,8) ,
62632	 => std_logic_vector(to_unsigned(31,8) ,
62633	 => std_logic_vector(to_unsigned(32,8) ,
62634	 => std_logic_vector(to_unsigned(29,8) ,
62635	 => std_logic_vector(to_unsigned(31,8) ,
62636	 => std_logic_vector(to_unsigned(32,8) ,
62637	 => std_logic_vector(to_unsigned(32,8) ,
62638	 => std_logic_vector(to_unsigned(13,8) ,
62639	 => std_logic_vector(to_unsigned(18,8) ,
62640	 => std_logic_vector(to_unsigned(35,8) ,
62641	 => std_logic_vector(to_unsigned(35,8) ,
62642	 => std_logic_vector(to_unsigned(32,8) ,
62643	 => std_logic_vector(to_unsigned(31,8) ,
62644	 => std_logic_vector(to_unsigned(30,8) ,
62645	 => std_logic_vector(to_unsigned(35,8) ,
62646	 => std_logic_vector(to_unsigned(39,8) ,
62647	 => std_logic_vector(to_unsigned(30,8) ,
62648	 => std_logic_vector(to_unsigned(30,8) ,
62649	 => std_logic_vector(to_unsigned(32,8) ,
62650	 => std_logic_vector(to_unsigned(35,8) ,
62651	 => std_logic_vector(to_unsigned(17,8) ,
62652	 => std_logic_vector(to_unsigned(12,8) ,
62653	 => std_logic_vector(to_unsigned(12,8) ,
62654	 => std_logic_vector(to_unsigned(9,8) ,
62655	 => std_logic_vector(to_unsigned(7,8) ,
62656	 => std_logic_vector(to_unsigned(7,8) ,
62657	 => std_logic_vector(to_unsigned(9,8) ,
62658	 => std_logic_vector(to_unsigned(9,8) ,
62659	 => std_logic_vector(to_unsigned(10,8) ,
62660	 => std_logic_vector(to_unsigned(11,8) ,
62661	 => std_logic_vector(to_unsigned(12,8) ,
62662	 => std_logic_vector(to_unsigned(10,8) ,
62663	 => std_logic_vector(to_unsigned(10,8) ,
62664	 => std_logic_vector(to_unsigned(9,8) ,
62665	 => std_logic_vector(to_unsigned(9,8) ,
62666	 => std_logic_vector(to_unsigned(8,8) ,
62667	 => std_logic_vector(to_unsigned(10,8) ,
62668	 => std_logic_vector(to_unsigned(3,8) ,
62669	 => std_logic_vector(to_unsigned(0,8) ,
62670	 => std_logic_vector(to_unsigned(1,8) ,
62671	 => std_logic_vector(to_unsigned(5,8) ,
62672	 => std_logic_vector(to_unsigned(9,8) ,
62673	 => std_logic_vector(to_unsigned(10,8) ,
62674	 => std_logic_vector(to_unsigned(9,8) ,
62675	 => std_logic_vector(to_unsigned(11,8) ,
62676	 => std_logic_vector(to_unsigned(12,8) ,
62677	 => std_logic_vector(to_unsigned(8,8) ,
62678	 => std_logic_vector(to_unsigned(6,8) ,
62679	 => std_logic_vector(to_unsigned(6,8) ,
62680	 => std_logic_vector(to_unsigned(5,8) ,
62681	 => std_logic_vector(to_unsigned(7,8) ,
62682	 => std_logic_vector(to_unsigned(5,8) ,
62683	 => std_logic_vector(to_unsigned(27,8) ,
62684	 => std_logic_vector(to_unsigned(11,8) ,
62685	 => std_logic_vector(to_unsigned(0,8) ,
62686	 => std_logic_vector(to_unsigned(0,8) ,
62687	 => std_logic_vector(to_unsigned(6,8) ,
62688	 => std_logic_vector(to_unsigned(65,8) ,
62689	 => std_logic_vector(to_unsigned(80,8) ,
62690	 => std_logic_vector(to_unsigned(13,8) ,
62691	 => std_logic_vector(to_unsigned(0,8) ,
62692	 => std_logic_vector(to_unsigned(1,8) ,
62693	 => std_logic_vector(to_unsigned(23,8) ,
62694	 => std_logic_vector(to_unsigned(18,8) ,
62695	 => std_logic_vector(to_unsigned(13,8) ,
62696	 => std_logic_vector(to_unsigned(17,8) ,
62697	 => std_logic_vector(to_unsigned(13,8) ,
62698	 => std_logic_vector(to_unsigned(17,8) ,
62699	 => std_logic_vector(to_unsigned(29,8) ,
62700	 => std_logic_vector(to_unsigned(18,8) ,
62701	 => std_logic_vector(to_unsigned(18,8) ,
62702	 => std_logic_vector(to_unsigned(22,8) ,
62703	 => std_logic_vector(to_unsigned(20,8) ,
62704	 => std_logic_vector(to_unsigned(17,8) ,
62705	 => std_logic_vector(to_unsigned(20,8) ,
62706	 => std_logic_vector(to_unsigned(35,8) ,
62707	 => std_logic_vector(to_unsigned(35,8) ,
62708	 => std_logic_vector(to_unsigned(32,8) ,
62709	 => std_logic_vector(to_unsigned(33,8) ,
62710	 => std_logic_vector(to_unsigned(27,8) ,
62711	 => std_logic_vector(to_unsigned(20,8) ,
62712	 => std_logic_vector(to_unsigned(20,8) ,
62713	 => std_logic_vector(to_unsigned(23,8) ,
62714	 => std_logic_vector(to_unsigned(20,8) ,
62715	 => std_logic_vector(to_unsigned(15,8) ,
62716	 => std_logic_vector(to_unsigned(20,8) ,
62717	 => std_logic_vector(to_unsigned(22,8) ,
62718	 => std_logic_vector(to_unsigned(14,8) ,
62719	 => std_logic_vector(to_unsigned(11,8) ,
62720	 => std_logic_vector(to_unsigned(12,8) ,
62721	 => std_logic_vector(to_unsigned(49,8) ,
62722	 => std_logic_vector(to_unsigned(67,8) ,
62723	 => std_logic_vector(to_unsigned(87,8) ,
62724	 => std_logic_vector(to_unsigned(60,8) ,
62725	 => std_logic_vector(to_unsigned(55,8) ,
62726	 => std_logic_vector(to_unsigned(65,8) ,
62727	 => std_logic_vector(to_unsigned(77,8) ,
62728	 => std_logic_vector(to_unsigned(72,8) ,
62729	 => std_logic_vector(to_unsigned(65,8) ,
62730	 => std_logic_vector(to_unsigned(59,8) ,
62731	 => std_logic_vector(to_unsigned(57,8) ,
62732	 => std_logic_vector(to_unsigned(51,8) ,
62733	 => std_logic_vector(to_unsigned(47,8) ,
62734	 => std_logic_vector(to_unsigned(45,8) ,
62735	 => std_logic_vector(to_unsigned(45,8) ,
62736	 => std_logic_vector(to_unsigned(53,8) ,
62737	 => std_logic_vector(to_unsigned(56,8) ,
62738	 => std_logic_vector(to_unsigned(55,8) ,
62739	 => std_logic_vector(to_unsigned(58,8) ,
62740	 => std_logic_vector(to_unsigned(57,8) ,
62741	 => std_logic_vector(to_unsigned(48,8) ,
62742	 => std_logic_vector(to_unsigned(47,8) ,
62743	 => std_logic_vector(to_unsigned(22,8) ,
62744	 => std_logic_vector(to_unsigned(18,8) ,
62745	 => std_logic_vector(to_unsigned(22,8) ,
62746	 => std_logic_vector(to_unsigned(22,8) ,
62747	 => std_logic_vector(to_unsigned(17,8) ,
62748	 => std_logic_vector(to_unsigned(22,8) ,
62749	 => std_logic_vector(to_unsigned(37,8) ,
62750	 => std_logic_vector(to_unsigned(33,8) ,
62751	 => std_logic_vector(to_unsigned(32,8) ,
62752	 => std_logic_vector(to_unsigned(45,8) ,
62753	 => std_logic_vector(to_unsigned(39,8) ,
62754	 => std_logic_vector(to_unsigned(34,8) ,
62755	 => std_logic_vector(to_unsigned(30,8) ,
62756	 => std_logic_vector(to_unsigned(32,8) ,
62757	 => std_logic_vector(to_unsigned(27,8) ,
62758	 => std_logic_vector(to_unsigned(23,8) ,
62759	 => std_logic_vector(to_unsigned(29,8) ,
62760	 => std_logic_vector(to_unsigned(41,8) ,
62761	 => std_logic_vector(to_unsigned(36,8) ,
62762	 => std_logic_vector(to_unsigned(35,8) ,
62763	 => std_logic_vector(to_unsigned(41,8) ,
62764	 => std_logic_vector(to_unsigned(55,8) ,
62765	 => std_logic_vector(to_unsigned(63,8) ,
62766	 => std_logic_vector(to_unsigned(62,8) ,
62767	 => std_logic_vector(to_unsigned(64,8) ,
62768	 => std_logic_vector(to_unsigned(63,8) ,
62769	 => std_logic_vector(to_unsigned(52,8) ,
62770	 => std_logic_vector(to_unsigned(40,8) ,
62771	 => std_logic_vector(to_unsigned(32,8) ,
62772	 => std_logic_vector(to_unsigned(28,8) ,
62773	 => std_logic_vector(to_unsigned(44,8) ,
62774	 => std_logic_vector(to_unsigned(59,8) ,
62775	 => std_logic_vector(to_unsigned(76,8) ,
62776	 => std_logic_vector(to_unsigned(80,8) ,
62777	 => std_logic_vector(to_unsigned(56,8) ,
62778	 => std_logic_vector(to_unsigned(54,8) ,
62779	 => std_logic_vector(to_unsigned(55,8) ,
62780	 => std_logic_vector(to_unsigned(50,8) ,
62781	 => std_logic_vector(to_unsigned(45,8) ,
62782	 => std_logic_vector(to_unsigned(53,8) ,
62783	 => std_logic_vector(to_unsigned(81,8) ,
62784	 => std_logic_vector(to_unsigned(78,8) ,
62785	 => std_logic_vector(to_unsigned(88,8) ,
62786	 => std_logic_vector(to_unsigned(85,8) ,
62787	 => std_logic_vector(to_unsigned(84,8) ,
62788	 => std_logic_vector(to_unsigned(90,8) ,
62789	 => std_logic_vector(to_unsigned(93,8) ,
62790	 => std_logic_vector(to_unsigned(90,8) ,
62791	 => std_logic_vector(to_unsigned(92,8) ,
62792	 => std_logic_vector(to_unsigned(84,8) ,
62793	 => std_logic_vector(to_unsigned(95,8) ,
62794	 => std_logic_vector(to_unsigned(136,8) ,
62795	 => std_logic_vector(to_unsigned(118,8) ,
62796	 => std_logic_vector(to_unsigned(109,8) ,
62797	 => std_logic_vector(to_unsigned(114,8) ,
62798	 => std_logic_vector(to_unsigned(124,8) ,
62799	 => std_logic_vector(to_unsigned(128,8) ,
62800	 => std_logic_vector(to_unsigned(121,8) ,
62801	 => std_logic_vector(to_unsigned(93,8) ,
62802	 => std_logic_vector(to_unsigned(59,8) ,
62803	 => std_logic_vector(to_unsigned(59,8) ,
62804	 => std_logic_vector(to_unsigned(79,8) ,
62805	 => std_logic_vector(to_unsigned(104,8) ,
62806	 => std_logic_vector(to_unsigned(86,8) ,
62807	 => std_logic_vector(to_unsigned(71,8) ,
62808	 => std_logic_vector(to_unsigned(82,8) ,
62809	 => std_logic_vector(to_unsigned(95,8) ,
62810	 => std_logic_vector(to_unsigned(87,8) ,
62811	 => std_logic_vector(to_unsigned(64,8) ,
62812	 => std_logic_vector(to_unsigned(64,8) ,
62813	 => std_logic_vector(to_unsigned(69,8) ,
62814	 => std_logic_vector(to_unsigned(35,8) ,
62815	 => std_logic_vector(to_unsigned(35,8) ,
62816	 => std_logic_vector(to_unsigned(40,8) ,
62817	 => std_logic_vector(to_unsigned(41,8) ,
62818	 => std_logic_vector(to_unsigned(53,8) ,
62819	 => std_logic_vector(to_unsigned(53,8) ,
62820	 => std_logic_vector(to_unsigned(59,8) ,
62821	 => std_logic_vector(to_unsigned(57,8) ,
62822	 => std_logic_vector(to_unsigned(41,8) ,
62823	 => std_logic_vector(to_unsigned(24,8) ,
62824	 => std_logic_vector(to_unsigned(29,8) ,
62825	 => std_logic_vector(to_unsigned(50,8) ,
62826	 => std_logic_vector(to_unsigned(45,8) ,
62827	 => std_logic_vector(to_unsigned(25,8) ,
62828	 => std_logic_vector(to_unsigned(51,8) ,
62829	 => std_logic_vector(to_unsigned(56,8) ,
62830	 => std_logic_vector(to_unsigned(39,8) ,
62831	 => std_logic_vector(to_unsigned(51,8) ,
62832	 => std_logic_vector(to_unsigned(46,8) ,
62833	 => std_logic_vector(to_unsigned(37,8) ,
62834	 => std_logic_vector(to_unsigned(38,8) ,
62835	 => std_logic_vector(to_unsigned(44,8) ,
62836	 => std_logic_vector(to_unsigned(64,8) ,
62837	 => std_logic_vector(to_unsigned(88,8) ,
62838	 => std_logic_vector(to_unsigned(88,8) ,
62839	 => std_logic_vector(to_unsigned(99,8) ,
62840	 => std_logic_vector(to_unsigned(48,8) ,
62841	 => std_logic_vector(to_unsigned(105,8) ,
62842	 => std_logic_vector(to_unsigned(111,8) ,
62843	 => std_logic_vector(to_unsigned(35,8) ,
62844	 => std_logic_vector(to_unsigned(30,8) ,
62845	 => std_logic_vector(to_unsigned(29,8) ,
62846	 => std_logic_vector(to_unsigned(41,8) ,
62847	 => std_logic_vector(to_unsigned(51,8) ,
62848	 => std_logic_vector(to_unsigned(26,8) ,
62849	 => std_logic_vector(to_unsigned(30,8) ,
62850	 => std_logic_vector(to_unsigned(45,8) ,
62851	 => std_logic_vector(to_unsigned(38,8) ,
62852	 => std_logic_vector(to_unsigned(27,8) ,
62853	 => std_logic_vector(to_unsigned(31,8) ,
62854	 => std_logic_vector(to_unsigned(58,8) ,
62855	 => std_logic_vector(to_unsigned(52,8) ,
62856	 => std_logic_vector(to_unsigned(47,8) ,
62857	 => std_logic_vector(to_unsigned(50,8) ,
62858	 => std_logic_vector(to_unsigned(56,8) ,
62859	 => std_logic_vector(to_unsigned(56,8) ,
62860	 => std_logic_vector(to_unsigned(43,8) ,
62861	 => std_logic_vector(to_unsigned(27,8) ,
62862	 => std_logic_vector(to_unsigned(22,8) ,
62863	 => std_logic_vector(to_unsigned(29,8) ,
62864	 => std_logic_vector(to_unsigned(23,8) ,
62865	 => std_logic_vector(to_unsigned(24,8) ,
62866	 => std_logic_vector(to_unsigned(24,8) ,
62867	 => std_logic_vector(to_unsigned(26,8) ,
62868	 => std_logic_vector(to_unsigned(58,8) ,
62869	 => std_logic_vector(to_unsigned(91,8) ,
62870	 => std_logic_vector(to_unsigned(80,8) ,
62871	 => std_logic_vector(to_unsigned(78,8) ,
62872	 => std_logic_vector(to_unsigned(84,8) ,
62873	 => std_logic_vector(to_unsigned(61,8) ,
62874	 => std_logic_vector(to_unsigned(67,8) ,
62875	 => std_logic_vector(to_unsigned(82,8) ,
62876	 => std_logic_vector(to_unsigned(55,8) ,
62877	 => std_logic_vector(to_unsigned(28,8) ,
62878	 => std_logic_vector(to_unsigned(19,8) ,
62879	 => std_logic_vector(to_unsigned(11,8) ,
62880	 => std_logic_vector(to_unsigned(29,8) ,
62881	 => std_logic_vector(to_unsigned(64,8) ,
62882	 => std_logic_vector(to_unsigned(44,8) ,
62883	 => std_logic_vector(to_unsigned(27,8) ,
62884	 => std_logic_vector(to_unsigned(31,8) ,
62885	 => std_logic_vector(to_unsigned(20,8) ,
62886	 => std_logic_vector(to_unsigned(12,8) ,
62887	 => std_logic_vector(to_unsigned(28,8) ,
62888	 => std_logic_vector(to_unsigned(41,8) ,
62889	 => std_logic_vector(to_unsigned(12,8) ,
62890	 => std_logic_vector(to_unsigned(22,8) ,
62891	 => std_logic_vector(to_unsigned(40,8) ,
62892	 => std_logic_vector(to_unsigned(43,8) ,
62893	 => std_logic_vector(to_unsigned(39,8) ,
62894	 => std_logic_vector(to_unsigned(44,8) ,
62895	 => std_logic_vector(to_unsigned(96,8) ,
62896	 => std_logic_vector(to_unsigned(59,8) ,
62897	 => std_logic_vector(to_unsigned(17,8) ,
62898	 => std_logic_vector(to_unsigned(33,8) ,
62899	 => std_logic_vector(to_unsigned(33,8) ,
62900	 => std_logic_vector(to_unsigned(20,8) ,
62901	 => std_logic_vector(to_unsigned(10,8) ,
62902	 => std_logic_vector(to_unsigned(8,8) ,
62903	 => std_logic_vector(to_unsigned(12,8) ,
62904	 => std_logic_vector(to_unsigned(10,8) ,
62905	 => std_logic_vector(to_unsigned(12,8) ,
62906	 => std_logic_vector(to_unsigned(56,8) ,
62907	 => std_logic_vector(to_unsigned(58,8) ,
62908	 => std_logic_vector(to_unsigned(35,8) ,
62909	 => std_logic_vector(to_unsigned(37,8) ,
62910	 => std_logic_vector(to_unsigned(46,8) ,
62911	 => std_logic_vector(to_unsigned(47,8) ,
62912	 => std_logic_vector(to_unsigned(47,8) ,
62913	 => std_logic_vector(to_unsigned(42,8) ,
62914	 => std_logic_vector(to_unsigned(46,8) ,
62915	 => std_logic_vector(to_unsigned(50,8) ,
62916	 => std_logic_vector(to_unsigned(53,8) ,
62917	 => std_logic_vector(to_unsigned(44,8) ,
62918	 => std_logic_vector(to_unsigned(45,8) ,
62919	 => std_logic_vector(to_unsigned(56,8) ,
62920	 => std_logic_vector(to_unsigned(49,8) ,
62921	 => std_logic_vector(to_unsigned(38,8) ,
62922	 => std_logic_vector(to_unsigned(26,8) ,
62923	 => std_logic_vector(to_unsigned(25,8) ,
62924	 => std_logic_vector(to_unsigned(43,8) ,
62925	 => std_logic_vector(to_unsigned(51,8) ,
62926	 => std_logic_vector(to_unsigned(51,8) ,
62927	 => std_logic_vector(to_unsigned(35,8) ,
62928	 => std_logic_vector(to_unsigned(30,8) ,
62929	 => std_logic_vector(to_unsigned(50,8) ,
62930	 => std_logic_vector(to_unsigned(29,8) ,
62931	 => std_logic_vector(to_unsigned(16,8) ,
62932	 => std_logic_vector(to_unsigned(26,8) ,
62933	 => std_logic_vector(to_unsigned(61,8) ,
62934	 => std_logic_vector(to_unsigned(71,8) ,
62935	 => std_logic_vector(to_unsigned(73,8) ,
62936	 => std_logic_vector(to_unsigned(85,8) ,
62937	 => std_logic_vector(to_unsigned(84,8) ,
62938	 => std_logic_vector(to_unsigned(85,8) ,
62939	 => std_logic_vector(to_unsigned(51,8) ,
62940	 => std_logic_vector(to_unsigned(20,8) ,
62941	 => std_logic_vector(to_unsigned(32,8) ,
62942	 => std_logic_vector(to_unsigned(61,8) ,
62943	 => std_logic_vector(to_unsigned(56,8) ,
62944	 => std_logic_vector(to_unsigned(41,8) ,
62945	 => std_logic_vector(to_unsigned(35,8) ,
62946	 => std_logic_vector(to_unsigned(35,8) ,
62947	 => std_logic_vector(to_unsigned(40,8) ,
62948	 => std_logic_vector(to_unsigned(41,8) ,
62949	 => std_logic_vector(to_unsigned(28,8) ,
62950	 => std_logic_vector(to_unsigned(22,8) ,
62951	 => std_logic_vector(to_unsigned(28,8) ,
62952	 => std_logic_vector(to_unsigned(22,8) ,
62953	 => std_logic_vector(to_unsigned(30,8) ,
62954	 => std_logic_vector(to_unsigned(41,8) ,
62955	 => std_logic_vector(to_unsigned(40,8) ,
62956	 => std_logic_vector(to_unsigned(45,8) ,
62957	 => std_logic_vector(to_unsigned(38,8) ,
62958	 => std_logic_vector(to_unsigned(35,8) ,
62959	 => std_logic_vector(to_unsigned(39,8) ,
62960	 => std_logic_vector(to_unsigned(26,8) ,
62961	 => std_logic_vector(to_unsigned(27,8) ,
62962	 => std_logic_vector(to_unsigned(30,8) ,
62963	 => std_logic_vector(to_unsigned(24,8) ,
62964	 => std_logic_vector(to_unsigned(29,8) ,
62965	 => std_logic_vector(to_unsigned(37,8) ,
62966	 => std_logic_vector(to_unsigned(35,8) ,
62967	 => std_logic_vector(to_unsigned(31,8) ,
62968	 => std_logic_vector(to_unsigned(35,8) ,
62969	 => std_logic_vector(to_unsigned(33,8) ,
62970	 => std_logic_vector(to_unsigned(32,8) ,
62971	 => std_logic_vector(to_unsigned(13,8) ,
62972	 => std_logic_vector(to_unsigned(13,8) ,
62973	 => std_logic_vector(to_unsigned(26,8) ,
62974	 => std_logic_vector(to_unsigned(25,8) ,
62975	 => std_logic_vector(to_unsigned(17,8) ,
62976	 => std_logic_vector(to_unsigned(18,8) ,
62977	 => std_logic_vector(to_unsigned(19,8) ,
62978	 => std_logic_vector(to_unsigned(12,8) ,
62979	 => std_logic_vector(to_unsigned(9,8) ,
62980	 => std_logic_vector(to_unsigned(12,8) ,
62981	 => std_logic_vector(to_unsigned(12,8) ,
62982	 => std_logic_vector(to_unsigned(11,8) ,
62983	 => std_logic_vector(to_unsigned(12,8) ,
62984	 => std_logic_vector(to_unsigned(11,8) ,
62985	 => std_logic_vector(to_unsigned(16,8) ,
62986	 => std_logic_vector(to_unsigned(9,8) ,
62987	 => std_logic_vector(to_unsigned(10,8) ,
62988	 => std_logic_vector(to_unsigned(9,8) ,
62989	 => std_logic_vector(to_unsigned(1,8) ,
62990	 => std_logic_vector(to_unsigned(0,8) ,
62991	 => std_logic_vector(to_unsigned(4,8) ,
62992	 => std_logic_vector(to_unsigned(15,8) ,
62993	 => std_logic_vector(to_unsigned(12,8) ,
62994	 => std_logic_vector(to_unsigned(9,8) ,
62995	 => std_logic_vector(to_unsigned(10,8) ,
62996	 => std_logic_vector(to_unsigned(13,8) ,
62997	 => std_logic_vector(to_unsigned(7,8) ,
62998	 => std_logic_vector(to_unsigned(6,8) ,
62999	 => std_logic_vector(to_unsigned(5,8) ,
63000	 => std_logic_vector(to_unsigned(4,8) ,
63001	 => std_logic_vector(to_unsigned(4,8) ,
63002	 => std_logic_vector(to_unsigned(4,8) ,
63003	 => std_logic_vector(to_unsigned(25,8) ,
63004	 => std_logic_vector(to_unsigned(4,8) ,
63005	 => std_logic_vector(to_unsigned(0,8) ,
63006	 => std_logic_vector(to_unsigned(0,8) ,
63007	 => std_logic_vector(to_unsigned(2,8) ,
63008	 => std_logic_vector(to_unsigned(13,8) ,
63009	 => std_logic_vector(to_unsigned(34,8) ,
63010	 => std_logic_vector(to_unsigned(9,8) ,
63011	 => std_logic_vector(to_unsigned(0,8) ,
63012	 => std_logic_vector(to_unsigned(0,8) ,
63013	 => std_logic_vector(to_unsigned(3,8) ,
63014	 => std_logic_vector(to_unsigned(8,8) ,
63015	 => std_logic_vector(to_unsigned(7,8) ,
63016	 => std_logic_vector(to_unsigned(9,8) ,
63017	 => std_logic_vector(to_unsigned(9,8) ,
63018	 => std_logic_vector(to_unsigned(17,8) ,
63019	 => std_logic_vector(to_unsigned(30,8) ,
63020	 => std_logic_vector(to_unsigned(29,8) ,
63021	 => std_logic_vector(to_unsigned(26,8) ,
63022	 => std_logic_vector(to_unsigned(28,8) ,
63023	 => std_logic_vector(to_unsigned(24,8) ,
63024	 => std_logic_vector(to_unsigned(21,8) ,
63025	 => std_logic_vector(to_unsigned(22,8) ,
63026	 => std_logic_vector(to_unsigned(37,8) ,
63027	 => std_logic_vector(to_unsigned(45,8) ,
63028	 => std_logic_vector(to_unsigned(50,8) ,
63029	 => std_logic_vector(to_unsigned(49,8) ,
63030	 => std_logic_vector(to_unsigned(43,8) ,
63031	 => std_logic_vector(to_unsigned(30,8) ,
63032	 => std_logic_vector(to_unsigned(21,8) ,
63033	 => std_logic_vector(to_unsigned(36,8) ,
63034	 => std_logic_vector(to_unsigned(35,8) ,
63035	 => std_logic_vector(to_unsigned(26,8) ,
63036	 => std_logic_vector(to_unsigned(32,8) ,
63037	 => std_logic_vector(to_unsigned(30,8) ,
63038	 => std_logic_vector(to_unsigned(22,8) ,
63039	 => std_logic_vector(to_unsigned(29,8) ,
63040	 => std_logic_vector(to_unsigned(20,8) ,
63041	 => std_logic_vector(to_unsigned(71,8) ,
63042	 => std_logic_vector(to_unsigned(76,8) ,
63043	 => std_logic_vector(to_unsigned(74,8) ,
63044	 => std_logic_vector(to_unsigned(68,8) ,
63045	 => std_logic_vector(to_unsigned(76,8) ,
63046	 => std_logic_vector(to_unsigned(82,8) ,
63047	 => std_logic_vector(to_unsigned(79,8) ,
63048	 => std_logic_vector(to_unsigned(69,8) ,
63049	 => std_logic_vector(to_unsigned(66,8) ,
63050	 => std_logic_vector(to_unsigned(58,8) ,
63051	 => std_logic_vector(to_unsigned(59,8) ,
63052	 => std_logic_vector(to_unsigned(61,8) ,
63053	 => std_logic_vector(to_unsigned(57,8) ,
63054	 => std_logic_vector(to_unsigned(59,8) ,
63055	 => std_logic_vector(to_unsigned(68,8) ,
63056	 => std_logic_vector(to_unsigned(69,8) ,
63057	 => std_logic_vector(to_unsigned(70,8) ,
63058	 => std_logic_vector(to_unsigned(64,8) ,
63059	 => std_logic_vector(to_unsigned(52,8) ,
63060	 => std_logic_vector(to_unsigned(51,8) ,
63061	 => std_logic_vector(to_unsigned(48,8) ,
63062	 => std_logic_vector(to_unsigned(45,8) ,
63063	 => std_logic_vector(to_unsigned(27,8) ,
63064	 => std_logic_vector(to_unsigned(18,8) ,
63065	 => std_logic_vector(to_unsigned(20,8) ,
63066	 => std_logic_vector(to_unsigned(25,8) ,
63067	 => std_logic_vector(to_unsigned(29,8) ,
63068	 => std_logic_vector(to_unsigned(30,8) ,
63069	 => std_logic_vector(to_unsigned(36,8) ,
63070	 => std_logic_vector(to_unsigned(45,8) ,
63071	 => std_logic_vector(to_unsigned(48,8) ,
63072	 => std_logic_vector(to_unsigned(45,8) ,
63073	 => std_logic_vector(to_unsigned(37,8) ,
63074	 => std_logic_vector(to_unsigned(35,8) ,
63075	 => std_logic_vector(to_unsigned(35,8) ,
63076	 => std_logic_vector(to_unsigned(37,8) ,
63077	 => std_logic_vector(to_unsigned(37,8) ,
63078	 => std_logic_vector(to_unsigned(27,8) ,
63079	 => std_logic_vector(to_unsigned(29,8) ,
63080	 => std_logic_vector(to_unsigned(41,8) ,
63081	 => std_logic_vector(to_unsigned(36,8) ,
63082	 => std_logic_vector(to_unsigned(35,8) ,
63083	 => std_logic_vector(to_unsigned(33,8) ,
63084	 => std_logic_vector(to_unsigned(44,8) ,
63085	 => std_logic_vector(to_unsigned(55,8) ,
63086	 => std_logic_vector(to_unsigned(65,8) ,
63087	 => std_logic_vector(to_unsigned(79,8) ,
63088	 => std_logic_vector(to_unsigned(68,8) ,
63089	 => std_logic_vector(to_unsigned(51,8) ,
63090	 => std_logic_vector(to_unsigned(40,8) ,
63091	 => std_logic_vector(to_unsigned(38,8) ,
63092	 => std_logic_vector(to_unsigned(30,8) ,
63093	 => std_logic_vector(to_unsigned(37,8) ,
63094	 => std_logic_vector(to_unsigned(53,8) ,
63095	 => std_logic_vector(to_unsigned(54,8) ,
63096	 => std_logic_vector(to_unsigned(51,8) ,
63097	 => std_logic_vector(to_unsigned(52,8) ,
63098	 => std_logic_vector(to_unsigned(52,8) ,
63099	 => std_logic_vector(to_unsigned(62,8) ,
63100	 => std_logic_vector(to_unsigned(68,8) ,
63101	 => std_logic_vector(to_unsigned(52,8) ,
63102	 => std_logic_vector(to_unsigned(59,8) ,
63103	 => std_logic_vector(to_unsigned(81,8) ,
63104	 => std_logic_vector(to_unsigned(63,8) ,
63105	 => std_logic_vector(to_unsigned(80,8) ,
63106	 => std_logic_vector(to_unsigned(74,8) ,
63107	 => std_logic_vector(to_unsigned(67,8) ,
63108	 => std_logic_vector(to_unsigned(96,8) ,
63109	 => std_logic_vector(to_unsigned(76,8) ,
63110	 => std_logic_vector(to_unsigned(90,8) ,
63111	 => std_logic_vector(to_unsigned(91,8) ,
63112	 => std_logic_vector(to_unsigned(71,8) ,
63113	 => std_logic_vector(to_unsigned(101,8) ,
63114	 => std_logic_vector(to_unsigned(134,8) ,
63115	 => std_logic_vector(to_unsigned(119,8) ,
63116	 => std_logic_vector(to_unsigned(109,8) ,
63117	 => std_logic_vector(to_unsigned(130,8) ,
63118	 => std_logic_vector(to_unsigned(133,8) ,
63119	 => std_logic_vector(to_unsigned(130,8) ,
63120	 => std_logic_vector(to_unsigned(114,8) ,
63121	 => std_logic_vector(to_unsigned(86,8) ,
63122	 => std_logic_vector(to_unsigned(74,8) ,
63123	 => std_logic_vector(to_unsigned(71,8) ,
63124	 => std_logic_vector(to_unsigned(62,8) ,
63125	 => std_logic_vector(to_unsigned(85,8) ,
63126	 => std_logic_vector(to_unsigned(99,8) ,
63127	 => std_logic_vector(to_unsigned(61,8) ,
63128	 => std_logic_vector(to_unsigned(47,8) ,
63129	 => std_logic_vector(to_unsigned(91,8) ,
63130	 => std_logic_vector(to_unsigned(92,8) ,
63131	 => std_logic_vector(to_unsigned(96,8) ,
63132	 => std_logic_vector(to_unsigned(80,8) ,
63133	 => std_logic_vector(to_unsigned(68,8) ,
63134	 => std_logic_vector(to_unsigned(46,8) ,
63135	 => std_logic_vector(to_unsigned(22,8) ,
63136	 => std_logic_vector(to_unsigned(21,8) ,
63137	 => std_logic_vector(to_unsigned(17,8) ,
63138	 => std_logic_vector(to_unsigned(29,8) ,
63139	 => std_logic_vector(to_unsigned(35,8) ,
63140	 => std_logic_vector(to_unsigned(41,8) ,
63141	 => std_logic_vector(to_unsigned(49,8) ,
63142	 => std_logic_vector(to_unsigned(52,8) ,
63143	 => std_logic_vector(to_unsigned(24,8) ,
63144	 => std_logic_vector(to_unsigned(17,8) ,
63145	 => std_logic_vector(to_unsigned(57,8) ,
63146	 => std_logic_vector(to_unsigned(58,8) ,
63147	 => std_logic_vector(to_unsigned(30,8) ,
63148	 => std_logic_vector(to_unsigned(34,8) ,
63149	 => std_logic_vector(to_unsigned(41,8) ,
63150	 => std_logic_vector(to_unsigned(46,8) ,
63151	 => std_logic_vector(to_unsigned(43,8) ,
63152	 => std_logic_vector(to_unsigned(39,8) ,
63153	 => std_logic_vector(to_unsigned(49,8) ,
63154	 => std_logic_vector(to_unsigned(52,8) ,
63155	 => std_logic_vector(to_unsigned(51,8) ,
63156	 => std_logic_vector(to_unsigned(71,8) ,
63157	 => std_logic_vector(to_unsigned(87,8) ,
63158	 => std_logic_vector(to_unsigned(91,8) ,
63159	 => std_logic_vector(to_unsigned(99,8) ,
63160	 => std_logic_vector(to_unsigned(72,8) ,
63161	 => std_logic_vector(to_unsigned(90,8) ,
63162	 => std_logic_vector(to_unsigned(79,8) ,
63163	 => std_logic_vector(to_unsigned(39,8) ,
63164	 => std_logic_vector(to_unsigned(25,8) ,
63165	 => std_logic_vector(to_unsigned(19,8) ,
63166	 => std_logic_vector(to_unsigned(27,8) ,
63167	 => std_logic_vector(to_unsigned(17,8) ,
63168	 => std_logic_vector(to_unsigned(19,8) ,
63169	 => std_logic_vector(to_unsigned(64,8) ,
63170	 => std_logic_vector(to_unsigned(67,8) ,
63171	 => std_logic_vector(to_unsigned(59,8) ,
63172	 => std_logic_vector(to_unsigned(74,8) ,
63173	 => std_logic_vector(to_unsigned(82,8) ,
63174	 => std_logic_vector(to_unsigned(68,8) ,
63175	 => std_logic_vector(to_unsigned(68,8) ,
63176	 => std_logic_vector(to_unsigned(82,8) ,
63177	 => std_logic_vector(to_unsigned(84,8) ,
63178	 => std_logic_vector(to_unsigned(56,8) ,
63179	 => std_logic_vector(to_unsigned(70,8) ,
63180	 => std_logic_vector(to_unsigned(48,8) ,
63181	 => std_logic_vector(to_unsigned(25,8) ,
63182	 => std_logic_vector(to_unsigned(51,8) ,
63183	 => std_logic_vector(to_unsigned(54,8) ,
63184	 => std_logic_vector(to_unsigned(25,8) ,
63185	 => std_logic_vector(to_unsigned(20,8) ,
63186	 => std_logic_vector(to_unsigned(25,8) ,
63187	 => std_logic_vector(to_unsigned(15,8) ,
63188	 => std_logic_vector(to_unsigned(39,8) ,
63189	 => std_logic_vector(to_unsigned(103,8) ,
63190	 => std_logic_vector(to_unsigned(57,8) ,
63191	 => std_logic_vector(to_unsigned(45,8) ,
63192	 => std_logic_vector(to_unsigned(82,8) ,
63193	 => std_logic_vector(to_unsigned(59,8) ,
63194	 => std_logic_vector(to_unsigned(68,8) ,
63195	 => std_logic_vector(to_unsigned(82,8) ,
63196	 => std_logic_vector(to_unsigned(52,8) ,
63197	 => std_logic_vector(to_unsigned(22,8) ,
63198	 => std_logic_vector(to_unsigned(19,8) ,
63199	 => std_logic_vector(to_unsigned(12,8) ,
63200	 => std_logic_vector(to_unsigned(32,8) ,
63201	 => std_logic_vector(to_unsigned(77,8) ,
63202	 => std_logic_vector(to_unsigned(47,8) ,
63203	 => std_logic_vector(to_unsigned(17,8) ,
63204	 => std_logic_vector(to_unsigned(23,8) ,
63205	 => std_logic_vector(to_unsigned(63,8) ,
63206	 => std_logic_vector(to_unsigned(61,8) ,
63207	 => std_logic_vector(to_unsigned(30,8) ,
63208	 => std_logic_vector(to_unsigned(25,8) ,
63209	 => std_logic_vector(to_unsigned(33,8) ,
63210	 => std_logic_vector(to_unsigned(51,8) ,
63211	 => std_logic_vector(to_unsigned(46,8) ,
63212	 => std_logic_vector(to_unsigned(38,8) ,
63213	 => std_logic_vector(to_unsigned(42,8) ,
63214	 => std_logic_vector(to_unsigned(86,8) ,
63215	 => std_logic_vector(to_unsigned(69,8) ,
63216	 => std_logic_vector(to_unsigned(47,8) ,
63217	 => std_logic_vector(to_unsigned(39,8) ,
63218	 => std_logic_vector(to_unsigned(25,8) ,
63219	 => std_logic_vector(to_unsigned(29,8) ,
63220	 => std_logic_vector(to_unsigned(41,8) ,
63221	 => std_logic_vector(to_unsigned(15,8) ,
63222	 => std_logic_vector(to_unsigned(9,8) ,
63223	 => std_logic_vector(to_unsigned(12,8) ,
63224	 => std_logic_vector(to_unsigned(10,8) ,
63225	 => std_logic_vector(to_unsigned(18,8) ,
63226	 => std_logic_vector(to_unsigned(59,8) ,
63227	 => std_logic_vector(to_unsigned(37,8) ,
63228	 => std_logic_vector(to_unsigned(32,8) ,
63229	 => std_logic_vector(to_unsigned(35,8) ,
63230	 => std_logic_vector(to_unsigned(45,8) ,
63231	 => std_logic_vector(to_unsigned(48,8) ,
63232	 => std_logic_vector(to_unsigned(35,8) ,
63233	 => std_logic_vector(to_unsigned(43,8) ,
63234	 => std_logic_vector(to_unsigned(51,8) ,
63235	 => std_logic_vector(to_unsigned(45,8) ,
63236	 => std_logic_vector(to_unsigned(51,8) ,
63237	 => std_logic_vector(to_unsigned(52,8) ,
63238	 => std_logic_vector(to_unsigned(78,8) ,
63239	 => std_logic_vector(to_unsigned(91,8) ,
63240	 => std_logic_vector(to_unsigned(72,8) ,
63241	 => std_logic_vector(to_unsigned(49,8) ,
63242	 => std_logic_vector(to_unsigned(34,8) ,
63243	 => std_logic_vector(to_unsigned(23,8) ,
63244	 => std_logic_vector(to_unsigned(30,8) ,
63245	 => std_logic_vector(to_unsigned(44,8) ,
63246	 => std_logic_vector(to_unsigned(39,8) ,
63247	 => std_logic_vector(to_unsigned(24,8) ,
63248	 => std_logic_vector(to_unsigned(27,8) ,
63249	 => std_logic_vector(to_unsigned(40,8) ,
63250	 => std_logic_vector(to_unsigned(51,8) ,
63251	 => std_logic_vector(to_unsigned(43,8) ,
63252	 => std_logic_vector(to_unsigned(60,8) ,
63253	 => std_logic_vector(to_unsigned(38,8) ,
63254	 => std_logic_vector(to_unsigned(15,8) ,
63255	 => std_logic_vector(to_unsigned(22,8) ,
63256	 => std_logic_vector(to_unsigned(31,8) ,
63257	 => std_logic_vector(to_unsigned(31,8) ,
63258	 => std_logic_vector(to_unsigned(49,8) ,
63259	 => std_logic_vector(to_unsigned(46,8) ,
63260	 => std_logic_vector(to_unsigned(17,8) ,
63261	 => std_logic_vector(to_unsigned(30,8) ,
63262	 => std_logic_vector(to_unsigned(44,8) ,
63263	 => std_logic_vector(to_unsigned(73,8) ,
63264	 => std_logic_vector(to_unsigned(70,8) ,
63265	 => std_logic_vector(to_unsigned(41,8) ,
63266	 => std_logic_vector(to_unsigned(45,8) ,
63267	 => std_logic_vector(to_unsigned(38,8) ,
63268	 => std_logic_vector(to_unsigned(37,8) ,
63269	 => std_logic_vector(to_unsigned(30,8) ,
63270	 => std_logic_vector(to_unsigned(15,8) ,
63271	 => std_logic_vector(to_unsigned(18,8) ,
63272	 => std_logic_vector(to_unsigned(20,8) ,
63273	 => std_logic_vector(to_unsigned(24,8) ,
63274	 => std_logic_vector(to_unsigned(30,8) ,
63275	 => std_logic_vector(to_unsigned(35,8) ,
63276	 => std_logic_vector(to_unsigned(30,8) ,
63277	 => std_logic_vector(to_unsigned(18,8) ,
63278	 => std_logic_vector(to_unsigned(47,8) ,
63279	 => std_logic_vector(to_unsigned(66,8) ,
63280	 => std_logic_vector(to_unsigned(25,8) ,
63281	 => std_logic_vector(to_unsigned(16,8) ,
63282	 => std_logic_vector(to_unsigned(18,8) ,
63283	 => std_logic_vector(to_unsigned(19,8) ,
63284	 => std_logic_vector(to_unsigned(30,8) ,
63285	 => std_logic_vector(to_unsigned(31,8) ,
63286	 => std_logic_vector(to_unsigned(30,8) ,
63287	 => std_logic_vector(to_unsigned(32,8) ,
63288	 => std_logic_vector(to_unsigned(28,8) ,
63289	 => std_logic_vector(to_unsigned(27,8) ,
63290	 => std_logic_vector(to_unsigned(23,8) ,
63291	 => std_logic_vector(to_unsigned(12,8) ,
63292	 => std_logic_vector(to_unsigned(27,8) ,
63293	 => std_logic_vector(to_unsigned(41,8) ,
63294	 => std_logic_vector(to_unsigned(42,8) ,
63295	 => std_logic_vector(to_unsigned(37,8) ,
63296	 => std_logic_vector(to_unsigned(41,8) ,
63297	 => std_logic_vector(to_unsigned(40,8) ,
63298	 => std_logic_vector(to_unsigned(18,8) ,
63299	 => std_logic_vector(to_unsigned(10,8) ,
63300	 => std_logic_vector(to_unsigned(15,8) ,
63301	 => std_logic_vector(to_unsigned(16,8) ,
63302	 => std_logic_vector(to_unsigned(14,8) ,
63303	 => std_logic_vector(to_unsigned(17,8) ,
63304	 => std_logic_vector(to_unsigned(16,8) ,
63305	 => std_logic_vector(to_unsigned(13,8) ,
63306	 => std_logic_vector(to_unsigned(14,8) ,
63307	 => std_logic_vector(to_unsigned(9,8) ,
63308	 => std_logic_vector(to_unsigned(10,8) ,
63309	 => std_logic_vector(to_unsigned(2,8) ,
63310	 => std_logic_vector(to_unsigned(0,8) ,
63311	 => std_logic_vector(to_unsigned(2,8) ,
63312	 => std_logic_vector(to_unsigned(12,8) ,
63313	 => std_logic_vector(to_unsigned(20,8) ,
63314	 => std_logic_vector(to_unsigned(20,8) ,
63315	 => std_logic_vector(to_unsigned(10,8) ,
63316	 => std_logic_vector(to_unsigned(8,8) ,
63317	 => std_logic_vector(to_unsigned(9,8) ,
63318	 => std_logic_vector(to_unsigned(8,8) ,
63319	 => std_logic_vector(to_unsigned(8,8) ,
63320	 => std_logic_vector(to_unsigned(6,8) ,
63321	 => std_logic_vector(to_unsigned(7,8) ,
63322	 => std_logic_vector(to_unsigned(7,8) ,
63323	 => std_logic_vector(to_unsigned(29,8) ,
63324	 => std_logic_vector(to_unsigned(6,8) ,
63325	 => std_logic_vector(to_unsigned(0,8) ,
63326	 => std_logic_vector(to_unsigned(1,8) ,
63327	 => std_logic_vector(to_unsigned(8,8) ,
63328	 => std_logic_vector(to_unsigned(38,8) ,
63329	 => std_logic_vector(to_unsigned(37,8) ,
63330	 => std_logic_vector(to_unsigned(12,8) ,
63331	 => std_logic_vector(to_unsigned(2,8) ,
63332	 => std_logic_vector(to_unsigned(0,8) ,
63333	 => std_logic_vector(to_unsigned(1,8) ,
63334	 => std_logic_vector(to_unsigned(5,8) ,
63335	 => std_logic_vector(to_unsigned(7,8) ,
63336	 => std_logic_vector(to_unsigned(6,8) ,
63337	 => std_logic_vector(to_unsigned(6,8) ,
63338	 => std_logic_vector(to_unsigned(15,8) ,
63339	 => std_logic_vector(to_unsigned(29,8) ,
63340	 => std_logic_vector(to_unsigned(10,8) ,
63341	 => std_logic_vector(to_unsigned(17,8) ,
63342	 => std_logic_vector(to_unsigned(20,8) ,
63343	 => std_logic_vector(to_unsigned(17,8) ,
63344	 => std_logic_vector(to_unsigned(22,8) ,
63345	 => std_logic_vector(to_unsigned(22,8) ,
63346	 => std_logic_vector(to_unsigned(23,8) ,
63347	 => std_logic_vector(to_unsigned(36,8) ,
63348	 => std_logic_vector(to_unsigned(48,8) ,
63349	 => std_logic_vector(to_unsigned(45,8) ,
63350	 => std_logic_vector(to_unsigned(47,8) ,
63351	 => std_logic_vector(to_unsigned(41,8) ,
63352	 => std_logic_vector(to_unsigned(17,8) ,
63353	 => std_logic_vector(to_unsigned(28,8) ,
63354	 => std_logic_vector(to_unsigned(35,8) ,
63355	 => std_logic_vector(to_unsigned(35,8) ,
63356	 => std_logic_vector(to_unsigned(41,8) ,
63357	 => std_logic_vector(to_unsigned(38,8) ,
63358	 => std_logic_vector(to_unsigned(35,8) ,
63359	 => std_logic_vector(to_unsigned(30,8) ,
63360	 => std_logic_vector(to_unsigned(15,8) ,
63361	 => std_logic_vector(to_unsigned(81,8) ,
63362	 => std_logic_vector(to_unsigned(79,8) ,
63363	 => std_logic_vector(to_unsigned(81,8) ,
63364	 => std_logic_vector(to_unsigned(87,8) ,
63365	 => std_logic_vector(to_unsigned(85,8) ,
63366	 => std_logic_vector(to_unsigned(80,8) ,
63367	 => std_logic_vector(to_unsigned(59,8) ,
63368	 => std_logic_vector(to_unsigned(53,8) ,
63369	 => std_logic_vector(to_unsigned(54,8) ,
63370	 => std_logic_vector(to_unsigned(56,8) ,
63371	 => std_logic_vector(to_unsigned(70,8) ,
63372	 => std_logic_vector(to_unsigned(64,8) ,
63373	 => std_logic_vector(to_unsigned(60,8) ,
63374	 => std_logic_vector(to_unsigned(68,8) ,
63375	 => std_logic_vector(to_unsigned(71,8) ,
63376	 => std_logic_vector(to_unsigned(70,8) ,
63377	 => std_logic_vector(to_unsigned(70,8) ,
63378	 => std_logic_vector(to_unsigned(64,8) ,
63379	 => std_logic_vector(to_unsigned(55,8) ,
63380	 => std_logic_vector(to_unsigned(50,8) ,
63381	 => std_logic_vector(to_unsigned(53,8) ,
63382	 => std_logic_vector(to_unsigned(48,8) ,
63383	 => std_logic_vector(to_unsigned(29,8) ,
63384	 => std_logic_vector(to_unsigned(24,8) ,
63385	 => std_logic_vector(to_unsigned(31,8) ,
63386	 => std_logic_vector(to_unsigned(33,8) ,
63387	 => std_logic_vector(to_unsigned(36,8) ,
63388	 => std_logic_vector(to_unsigned(42,8) ,
63389	 => std_logic_vector(to_unsigned(40,8) ,
63390	 => std_logic_vector(to_unsigned(39,8) ,
63391	 => std_logic_vector(to_unsigned(42,8) ,
63392	 => std_logic_vector(to_unsigned(35,8) ,
63393	 => std_logic_vector(to_unsigned(33,8) ,
63394	 => std_logic_vector(to_unsigned(34,8) ,
63395	 => std_logic_vector(to_unsigned(30,8) ,
63396	 => std_logic_vector(to_unsigned(35,8) ,
63397	 => std_logic_vector(to_unsigned(37,8) ,
63398	 => std_logic_vector(to_unsigned(25,8) ,
63399	 => std_logic_vector(to_unsigned(27,8) ,
63400	 => std_logic_vector(to_unsigned(32,8) ,
63401	 => std_logic_vector(to_unsigned(31,8) ,
63402	 => std_logic_vector(to_unsigned(35,8) ,
63403	 => std_logic_vector(to_unsigned(36,8) ,
63404	 => std_logic_vector(to_unsigned(41,8) ,
63405	 => std_logic_vector(to_unsigned(39,8) ,
63406	 => std_logic_vector(to_unsigned(56,8) ,
63407	 => std_logic_vector(to_unsigned(72,8) ,
63408	 => std_logic_vector(to_unsigned(64,8) ,
63409	 => std_logic_vector(to_unsigned(48,8) ,
63410	 => std_logic_vector(to_unsigned(42,8) ,
63411	 => std_logic_vector(to_unsigned(37,8) ,
63412	 => std_logic_vector(to_unsigned(32,8) ,
63413	 => std_logic_vector(to_unsigned(41,8) ,
63414	 => std_logic_vector(to_unsigned(66,8) ,
63415	 => std_logic_vector(to_unsigned(57,8) ,
63416	 => std_logic_vector(to_unsigned(54,8) ,
63417	 => std_logic_vector(to_unsigned(54,8) ,
63418	 => std_logic_vector(to_unsigned(51,8) ,
63419	 => std_logic_vector(to_unsigned(62,8) ,
63420	 => std_logic_vector(to_unsigned(73,8) ,
63421	 => std_logic_vector(to_unsigned(55,8) ,
63422	 => std_logic_vector(to_unsigned(59,8) ,
63423	 => std_logic_vector(to_unsigned(84,8) ,
63424	 => std_logic_vector(to_unsigned(80,8) ,
63425	 => std_logic_vector(to_unsigned(88,8) ,
63426	 => std_logic_vector(to_unsigned(91,8) ,
63427	 => std_logic_vector(to_unsigned(88,8) ,
63428	 => std_logic_vector(to_unsigned(99,8) ,
63429	 => std_logic_vector(to_unsigned(81,8) ,
63430	 => std_logic_vector(to_unsigned(97,8) ,
63431	 => std_logic_vector(to_unsigned(99,8) ,
63432	 => std_logic_vector(to_unsigned(70,8) ,
63433	 => std_logic_vector(to_unsigned(105,8) ,
63434	 => std_logic_vector(to_unsigned(131,8) ,
63435	 => std_logic_vector(to_unsigned(128,8) ,
63436	 => std_logic_vector(to_unsigned(122,8) ,
63437	 => std_logic_vector(to_unsigned(125,8) ,
63438	 => std_logic_vector(to_unsigned(121,8) ,
63439	 => std_logic_vector(to_unsigned(121,8) ,
63440	 => std_logic_vector(to_unsigned(96,8) ,
63441	 => std_logic_vector(to_unsigned(96,8) ,
63442	 => std_logic_vector(to_unsigned(92,8) ,
63443	 => std_logic_vector(to_unsigned(80,8) ,
63444	 => std_logic_vector(to_unsigned(60,8) ,
63445	 => std_logic_vector(to_unsigned(45,8) ,
63446	 => std_logic_vector(to_unsigned(39,8) ,
63447	 => std_logic_vector(to_unsigned(52,8) ,
63448	 => std_logic_vector(to_unsigned(127,8) ,
63449	 => std_logic_vector(to_unsigned(136,8) ,
63450	 => std_logic_vector(to_unsigned(90,8) ,
63451	 => std_logic_vector(to_unsigned(84,8) ,
63452	 => std_logic_vector(to_unsigned(77,8) ,
63453	 => std_logic_vector(to_unsigned(78,8) ,
63454	 => std_logic_vector(to_unsigned(86,8) ,
63455	 => std_logic_vector(to_unsigned(52,8) ,
63456	 => std_logic_vector(to_unsigned(41,8) ,
63457	 => std_logic_vector(to_unsigned(30,8) ,
63458	 => std_logic_vector(to_unsigned(20,8) ,
63459	 => std_logic_vector(to_unsigned(17,8) ,
63460	 => std_logic_vector(to_unsigned(19,8) ,
63461	 => std_logic_vector(to_unsigned(17,8) ,
63462	 => std_logic_vector(to_unsigned(30,8) ,
63463	 => std_logic_vector(to_unsigned(40,8) ,
63464	 => std_logic_vector(to_unsigned(53,8) ,
63465	 => std_logic_vector(to_unsigned(76,8) ,
63466	 => std_logic_vector(to_unsigned(50,8) ,
63467	 => std_logic_vector(to_unsigned(27,8) ,
63468	 => std_logic_vector(to_unsigned(30,8) ,
63469	 => std_logic_vector(to_unsigned(40,8) ,
63470	 => std_logic_vector(to_unsigned(37,8) ,
63471	 => std_logic_vector(to_unsigned(47,8) ,
63472	 => std_logic_vector(to_unsigned(62,8) ,
63473	 => std_logic_vector(to_unsigned(67,8) ,
63474	 => std_logic_vector(to_unsigned(62,8) ,
63475	 => std_logic_vector(to_unsigned(62,8) ,
63476	 => std_logic_vector(to_unsigned(76,8) ,
63477	 => std_logic_vector(to_unsigned(76,8) ,
63478	 => std_logic_vector(to_unsigned(65,8) ,
63479	 => std_logic_vector(to_unsigned(55,8) ,
63480	 => std_logic_vector(to_unsigned(60,8) ,
63481	 => std_logic_vector(to_unsigned(78,8) ,
63482	 => std_logic_vector(to_unsigned(51,8) ,
63483	 => std_logic_vector(to_unsigned(29,8) ,
63484	 => std_logic_vector(to_unsigned(27,8) ,
63485	 => std_logic_vector(to_unsigned(32,8) ,
63486	 => std_logic_vector(to_unsigned(39,8) ,
63487	 => std_logic_vector(to_unsigned(36,8) ,
63488	 => std_logic_vector(to_unsigned(34,8) ,
63489	 => std_logic_vector(to_unsigned(27,8) ,
63490	 => std_logic_vector(to_unsigned(32,8) ,
63491	 => std_logic_vector(to_unsigned(34,8) ,
63492	 => std_logic_vector(to_unsigned(38,8) ,
63493	 => std_logic_vector(to_unsigned(88,8) ,
63494	 => std_logic_vector(to_unsigned(90,8) ,
63495	 => std_logic_vector(to_unsigned(93,8) ,
63496	 => std_logic_vector(to_unsigned(85,8) ,
63497	 => std_logic_vector(to_unsigned(101,8) ,
63498	 => std_logic_vector(to_unsigned(37,8) ,
63499	 => std_logic_vector(to_unsigned(65,8) ,
63500	 => std_logic_vector(to_unsigned(53,8) ,
63501	 => std_logic_vector(to_unsigned(24,8) ,
63502	 => std_logic_vector(to_unsigned(29,8) ,
63503	 => std_logic_vector(to_unsigned(22,8) ,
63504	 => std_logic_vector(to_unsigned(23,8) ,
63505	 => std_logic_vector(to_unsigned(35,8) ,
63506	 => std_logic_vector(to_unsigned(43,8) ,
63507	 => std_logic_vector(to_unsigned(19,8) ,
63508	 => std_logic_vector(to_unsigned(32,8) ,
63509	 => std_logic_vector(to_unsigned(105,8) ,
63510	 => std_logic_vector(to_unsigned(47,8) ,
63511	 => std_logic_vector(to_unsigned(27,8) ,
63512	 => std_logic_vector(to_unsigned(85,8) ,
63513	 => std_logic_vector(to_unsigned(25,8) ,
63514	 => std_logic_vector(to_unsigned(34,8) ,
63515	 => std_logic_vector(to_unsigned(87,8) ,
63516	 => std_logic_vector(to_unsigned(50,8) ,
63517	 => std_logic_vector(to_unsigned(17,8) ,
63518	 => std_logic_vector(to_unsigned(14,8) ,
63519	 => std_logic_vector(to_unsigned(7,8) ,
63520	 => std_logic_vector(to_unsigned(27,8) ,
63521	 => std_logic_vector(to_unsigned(45,8) ,
63522	 => std_logic_vector(to_unsigned(41,8) ,
63523	 => std_logic_vector(to_unsigned(51,8) ,
63524	 => std_logic_vector(to_unsigned(35,8) ,
63525	 => std_logic_vector(to_unsigned(46,8) ,
63526	 => std_logic_vector(to_unsigned(36,8) ,
63527	 => std_logic_vector(to_unsigned(16,8) ,
63528	 => std_logic_vector(to_unsigned(17,8) ,
63529	 => std_logic_vector(to_unsigned(51,8) ,
63530	 => std_logic_vector(to_unsigned(86,8) ,
63531	 => std_logic_vector(to_unsigned(43,8) ,
63532	 => std_logic_vector(to_unsigned(43,8) ,
63533	 => std_logic_vector(to_unsigned(91,8) ,
63534	 => std_logic_vector(to_unsigned(88,8) ,
63535	 => std_logic_vector(to_unsigned(44,8) ,
63536	 => std_logic_vector(to_unsigned(35,8) ,
63537	 => std_logic_vector(to_unsigned(23,8) ,
63538	 => std_logic_vector(to_unsigned(27,8) ,
63539	 => std_logic_vector(to_unsigned(45,8) ,
63540	 => std_logic_vector(to_unsigned(32,8) ,
63541	 => std_logic_vector(to_unsigned(12,8) ,
63542	 => std_logic_vector(to_unsigned(9,8) ,
63543	 => std_logic_vector(to_unsigned(12,8) ,
63544	 => std_logic_vector(to_unsigned(12,8) ,
63545	 => std_logic_vector(to_unsigned(18,8) ,
63546	 => std_logic_vector(to_unsigned(37,8) ,
63547	 => std_logic_vector(to_unsigned(29,8) ,
63548	 => std_logic_vector(to_unsigned(38,8) ,
63549	 => std_logic_vector(to_unsigned(42,8) ,
63550	 => std_logic_vector(to_unsigned(44,8) ,
63551	 => std_logic_vector(to_unsigned(54,8) ,
63552	 => std_logic_vector(to_unsigned(34,8) ,
63553	 => std_logic_vector(to_unsigned(49,8) ,
63554	 => std_logic_vector(to_unsigned(69,8) ,
63555	 => std_logic_vector(to_unsigned(51,8) ,
63556	 => std_logic_vector(to_unsigned(51,8) ,
63557	 => std_logic_vector(to_unsigned(47,8) ,
63558	 => std_logic_vector(to_unsigned(68,8) ,
63559	 => std_logic_vector(to_unsigned(93,8) ,
63560	 => std_logic_vector(to_unsigned(97,8) ,
63561	 => std_logic_vector(to_unsigned(70,8) ,
63562	 => std_logic_vector(to_unsigned(35,8) ,
63563	 => std_logic_vector(to_unsigned(19,8) ,
63564	 => std_logic_vector(to_unsigned(17,8) ,
63565	 => std_logic_vector(to_unsigned(24,8) ,
63566	 => std_logic_vector(to_unsigned(24,8) ,
63567	 => std_logic_vector(to_unsigned(23,8) ,
63568	 => std_logic_vector(to_unsigned(30,8) ,
63569	 => std_logic_vector(to_unsigned(51,8) ,
63570	 => std_logic_vector(to_unsigned(47,8) ,
63571	 => std_logic_vector(to_unsigned(40,8) ,
63572	 => std_logic_vector(to_unsigned(38,8) ,
63573	 => std_logic_vector(to_unsigned(35,8) ,
63574	 => std_logic_vector(to_unsigned(26,8) ,
63575	 => std_logic_vector(to_unsigned(23,8) ,
63576	 => std_logic_vector(to_unsigned(17,8) ,
63577	 => std_logic_vector(to_unsigned(12,8) ,
63578	 => std_logic_vector(to_unsigned(22,8) ,
63579	 => std_logic_vector(to_unsigned(59,8) ,
63580	 => std_logic_vector(to_unsigned(36,8) ,
63581	 => std_logic_vector(to_unsigned(35,8) ,
63582	 => std_logic_vector(to_unsigned(29,8) ,
63583	 => std_logic_vector(to_unsigned(44,8) ,
63584	 => std_logic_vector(to_unsigned(76,8) ,
63585	 => std_logic_vector(to_unsigned(40,8) ,
63586	 => std_logic_vector(to_unsigned(40,8) ,
63587	 => std_logic_vector(to_unsigned(41,8) ,
63588	 => std_logic_vector(to_unsigned(40,8) ,
63589	 => std_logic_vector(to_unsigned(33,8) ,
63590	 => std_logic_vector(to_unsigned(32,8) ,
63591	 => std_logic_vector(to_unsigned(29,8) ,
63592	 => std_logic_vector(to_unsigned(27,8) ,
63593	 => std_logic_vector(to_unsigned(30,8) ,
63594	 => std_logic_vector(to_unsigned(16,8) ,
63595	 => std_logic_vector(to_unsigned(17,8) ,
63596	 => std_logic_vector(to_unsigned(18,8) ,
63597	 => std_logic_vector(to_unsigned(13,8) ,
63598	 => std_logic_vector(to_unsigned(35,8) ,
63599	 => std_logic_vector(to_unsigned(49,8) ,
63600	 => std_logic_vector(to_unsigned(13,8) ,
63601	 => std_logic_vector(to_unsigned(8,8) ,
63602	 => std_logic_vector(to_unsigned(16,8) ,
63603	 => std_logic_vector(to_unsigned(29,8) ,
63604	 => std_logic_vector(to_unsigned(37,8) ,
63605	 => std_logic_vector(to_unsigned(30,8) ,
63606	 => std_logic_vector(to_unsigned(30,8) ,
63607	 => std_logic_vector(to_unsigned(35,8) ,
63608	 => std_logic_vector(to_unsigned(37,8) ,
63609	 => std_logic_vector(to_unsigned(24,8) ,
63610	 => std_logic_vector(to_unsigned(17,8) ,
63611	 => std_logic_vector(to_unsigned(13,8) ,
63612	 => std_logic_vector(to_unsigned(41,8) ,
63613	 => std_logic_vector(to_unsigned(45,8) ,
63614	 => std_logic_vector(to_unsigned(37,8) ,
63615	 => std_logic_vector(to_unsigned(41,8) ,
63616	 => std_logic_vector(to_unsigned(30,8) ,
63617	 => std_logic_vector(to_unsigned(18,8) ,
63618	 => std_logic_vector(to_unsigned(20,8) ,
63619	 => std_logic_vector(to_unsigned(22,8) ,
63620	 => std_logic_vector(to_unsigned(22,8) ,
63621	 => std_logic_vector(to_unsigned(25,8) ,
63622	 => std_logic_vector(to_unsigned(27,8) ,
63623	 => std_logic_vector(to_unsigned(22,8) ,
63624	 => std_logic_vector(to_unsigned(18,8) ,
63625	 => std_logic_vector(to_unsigned(20,8) ,
63626	 => std_logic_vector(to_unsigned(24,8) ,
63627	 => std_logic_vector(to_unsigned(13,8) ,
63628	 => std_logic_vector(to_unsigned(12,8) ,
63629	 => std_logic_vector(to_unsigned(5,8) ,
63630	 => std_logic_vector(to_unsigned(0,8) ,
63631	 => std_logic_vector(to_unsigned(1,8) ,
63632	 => std_logic_vector(to_unsigned(5,8) ,
63633	 => std_logic_vector(to_unsigned(13,8) ,
63634	 => std_logic_vector(to_unsigned(11,8) ,
63635	 => std_logic_vector(to_unsigned(10,8) ,
63636	 => std_logic_vector(to_unsigned(12,8) ,
63637	 => std_logic_vector(to_unsigned(9,8) ,
63638	 => std_logic_vector(to_unsigned(8,8) ,
63639	 => std_logic_vector(to_unsigned(8,8) ,
63640	 => std_logic_vector(to_unsigned(3,8) ,
63641	 => std_logic_vector(to_unsigned(5,8) ,
63642	 => std_logic_vector(to_unsigned(6,8) ,
63643	 => std_logic_vector(to_unsigned(27,8) ,
63644	 => std_logic_vector(to_unsigned(5,8) ,
63645	 => std_logic_vector(to_unsigned(1,8) ,
63646	 => std_logic_vector(to_unsigned(1,8) ,
63647	 => std_logic_vector(to_unsigned(9,8) ,
63648	 => std_logic_vector(to_unsigned(49,8) ,
63649	 => std_logic_vector(to_unsigned(59,8) ,
63650	 => std_logic_vector(to_unsigned(60,8) ,
63651	 => std_logic_vector(to_unsigned(35,8) ,
63652	 => std_logic_vector(to_unsigned(2,8) ,
63653	 => std_logic_vector(to_unsigned(0,8) ,
63654	 => std_logic_vector(to_unsigned(2,8) ,
63655	 => std_logic_vector(to_unsigned(6,8) ,
63656	 => std_logic_vector(to_unsigned(8,8) ,
63657	 => std_logic_vector(to_unsigned(7,8) ,
63658	 => std_logic_vector(to_unsigned(8,8) ,
63659	 => std_logic_vector(to_unsigned(20,8) ,
63660	 => std_logic_vector(to_unsigned(17,8) ,
63661	 => std_logic_vector(to_unsigned(20,8) ,
63662	 => std_logic_vector(to_unsigned(19,8) ,
63663	 => std_logic_vector(to_unsigned(24,8) ,
63664	 => std_logic_vector(to_unsigned(12,8) ,
63665	 => std_logic_vector(to_unsigned(17,8) ,
63666	 => std_logic_vector(to_unsigned(7,8) ,
63667	 => std_logic_vector(to_unsigned(4,8) ,
63668	 => std_logic_vector(to_unsigned(10,8) ,
63669	 => std_logic_vector(to_unsigned(13,8) ,
63670	 => std_logic_vector(to_unsigned(16,8) ,
63671	 => std_logic_vector(to_unsigned(19,8) ,
63672	 => std_logic_vector(to_unsigned(15,8) ,
63673	 => std_logic_vector(to_unsigned(17,8) ,
63674	 => std_logic_vector(to_unsigned(26,8) ,
63675	 => std_logic_vector(to_unsigned(24,8) ,
63676	 => std_logic_vector(to_unsigned(31,8) ,
63677	 => std_logic_vector(to_unsigned(34,8) ,
63678	 => std_logic_vector(to_unsigned(25,8) ,
63679	 => std_logic_vector(to_unsigned(20,8) ,
63680	 => std_logic_vector(to_unsigned(10,8) ,
63681	 => std_logic_vector(to_unsigned(93,8) ,
63682	 => std_logic_vector(to_unsigned(95,8) ,
63683	 => std_logic_vector(to_unsigned(86,8) ,
63684	 => std_logic_vector(to_unsigned(87,8) ,
63685	 => std_logic_vector(to_unsigned(82,8) ,
63686	 => std_logic_vector(to_unsigned(85,8) ,
63687	 => std_logic_vector(to_unsigned(80,8) ,
63688	 => std_logic_vector(to_unsigned(73,8) ,
63689	 => std_logic_vector(to_unsigned(70,8) ,
63690	 => std_logic_vector(to_unsigned(70,8) ,
63691	 => std_logic_vector(to_unsigned(71,8) ,
63692	 => std_logic_vector(to_unsigned(69,8) ,
63693	 => std_logic_vector(to_unsigned(71,8) ,
63694	 => std_logic_vector(to_unsigned(76,8) ,
63695	 => std_logic_vector(to_unsigned(67,8) ,
63696	 => std_logic_vector(to_unsigned(71,8) ,
63697	 => std_logic_vector(to_unsigned(71,8) ,
63698	 => std_logic_vector(to_unsigned(64,8) ,
63699	 => std_logic_vector(to_unsigned(54,8) ,
63700	 => std_logic_vector(to_unsigned(50,8) ,
63701	 => std_logic_vector(to_unsigned(41,8) ,
63702	 => std_logic_vector(to_unsigned(42,8) ,
63703	 => std_logic_vector(to_unsigned(34,8) ,
63704	 => std_logic_vector(to_unsigned(31,8) ,
63705	 => std_logic_vector(to_unsigned(38,8) ,
63706	 => std_logic_vector(to_unsigned(41,8) ,
63707	 => std_logic_vector(to_unsigned(57,8) ,
63708	 => std_logic_vector(to_unsigned(59,8) ,
63709	 => std_logic_vector(to_unsigned(46,8) ,
63710	 => std_logic_vector(to_unsigned(35,8) ,
63711	 => std_logic_vector(to_unsigned(35,8) ,
63712	 => std_logic_vector(to_unsigned(37,8) ,
63713	 => std_logic_vector(to_unsigned(37,8) ,
63714	 => std_logic_vector(to_unsigned(30,8) ,
63715	 => std_logic_vector(to_unsigned(25,8) ,
63716	 => std_logic_vector(to_unsigned(34,8) ,
63717	 => std_logic_vector(to_unsigned(32,8) ,
63718	 => std_logic_vector(to_unsigned(18,8) ,
63719	 => std_logic_vector(to_unsigned(19,8) ,
63720	 => std_logic_vector(to_unsigned(19,8) ,
63721	 => std_logic_vector(to_unsigned(23,8) ,
63722	 => std_logic_vector(to_unsigned(28,8) ,
63723	 => std_logic_vector(to_unsigned(42,8) ,
63724	 => std_logic_vector(to_unsigned(47,8) ,
63725	 => std_logic_vector(to_unsigned(51,8) ,
63726	 => std_logic_vector(to_unsigned(56,8) ,
63727	 => std_logic_vector(to_unsigned(60,8) ,
63728	 => std_logic_vector(to_unsigned(61,8) ,
63729	 => std_logic_vector(to_unsigned(50,8) ,
63730	 => std_logic_vector(to_unsigned(37,8) ,
63731	 => std_logic_vector(to_unsigned(35,8) ,
63732	 => std_logic_vector(to_unsigned(29,8) ,
63733	 => std_logic_vector(to_unsigned(41,8) ,
63734	 => std_logic_vector(to_unsigned(63,8) ,
63735	 => std_logic_vector(to_unsigned(62,8) ,
63736	 => std_logic_vector(to_unsigned(74,8) ,
63737	 => std_logic_vector(to_unsigned(65,8) ,
63738	 => std_logic_vector(to_unsigned(58,8) ,
63739	 => std_logic_vector(to_unsigned(54,8) ,
63740	 => std_logic_vector(to_unsigned(46,8) ,
63741	 => std_logic_vector(to_unsigned(49,8) ,
63742	 => std_logic_vector(to_unsigned(63,8) ,
63743	 => std_logic_vector(to_unsigned(84,8) ,
63744	 => std_logic_vector(to_unsigned(68,8) ,
63745	 => std_logic_vector(to_unsigned(87,8) ,
63746	 => std_logic_vector(to_unsigned(80,8) ,
63747	 => std_logic_vector(to_unsigned(88,8) ,
63748	 => std_logic_vector(to_unsigned(96,8) ,
63749	 => std_logic_vector(to_unsigned(97,8) ,
63750	 => std_logic_vector(to_unsigned(103,8) ,
63751	 => std_logic_vector(to_unsigned(93,8) ,
63752	 => std_logic_vector(to_unsigned(101,8) ,
63753	 => std_logic_vector(to_unsigned(108,8) ,
63754	 => std_logic_vector(to_unsigned(128,8) ,
63755	 => std_logic_vector(to_unsigned(133,8) ,
63756	 => std_logic_vector(to_unsigned(111,8) ,
63757	 => std_logic_vector(to_unsigned(115,8) ,
63758	 => std_logic_vector(to_unsigned(114,8) ,
63759	 => std_logic_vector(to_unsigned(101,8) ,
63760	 => std_logic_vector(to_unsigned(104,8) ,
63761	 => std_logic_vector(to_unsigned(108,8) ,
63762	 => std_logic_vector(to_unsigned(97,8) ,
63763	 => std_logic_vector(to_unsigned(96,8) ,
63764	 => std_logic_vector(to_unsigned(96,8) ,
63765	 => std_logic_vector(to_unsigned(65,8) ,
63766	 => std_logic_vector(to_unsigned(51,8) ,
63767	 => std_logic_vector(to_unsigned(103,8) ,
63768	 => std_logic_vector(to_unsigned(149,8) ,
63769	 => std_logic_vector(to_unsigned(104,8) ,
63770	 => std_logic_vector(to_unsigned(44,8) ,
63771	 => std_logic_vector(to_unsigned(46,8) ,
63772	 => std_logic_vector(to_unsigned(64,8) ,
63773	 => std_logic_vector(to_unsigned(64,8) ,
63774	 => std_logic_vector(to_unsigned(70,8) ,
63775	 => std_logic_vector(to_unsigned(72,8) ,
63776	 => std_logic_vector(to_unsigned(84,8) ,
63777	 => std_logic_vector(to_unsigned(115,8) ,
63778	 => std_logic_vector(to_unsigned(100,8) ,
63779	 => std_logic_vector(to_unsigned(67,8) ,
63780	 => std_logic_vector(to_unsigned(50,8) ,
63781	 => std_logic_vector(to_unsigned(34,8) ,
63782	 => std_logic_vector(to_unsigned(41,8) ,
63783	 => std_logic_vector(to_unsigned(77,8) ,
63784	 => std_logic_vector(to_unsigned(86,8) ,
63785	 => std_logic_vector(to_unsigned(62,8) ,
63786	 => std_logic_vector(to_unsigned(54,8) ,
63787	 => std_logic_vector(to_unsigned(23,8) ,
63788	 => std_logic_vector(to_unsigned(37,8) ,
63789	 => std_logic_vector(to_unsigned(61,8) ,
63790	 => std_logic_vector(to_unsigned(25,8) ,
63791	 => std_logic_vector(to_unsigned(80,8) ,
63792	 => std_logic_vector(to_unsigned(138,8) ,
63793	 => std_logic_vector(to_unsigned(105,8) ,
63794	 => std_logic_vector(to_unsigned(96,8) ,
63795	 => std_logic_vector(to_unsigned(86,8) ,
63796	 => std_logic_vector(to_unsigned(60,8) ,
63797	 => std_logic_vector(to_unsigned(45,8) ,
63798	 => std_logic_vector(to_unsigned(40,8) ,
63799	 => std_logic_vector(to_unsigned(30,8) ,
63800	 => std_logic_vector(to_unsigned(36,8) ,
63801	 => std_logic_vector(to_unsigned(65,8) ,
63802	 => std_logic_vector(to_unsigned(50,8) ,
63803	 => std_logic_vector(to_unsigned(34,8) ,
63804	 => std_logic_vector(to_unsigned(30,8) ,
63805	 => std_logic_vector(to_unsigned(31,8) ,
63806	 => std_logic_vector(to_unsigned(40,8) ,
63807	 => std_logic_vector(to_unsigned(44,8) ,
63808	 => std_logic_vector(to_unsigned(27,8) ,
63809	 => std_logic_vector(to_unsigned(13,8) ,
63810	 => std_logic_vector(to_unsigned(16,8) ,
63811	 => std_logic_vector(to_unsigned(16,8) ,
63812	 => std_logic_vector(to_unsigned(25,8) ,
63813	 => std_logic_vector(to_unsigned(67,8) ,
63814	 => std_logic_vector(to_unsigned(91,8) ,
63815	 => std_logic_vector(to_unsigned(82,8) ,
63816	 => std_logic_vector(to_unsigned(76,8) ,
63817	 => std_logic_vector(to_unsigned(90,8) ,
63818	 => std_logic_vector(to_unsigned(57,8) ,
63819	 => std_logic_vector(to_unsigned(65,8) ,
63820	 => std_logic_vector(to_unsigned(29,8) ,
63821	 => std_logic_vector(to_unsigned(12,8) ,
63822	 => std_logic_vector(to_unsigned(14,8) ,
63823	 => std_logic_vector(to_unsigned(10,8) ,
63824	 => std_logic_vector(to_unsigned(13,8) ,
63825	 => std_logic_vector(to_unsigned(18,8) ,
63826	 => std_logic_vector(to_unsigned(23,8) ,
63827	 => std_logic_vector(to_unsigned(16,8) ,
63828	 => std_logic_vector(to_unsigned(37,8) ,
63829	 => std_logic_vector(to_unsigned(92,8) ,
63830	 => std_logic_vector(to_unsigned(78,8) ,
63831	 => std_logic_vector(to_unsigned(77,8) ,
63832	 => std_logic_vector(to_unsigned(82,8) ,
63833	 => std_logic_vector(to_unsigned(51,8) ,
63834	 => std_logic_vector(to_unsigned(56,8) ,
63835	 => std_logic_vector(to_unsigned(88,8) ,
63836	 => std_logic_vector(to_unsigned(50,8) ,
63837	 => std_logic_vector(to_unsigned(21,8) ,
63838	 => std_logic_vector(to_unsigned(11,8) ,
63839	 => std_logic_vector(to_unsigned(7,8) ,
63840	 => std_logic_vector(to_unsigned(20,8) ,
63841	 => std_logic_vector(to_unsigned(18,8) ,
63842	 => std_logic_vector(to_unsigned(21,8) ,
63843	 => std_logic_vector(to_unsigned(32,8) ,
63844	 => std_logic_vector(to_unsigned(32,8) ,
63845	 => std_logic_vector(to_unsigned(32,8) ,
63846	 => std_logic_vector(to_unsigned(18,8) ,
63847	 => std_logic_vector(to_unsigned(12,8) ,
63848	 => std_logic_vector(to_unsigned(24,8) ,
63849	 => std_logic_vector(to_unsigned(55,8) ,
63850	 => std_logic_vector(to_unsigned(76,8) ,
63851	 => std_logic_vector(to_unsigned(45,8) ,
63852	 => std_logic_vector(to_unsigned(86,8) ,
63853	 => std_logic_vector(to_unsigned(72,8) ,
63854	 => std_logic_vector(to_unsigned(39,8) ,
63855	 => std_logic_vector(to_unsigned(51,8) ,
63856	 => std_logic_vector(to_unsigned(22,8) ,
63857	 => std_logic_vector(to_unsigned(21,8) ,
63858	 => std_logic_vector(to_unsigned(41,8) ,
63859	 => std_logic_vector(to_unsigned(30,8) ,
63860	 => std_logic_vector(to_unsigned(32,8) ,
63861	 => std_logic_vector(to_unsigned(20,8) ,
63862	 => std_logic_vector(to_unsigned(10,8) ,
63863	 => std_logic_vector(to_unsigned(14,8) ,
63864	 => std_logic_vector(to_unsigned(10,8) ,
63865	 => std_logic_vector(to_unsigned(20,8) ,
63866	 => std_logic_vector(to_unsigned(40,8) ,
63867	 => std_logic_vector(to_unsigned(11,8) ,
63868	 => std_logic_vector(to_unsigned(22,8) ,
63869	 => std_logic_vector(to_unsigned(15,8) ,
63870	 => std_logic_vector(to_unsigned(40,8) ,
63871	 => std_logic_vector(to_unsigned(63,8) ,
63872	 => std_logic_vector(to_unsigned(57,8) ,
63873	 => std_logic_vector(to_unsigned(61,8) ,
63874	 => std_logic_vector(to_unsigned(72,8) ,
63875	 => std_logic_vector(to_unsigned(66,8) ,
63876	 => std_logic_vector(to_unsigned(49,8) ,
63877	 => std_logic_vector(to_unsigned(39,8) ,
63878	 => std_logic_vector(to_unsigned(39,8) ,
63879	 => std_logic_vector(to_unsigned(43,8) ,
63880	 => std_logic_vector(to_unsigned(73,8) ,
63881	 => std_logic_vector(to_unsigned(74,8) ,
63882	 => std_logic_vector(to_unsigned(24,8) ,
63883	 => std_logic_vector(to_unsigned(19,8) ,
63884	 => std_logic_vector(to_unsigned(15,8) ,
63885	 => std_logic_vector(to_unsigned(10,8) ,
63886	 => std_logic_vector(to_unsigned(15,8) ,
63887	 => std_logic_vector(to_unsigned(19,8) ,
63888	 => std_logic_vector(to_unsigned(43,8) ,
63889	 => std_logic_vector(to_unsigned(69,8) ,
63890	 => std_logic_vector(to_unsigned(24,8) ,
63891	 => std_logic_vector(to_unsigned(16,8) ,
63892	 => std_logic_vector(to_unsigned(30,8) ,
63893	 => std_logic_vector(to_unsigned(45,8) ,
63894	 => std_logic_vector(to_unsigned(35,8) ,
63895	 => std_logic_vector(to_unsigned(35,8) ,
63896	 => std_logic_vector(to_unsigned(35,8) ,
63897	 => std_logic_vector(to_unsigned(32,8) ,
63898	 => std_logic_vector(to_unsigned(42,8) ,
63899	 => std_logic_vector(to_unsigned(49,8) ,
63900	 => std_logic_vector(to_unsigned(29,8) ,
63901	 => std_logic_vector(to_unsigned(29,8) ,
63902	 => std_logic_vector(to_unsigned(37,8) ,
63903	 => std_logic_vector(to_unsigned(35,8) ,
63904	 => std_logic_vector(to_unsigned(52,8) ,
63905	 => std_logic_vector(to_unsigned(51,8) ,
63906	 => std_logic_vector(to_unsigned(39,8) ,
63907	 => std_logic_vector(to_unsigned(41,8) ,
63908	 => std_logic_vector(to_unsigned(40,8) ,
63909	 => std_logic_vector(to_unsigned(24,8) ,
63910	 => std_logic_vector(to_unsigned(19,8) ,
63911	 => std_logic_vector(to_unsigned(21,8) ,
63912	 => std_logic_vector(to_unsigned(27,8) ,
63913	 => std_logic_vector(to_unsigned(33,8) ,
63914	 => std_logic_vector(to_unsigned(18,8) ,
63915	 => std_logic_vector(to_unsigned(14,8) ,
63916	 => std_logic_vector(to_unsigned(18,8) ,
63917	 => std_logic_vector(to_unsigned(20,8) ,
63918	 => std_logic_vector(to_unsigned(26,8) ,
63919	 => std_logic_vector(to_unsigned(25,8) ,
63920	 => std_logic_vector(to_unsigned(11,8) ,
63921	 => std_logic_vector(to_unsigned(9,8) ,
63922	 => std_logic_vector(to_unsigned(18,8) ,
63923	 => std_logic_vector(to_unsigned(32,8) ,
63924	 => std_logic_vector(to_unsigned(34,8) ,
63925	 => std_logic_vector(to_unsigned(32,8) ,
63926	 => std_logic_vector(to_unsigned(32,8) ,
63927	 => std_logic_vector(to_unsigned(23,8) ,
63928	 => std_logic_vector(to_unsigned(27,8) ,
63929	 => std_logic_vector(to_unsigned(30,8) ,
63930	 => std_logic_vector(to_unsigned(22,8) ,
63931	 => std_logic_vector(to_unsigned(30,8) ,
63932	 => std_logic_vector(to_unsigned(42,8) ,
63933	 => std_logic_vector(to_unsigned(44,8) ,
63934	 => std_logic_vector(to_unsigned(40,8) ,
63935	 => std_logic_vector(to_unsigned(41,8) ,
63936	 => std_logic_vector(to_unsigned(26,8) ,
63937	 => std_logic_vector(to_unsigned(15,8) ,
63938	 => std_logic_vector(to_unsigned(28,8) ,
63939	 => std_logic_vector(to_unsigned(36,8) ,
63940	 => std_logic_vector(to_unsigned(30,8) ,
63941	 => std_logic_vector(to_unsigned(33,8) ,
63942	 => std_logic_vector(to_unsigned(31,8) ,
63943	 => std_logic_vector(to_unsigned(20,8) ,
63944	 => std_logic_vector(to_unsigned(22,8) ,
63945	 => std_logic_vector(to_unsigned(27,8) ,
63946	 => std_logic_vector(to_unsigned(21,8) ,
63947	 => std_logic_vector(to_unsigned(22,8) ,
63948	 => std_logic_vector(to_unsigned(22,8) ,
63949	 => std_logic_vector(to_unsigned(17,8) ,
63950	 => std_logic_vector(to_unsigned(2,8) ,
63951	 => std_logic_vector(to_unsigned(0,8) ,
63952	 => std_logic_vector(to_unsigned(3,8) ,
63953	 => std_logic_vector(to_unsigned(14,8) ,
63954	 => std_logic_vector(to_unsigned(11,8) ,
63955	 => std_logic_vector(to_unsigned(12,8) ,
63956	 => std_logic_vector(to_unsigned(10,8) ,
63957	 => std_logic_vector(to_unsigned(6,8) ,
63958	 => std_logic_vector(to_unsigned(6,8) ,
63959	 => std_logic_vector(to_unsigned(5,8) ,
63960	 => std_logic_vector(to_unsigned(3,8) ,
63961	 => std_logic_vector(to_unsigned(3,8) ,
63962	 => std_logic_vector(to_unsigned(4,8) ,
63963	 => std_logic_vector(to_unsigned(33,8) ,
63964	 => std_logic_vector(to_unsigned(9,8) ,
63965	 => std_logic_vector(to_unsigned(0,8) ,
63966	 => std_logic_vector(to_unsigned(0,8) ,
63967	 => std_logic_vector(to_unsigned(3,8) ,
63968	 => std_logic_vector(to_unsigned(16,8) ,
63969	 => std_logic_vector(to_unsigned(23,8) ,
63970	 => std_logic_vector(to_unsigned(5,8) ,
63971	 => std_logic_vector(to_unsigned(7,8) ,
63972	 => std_logic_vector(to_unsigned(4,8) ,
63973	 => std_logic_vector(to_unsigned(0,8) ,
63974	 => std_logic_vector(to_unsigned(0,8) ,
63975	 => std_logic_vector(to_unsigned(6,8) ,
63976	 => std_logic_vector(to_unsigned(35,8) ,
63977	 => std_logic_vector(to_unsigned(30,8) ,
63978	 => std_logic_vector(to_unsigned(8,8) ,
63979	 => std_logic_vector(to_unsigned(6,8) ,
63980	 => std_logic_vector(to_unsigned(12,8) ,
63981	 => std_logic_vector(to_unsigned(13,8) ,
63982	 => std_logic_vector(to_unsigned(16,8) ,
63983	 => std_logic_vector(to_unsigned(17,8) ,
63984	 => std_logic_vector(to_unsigned(19,8) ,
63985	 => std_logic_vector(to_unsigned(17,8) ,
63986	 => std_logic_vector(to_unsigned(6,8) ,
63987	 => std_logic_vector(to_unsigned(3,8) ,
63988	 => std_logic_vector(to_unsigned(3,8) ,
63989	 => std_logic_vector(to_unsigned(4,8) ,
63990	 => std_logic_vector(to_unsigned(4,8) ,
63991	 => std_logic_vector(to_unsigned(4,8) ,
63992	 => std_logic_vector(to_unsigned(11,8) ,
63993	 => std_logic_vector(to_unsigned(10,8) ,
63994	 => std_logic_vector(to_unsigned(17,8) ,
63995	 => std_logic_vector(to_unsigned(23,8) ,
63996	 => std_logic_vector(to_unsigned(19,8) ,
63997	 => std_logic_vector(to_unsigned(25,8) ,
63998	 => std_logic_vector(to_unsigned(19,8) ,
63999	 => std_logic_vector(to_unsigned(16,8) ,
64000	 => std_logic_vector(to_unsigned(11,8) ,
64001	 => std_logic_vector(to_unsigned(97,8) ,
64002	 => std_logic_vector(to_unsigned(99,8) ,
64003	 => std_logic_vector(to_unsigned(93,8) ,
64004	 => std_logic_vector(to_unsigned(86,8) ,
64005	 => std_logic_vector(to_unsigned(90,8) ,
64006	 => std_logic_vector(to_unsigned(84,8) ,
64007	 => std_logic_vector(to_unsigned(69,8) ,
64008	 => std_logic_vector(to_unsigned(56,8) ,
64009	 => std_logic_vector(to_unsigned(67,8) ,
64010	 => std_logic_vector(to_unsigned(79,8) ,
64011	 => std_logic_vector(to_unsigned(82,8) ,
64012	 => std_logic_vector(to_unsigned(78,8) ,
64013	 => std_logic_vector(to_unsigned(68,8) ,
64014	 => std_logic_vector(to_unsigned(69,8) ,
64015	 => std_logic_vector(to_unsigned(71,8) ,
64016	 => std_logic_vector(to_unsigned(73,8) ,
64017	 => std_logic_vector(to_unsigned(70,8) ,
64018	 => std_logic_vector(to_unsigned(56,8) ,
64019	 => std_logic_vector(to_unsigned(49,8) ,
64020	 => std_logic_vector(to_unsigned(41,8) ,
64021	 => std_logic_vector(to_unsigned(28,8) ,
64022	 => std_logic_vector(to_unsigned(36,8) ,
64023	 => std_logic_vector(to_unsigned(36,8) ,
64024	 => std_logic_vector(to_unsigned(38,8) ,
64025	 => std_logic_vector(to_unsigned(43,8) ,
64026	 => std_logic_vector(to_unsigned(45,8) ,
64027	 => std_logic_vector(to_unsigned(49,8) ,
64028	 => std_logic_vector(to_unsigned(45,8) ,
64029	 => std_logic_vector(to_unsigned(46,8) ,
64030	 => std_logic_vector(to_unsigned(41,8) ,
64031	 => std_logic_vector(to_unsigned(31,8) ,
64032	 => std_logic_vector(to_unsigned(32,8) ,
64033	 => std_logic_vector(to_unsigned(35,8) ,
64034	 => std_logic_vector(to_unsigned(33,8) ,
64035	 => std_logic_vector(to_unsigned(28,8) ,
64036	 => std_logic_vector(to_unsigned(27,8) ,
64037	 => std_logic_vector(to_unsigned(33,8) ,
64038	 => std_logic_vector(to_unsigned(24,8) ,
64039	 => std_logic_vector(to_unsigned(19,8) ,
64040	 => std_logic_vector(to_unsigned(23,8) ,
64041	 => std_logic_vector(to_unsigned(22,8) ,
64042	 => std_logic_vector(to_unsigned(25,8) ,
64043	 => std_logic_vector(to_unsigned(46,8) ,
64044	 => std_logic_vector(to_unsigned(43,8) ,
64045	 => std_logic_vector(to_unsigned(42,8) ,
64046	 => std_logic_vector(to_unsigned(55,8) ,
64047	 => std_logic_vector(to_unsigned(70,8) ,
64048	 => std_logic_vector(to_unsigned(64,8) ,
64049	 => std_logic_vector(to_unsigned(45,8) ,
64050	 => std_logic_vector(to_unsigned(37,8) ,
64051	 => std_logic_vector(to_unsigned(37,8) ,
64052	 => std_logic_vector(to_unsigned(26,8) ,
64053	 => std_logic_vector(to_unsigned(36,8) ,
64054	 => std_logic_vector(to_unsigned(52,8) ,
64055	 => std_logic_vector(to_unsigned(66,8) ,
64056	 => std_logic_vector(to_unsigned(93,8) ,
64057	 => std_logic_vector(to_unsigned(66,8) ,
64058	 => std_logic_vector(to_unsigned(52,8) ,
64059	 => std_logic_vector(to_unsigned(63,8) ,
64060	 => std_logic_vector(to_unsigned(71,8) ,
64061	 => std_logic_vector(to_unsigned(54,8) ,
64062	 => std_logic_vector(to_unsigned(62,8) ,
64063	 => std_logic_vector(to_unsigned(91,8) ,
64064	 => std_logic_vector(to_unsigned(79,8) ,
64065	 => std_logic_vector(to_unsigned(84,8) ,
64066	 => std_logic_vector(to_unsigned(65,8) ,
64067	 => std_logic_vector(to_unsigned(81,8) ,
64068	 => std_logic_vector(to_unsigned(109,8) ,
64069	 => std_logic_vector(to_unsigned(104,8) ,
64070	 => std_logic_vector(to_unsigned(119,8) ,
64071	 => std_logic_vector(to_unsigned(96,8) ,
64072	 => std_logic_vector(to_unsigned(85,8) ,
64073	 => std_logic_vector(to_unsigned(109,8) ,
64074	 => std_logic_vector(to_unsigned(133,8) ,
64075	 => std_logic_vector(to_unsigned(124,8) ,
64076	 => std_logic_vector(to_unsigned(116,8) ,
64077	 => std_logic_vector(to_unsigned(103,8) ,
64078	 => std_logic_vector(to_unsigned(90,8) ,
64079	 => std_logic_vector(to_unsigned(101,8) ,
64080	 => std_logic_vector(to_unsigned(104,8) ,
64081	 => std_logic_vector(to_unsigned(84,8) ,
64082	 => std_logic_vector(to_unsigned(109,8) ,
64083	 => std_logic_vector(to_unsigned(107,8) ,
64084	 => std_logic_vector(to_unsigned(70,8) ,
64085	 => std_logic_vector(to_unsigned(64,8) ,
64086	 => std_logic_vector(to_unsigned(66,8) ,
64087	 => std_logic_vector(to_unsigned(86,8) ,
64088	 => std_logic_vector(to_unsigned(82,8) ,
64089	 => std_logic_vector(to_unsigned(44,8) ,
64090	 => std_logic_vector(to_unsigned(36,8) ,
64091	 => std_logic_vector(to_unsigned(53,8) ,
64092	 => std_logic_vector(to_unsigned(70,8) ,
64093	 => std_logic_vector(to_unsigned(87,8) ,
64094	 => std_logic_vector(to_unsigned(64,8) ,
64095	 => std_logic_vector(to_unsigned(61,8) ,
64096	 => std_logic_vector(to_unsigned(80,8) ,
64097	 => std_logic_vector(to_unsigned(130,8) ,
64098	 => std_logic_vector(to_unsigned(151,8) ,
64099	 => std_logic_vector(to_unsigned(136,8) ,
64100	 => std_logic_vector(to_unsigned(131,8) ,
64101	 => std_logic_vector(to_unsigned(115,8) ,
64102	 => std_logic_vector(to_unsigned(86,8) ,
64103	 => std_logic_vector(to_unsigned(74,8) ,
64104	 => std_logic_vector(to_unsigned(54,8) ,
64105	 => std_logic_vector(to_unsigned(42,8) ,
64106	 => std_logic_vector(to_unsigned(45,8) ,
64107	 => std_logic_vector(to_unsigned(27,8) ,
64108	 => std_logic_vector(to_unsigned(23,8) ,
64109	 => std_logic_vector(to_unsigned(31,8) ,
64110	 => std_logic_vector(to_unsigned(17,8) ,
64111	 => std_logic_vector(to_unsigned(72,8) ,
64112	 => std_logic_vector(to_unsigned(177,8) ,
64113	 => std_logic_vector(to_unsigned(154,8) ,
64114	 => std_logic_vector(to_unsigned(149,8) ,
64115	 => std_logic_vector(to_unsigned(138,8) ,
64116	 => std_logic_vector(to_unsigned(68,8) ,
64117	 => std_logic_vector(to_unsigned(68,8) ,
64118	 => std_logic_vector(to_unsigned(71,8) ,
64119	 => std_logic_vector(to_unsigned(59,8) ,
64120	 => std_logic_vector(to_unsigned(81,8) ,
64121	 => std_logic_vector(to_unsigned(82,8) ,
64122	 => std_logic_vector(to_unsigned(87,8) ,
64123	 => std_logic_vector(to_unsigned(76,8) ,
64124	 => std_logic_vector(to_unsigned(50,8) ,
64125	 => std_logic_vector(to_unsigned(49,8) ,
64126	 => std_logic_vector(to_unsigned(29,8) ,
64127	 => std_logic_vector(to_unsigned(18,8) ,
64128	 => std_logic_vector(to_unsigned(18,8) ,
64129	 => std_logic_vector(to_unsigned(17,8) ,
64130	 => std_logic_vector(to_unsigned(23,8) ,
64131	 => std_logic_vector(to_unsigned(23,8) ,
64132	 => std_logic_vector(to_unsigned(31,8) ,
64133	 => std_logic_vector(to_unsigned(82,8) ,
64134	 => std_logic_vector(to_unsigned(100,8) ,
64135	 => std_logic_vector(to_unsigned(87,8) ,
64136	 => std_logic_vector(to_unsigned(79,8) ,
64137	 => std_logic_vector(to_unsigned(67,8) ,
64138	 => std_logic_vector(to_unsigned(85,8) ,
64139	 => std_logic_vector(to_unsigned(97,8) ,
64140	 => std_logic_vector(to_unsigned(41,8) ,
64141	 => std_logic_vector(to_unsigned(9,8) ,
64142	 => std_logic_vector(to_unsigned(9,8) ,
64143	 => std_logic_vector(to_unsigned(6,8) ,
64144	 => std_logic_vector(to_unsigned(10,8) ,
64145	 => std_logic_vector(to_unsigned(11,8) ,
64146	 => std_logic_vector(to_unsigned(20,8) ,
64147	 => std_logic_vector(to_unsigned(6,8) ,
64148	 => std_logic_vector(to_unsigned(25,8) ,
64149	 => std_logic_vector(to_unsigned(100,8) ,
64150	 => std_logic_vector(to_unsigned(86,8) ,
64151	 => std_logic_vector(to_unsigned(84,8) ,
64152	 => std_logic_vector(to_unsigned(86,8) ,
64153	 => std_logic_vector(to_unsigned(99,8) ,
64154	 => std_logic_vector(to_unsigned(90,8) ,
64155	 => std_logic_vector(to_unsigned(87,8) ,
64156	 => std_logic_vector(to_unsigned(54,8) ,
64157	 => std_logic_vector(to_unsigned(16,8) ,
64158	 => std_logic_vector(to_unsigned(11,8) ,
64159	 => std_logic_vector(to_unsigned(10,8) ,
64160	 => std_logic_vector(to_unsigned(23,8) ,
64161	 => std_logic_vector(to_unsigned(26,8) ,
64162	 => std_logic_vector(to_unsigned(9,8) ,
64163	 => std_logic_vector(to_unsigned(8,8) ,
64164	 => std_logic_vector(to_unsigned(32,8) ,
64165	 => std_logic_vector(to_unsigned(24,8) ,
64166	 => std_logic_vector(to_unsigned(15,8) ,
64167	 => std_logic_vector(to_unsigned(12,8) ,
64168	 => std_logic_vector(to_unsigned(22,8) ,
64169	 => std_logic_vector(to_unsigned(60,8) ,
64170	 => std_logic_vector(to_unsigned(92,8) ,
64171	 => std_logic_vector(to_unsigned(92,8) ,
64172	 => std_logic_vector(to_unsigned(74,8) ,
64173	 => std_logic_vector(to_unsigned(53,8) ,
64174	 => std_logic_vector(to_unsigned(35,8) ,
64175	 => std_logic_vector(to_unsigned(34,8) ,
64176	 => std_logic_vector(to_unsigned(54,8) ,
64177	 => std_logic_vector(to_unsigned(48,8) ,
64178	 => std_logic_vector(to_unsigned(29,8) ,
64179	 => std_logic_vector(to_unsigned(30,8) ,
64180	 => std_logic_vector(to_unsigned(63,8) ,
64181	 => std_logic_vector(to_unsigned(24,8) ,
64182	 => std_logic_vector(to_unsigned(11,8) ,
64183	 => std_logic_vector(to_unsigned(13,8) ,
64184	 => std_logic_vector(to_unsigned(10,8) ,
64185	 => std_logic_vector(to_unsigned(28,8) ,
64186	 => std_logic_vector(to_unsigned(49,8) ,
64187	 => std_logic_vector(to_unsigned(16,8) ,
64188	 => std_logic_vector(to_unsigned(18,8) ,
64189	 => std_logic_vector(to_unsigned(7,8) ,
64190	 => std_logic_vector(to_unsigned(32,8) ,
64191	 => std_logic_vector(to_unsigned(62,8) ,
64192	 => std_logic_vector(to_unsigned(26,8) ,
64193	 => std_logic_vector(to_unsigned(31,8) ,
64194	 => std_logic_vector(to_unsigned(32,8) ,
64195	 => std_logic_vector(to_unsigned(55,8) ,
64196	 => std_logic_vector(to_unsigned(63,8) ,
64197	 => std_logic_vector(to_unsigned(30,8) ,
64198	 => std_logic_vector(to_unsigned(36,8) ,
64199	 => std_logic_vector(to_unsigned(32,8) ,
64200	 => std_logic_vector(to_unsigned(47,8) ,
64201	 => std_logic_vector(to_unsigned(59,8) ,
64202	 => std_logic_vector(to_unsigned(23,8) ,
64203	 => std_logic_vector(to_unsigned(25,8) ,
64204	 => std_logic_vector(to_unsigned(28,8) ,
64205	 => std_logic_vector(to_unsigned(18,8) ,
64206	 => std_logic_vector(to_unsigned(16,8) ,
64207	 => std_logic_vector(to_unsigned(22,8) ,
64208	 => std_logic_vector(to_unsigned(80,8) ,
64209	 => std_logic_vector(to_unsigned(68,8) ,
64210	 => std_logic_vector(to_unsigned(22,8) ,
64211	 => std_logic_vector(to_unsigned(15,8) ,
64212	 => std_logic_vector(to_unsigned(30,8) ,
64213	 => std_logic_vector(to_unsigned(41,8) ,
64214	 => std_logic_vector(to_unsigned(37,8) ,
64215	 => std_logic_vector(to_unsigned(45,8) ,
64216	 => std_logic_vector(to_unsigned(43,8) ,
64217	 => std_logic_vector(to_unsigned(38,8) ,
64218	 => std_logic_vector(to_unsigned(45,8) ,
64219	 => std_logic_vector(to_unsigned(44,8) ,
64220	 => std_logic_vector(to_unsigned(30,8) ,
64221	 => std_logic_vector(to_unsigned(30,8) ,
64222	 => std_logic_vector(to_unsigned(30,8) ,
64223	 => std_logic_vector(to_unsigned(30,8) ,
64224	 => std_logic_vector(to_unsigned(42,8) ,
64225	 => std_logic_vector(to_unsigned(51,8) ,
64226	 => std_logic_vector(to_unsigned(45,8) ,
64227	 => std_logic_vector(to_unsigned(32,8) ,
64228	 => std_logic_vector(to_unsigned(31,8) ,
64229	 => std_logic_vector(to_unsigned(41,8) ,
64230	 => std_logic_vector(to_unsigned(30,8) ,
64231	 => std_logic_vector(to_unsigned(22,8) ,
64232	 => std_logic_vector(to_unsigned(25,8) ,
64233	 => std_logic_vector(to_unsigned(38,8) ,
64234	 => std_logic_vector(to_unsigned(12,8) ,
64235	 => std_logic_vector(to_unsigned(8,8) ,
64236	 => std_logic_vector(to_unsigned(12,8) ,
64237	 => std_logic_vector(to_unsigned(14,8) ,
64238	 => std_logic_vector(to_unsigned(16,8) ,
64239	 => std_logic_vector(to_unsigned(15,8) ,
64240	 => std_logic_vector(to_unsigned(15,8) ,
64241	 => std_logic_vector(to_unsigned(22,8) ,
64242	 => std_logic_vector(to_unsigned(19,8) ,
64243	 => std_logic_vector(to_unsigned(22,8) ,
64244	 => std_logic_vector(to_unsigned(21,8) ,
64245	 => std_logic_vector(to_unsigned(25,8) ,
64246	 => std_logic_vector(to_unsigned(27,8) ,
64247	 => std_logic_vector(to_unsigned(14,8) ,
64248	 => std_logic_vector(to_unsigned(15,8) ,
64249	 => std_logic_vector(to_unsigned(31,8) ,
64250	 => std_logic_vector(to_unsigned(30,8) ,
64251	 => std_logic_vector(to_unsigned(40,8) ,
64252	 => std_logic_vector(to_unsigned(39,8) ,
64253	 => std_logic_vector(to_unsigned(37,8) ,
64254	 => std_logic_vector(to_unsigned(35,8) ,
64255	 => std_logic_vector(to_unsigned(41,8) ,
64256	 => std_logic_vector(to_unsigned(29,8) ,
64257	 => std_logic_vector(to_unsigned(20,8) ,
64258	 => std_logic_vector(to_unsigned(27,8) ,
64259	 => std_logic_vector(to_unsigned(34,8) ,
64260	 => std_logic_vector(to_unsigned(30,8) ,
64261	 => std_logic_vector(to_unsigned(28,8) ,
64262	 => std_logic_vector(to_unsigned(25,8) ,
64263	 => std_logic_vector(to_unsigned(26,8) ,
64264	 => std_logic_vector(to_unsigned(32,8) ,
64265	 => std_logic_vector(to_unsigned(31,8) ,
64266	 => std_logic_vector(to_unsigned(19,8) ,
64267	 => std_logic_vector(to_unsigned(19,8) ,
64268	 => std_logic_vector(to_unsigned(29,8) ,
64269	 => std_logic_vector(to_unsigned(35,8) ,
64270	 => std_logic_vector(to_unsigned(8,8) ,
64271	 => std_logic_vector(to_unsigned(0,8) ,
64272	 => std_logic_vector(to_unsigned(2,8) ,
64273	 => std_logic_vector(to_unsigned(32,8) ,
64274	 => std_logic_vector(to_unsigned(37,8) ,
64275	 => std_logic_vector(to_unsigned(22,8) ,
64276	 => std_logic_vector(to_unsigned(21,8) ,
64277	 => std_logic_vector(to_unsigned(16,8) ,
64278	 => std_logic_vector(to_unsigned(12,8) ,
64279	 => std_logic_vector(to_unsigned(15,8) ,
64280	 => std_logic_vector(to_unsigned(11,8) ,
64281	 => std_logic_vector(to_unsigned(11,8) ,
64282	 => std_logic_vector(to_unsigned(16,8) ,
64283	 => std_logic_vector(to_unsigned(24,8) ,
64284	 => std_logic_vector(to_unsigned(6,8) ,
64285	 => std_logic_vector(to_unsigned(0,8) ,
64286	 => std_logic_vector(to_unsigned(0,8) ,
64287	 => std_logic_vector(to_unsigned(13,8) ,
64288	 => std_logic_vector(to_unsigned(42,8) ,
64289	 => std_logic_vector(to_unsigned(37,8) ,
64290	 => std_logic_vector(to_unsigned(20,8) ,
64291	 => std_logic_vector(to_unsigned(18,8) ,
64292	 => std_logic_vector(to_unsigned(30,8) ,
64293	 => std_logic_vector(to_unsigned(3,8) ,
64294	 => std_logic_vector(to_unsigned(0,8) ,
64295	 => std_logic_vector(to_unsigned(4,8) ,
64296	 => std_logic_vector(to_unsigned(29,8) ,
64297	 => std_logic_vector(to_unsigned(57,8) ,
64298	 => std_logic_vector(to_unsigned(49,8) ,
64299	 => std_logic_vector(to_unsigned(16,8) ,
64300	 => std_logic_vector(to_unsigned(5,8) ,
64301	 => std_logic_vector(to_unsigned(9,8) ,
64302	 => std_logic_vector(to_unsigned(8,8) ,
64303	 => std_logic_vector(to_unsigned(7,8) ,
64304	 => std_logic_vector(to_unsigned(9,8) ,
64305	 => std_logic_vector(to_unsigned(11,8) ,
64306	 => std_logic_vector(to_unsigned(9,8) ,
64307	 => std_logic_vector(to_unsigned(9,8) ,
64308	 => std_logic_vector(to_unsigned(9,8) ,
64309	 => std_logic_vector(to_unsigned(8,8) ,
64310	 => std_logic_vector(to_unsigned(8,8) ,
64311	 => std_logic_vector(to_unsigned(8,8) ,
64312	 => std_logic_vector(to_unsigned(20,8) ,
64313	 => std_logic_vector(to_unsigned(25,8) ,
64314	 => std_logic_vector(to_unsigned(29,8) ,
64315	 => std_logic_vector(to_unsigned(36,8) ,
64316	 => std_logic_vector(to_unsigned(27,8) ,
64317	 => std_logic_vector(to_unsigned(26,8) ,
64318	 => std_logic_vector(to_unsigned(21,8) ,
64319	 => std_logic_vector(to_unsigned(16,8) ,
64320	 => std_logic_vector(to_unsigned(8,8) ,
64321	 => std_logic_vector(to_unsigned(101,8) ,
64322	 => std_logic_vector(to_unsigned(95,8) ,
64323	 => std_logic_vector(to_unsigned(101,8) ,
64324	 => std_logic_vector(to_unsigned(95,8) ,
64325	 => std_logic_vector(to_unsigned(85,8) ,
64326	 => std_logic_vector(to_unsigned(67,8) ,
64327	 => std_logic_vector(to_unsigned(43,8) ,
64328	 => std_logic_vector(to_unsigned(53,8) ,
64329	 => std_logic_vector(to_unsigned(79,8) ,
64330	 => std_logic_vector(to_unsigned(87,8) ,
64331	 => std_logic_vector(to_unsigned(85,8) ,
64332	 => std_logic_vector(to_unsigned(79,8) ,
64333	 => std_logic_vector(to_unsigned(73,8) ,
64334	 => std_logic_vector(to_unsigned(69,8) ,
64335	 => std_logic_vector(to_unsigned(64,8) ,
64336	 => std_logic_vector(to_unsigned(61,8) ,
64337	 => std_logic_vector(to_unsigned(54,8) ,
64338	 => std_logic_vector(to_unsigned(53,8) ,
64339	 => std_logic_vector(to_unsigned(42,8) ,
64340	 => std_logic_vector(to_unsigned(29,8) ,
64341	 => std_logic_vector(to_unsigned(21,8) ,
64342	 => std_logic_vector(to_unsigned(29,8) ,
64343	 => std_logic_vector(to_unsigned(45,8) ,
64344	 => std_logic_vector(to_unsigned(50,8) ,
64345	 => std_logic_vector(to_unsigned(41,8) ,
64346	 => std_logic_vector(to_unsigned(37,8) ,
64347	 => std_logic_vector(to_unsigned(33,8) ,
64348	 => std_logic_vector(to_unsigned(30,8) ,
64349	 => std_logic_vector(to_unsigned(35,8) ,
64350	 => std_logic_vector(to_unsigned(35,8) ,
64351	 => std_logic_vector(to_unsigned(32,8) ,
64352	 => std_logic_vector(to_unsigned(32,8) ,
64353	 => std_logic_vector(to_unsigned(35,8) ,
64354	 => std_logic_vector(to_unsigned(32,8) ,
64355	 => std_logic_vector(to_unsigned(26,8) ,
64356	 => std_logic_vector(to_unsigned(29,8) ,
64357	 => std_logic_vector(to_unsigned(29,8) ,
64358	 => std_logic_vector(to_unsigned(20,8) ,
64359	 => std_logic_vector(to_unsigned(23,8) ,
64360	 => std_logic_vector(to_unsigned(23,8) ,
64361	 => std_logic_vector(to_unsigned(24,8) ,
64362	 => std_logic_vector(to_unsigned(25,8) ,
64363	 => std_logic_vector(to_unsigned(34,8) ,
64364	 => std_logic_vector(to_unsigned(45,8) ,
64365	 => std_logic_vector(to_unsigned(40,8) ,
64366	 => std_logic_vector(to_unsigned(45,8) ,
64367	 => std_logic_vector(to_unsigned(63,8) ,
64368	 => std_logic_vector(to_unsigned(66,8) ,
64369	 => std_logic_vector(to_unsigned(44,8) ,
64370	 => std_logic_vector(to_unsigned(35,8) ,
64371	 => std_logic_vector(to_unsigned(29,8) ,
64372	 => std_logic_vector(to_unsigned(24,8) ,
64373	 => std_logic_vector(to_unsigned(40,8) ,
64374	 => std_logic_vector(to_unsigned(51,8) ,
64375	 => std_logic_vector(to_unsigned(78,8) ,
64376	 => std_logic_vector(to_unsigned(125,8) ,
64377	 => std_logic_vector(to_unsigned(77,8) ,
64378	 => std_logic_vector(to_unsigned(47,8) ,
64379	 => std_logic_vector(to_unsigned(52,8) ,
64380	 => std_logic_vector(to_unsigned(51,8) ,
64381	 => std_logic_vector(to_unsigned(41,8) ,
64382	 => std_logic_vector(to_unsigned(56,8) ,
64383	 => std_logic_vector(to_unsigned(69,8) ,
64384	 => std_logic_vector(to_unsigned(69,8) ,
64385	 => std_logic_vector(to_unsigned(88,8) ,
64386	 => std_logic_vector(to_unsigned(73,8) ,
64387	 => std_logic_vector(to_unsigned(68,8) ,
64388	 => std_logic_vector(to_unsigned(91,8) ,
64389	 => std_logic_vector(to_unsigned(104,8) ,
64390	 => std_logic_vector(to_unsigned(115,8) ,
64391	 => std_logic_vector(to_unsigned(105,8) ,
64392	 => std_logic_vector(to_unsigned(100,8) ,
64393	 => std_logic_vector(to_unsigned(122,8) ,
64394	 => std_logic_vector(to_unsigned(127,8) ,
64395	 => std_logic_vector(to_unsigned(122,8) ,
64396	 => std_logic_vector(to_unsigned(111,8) ,
64397	 => std_logic_vector(to_unsigned(100,8) ,
64398	 => std_logic_vector(to_unsigned(95,8) ,
64399	 => std_logic_vector(to_unsigned(82,8) ,
64400	 => std_logic_vector(to_unsigned(80,8) ,
64401	 => std_logic_vector(to_unsigned(77,8) ,
64402	 => std_logic_vector(to_unsigned(105,8) ,
64403	 => std_logic_vector(to_unsigned(81,8) ,
64404	 => std_logic_vector(to_unsigned(45,8) ,
64405	 => std_logic_vector(to_unsigned(66,8) ,
64406	 => std_logic_vector(to_unsigned(65,8) ,
64407	 => std_logic_vector(to_unsigned(69,8) ,
64408	 => std_logic_vector(to_unsigned(82,8) ,
64409	 => std_logic_vector(to_unsigned(40,8) ,
64410	 => std_logic_vector(to_unsigned(34,8) ,
64411	 => std_logic_vector(to_unsigned(59,8) ,
64412	 => std_logic_vector(to_unsigned(79,8) ,
64413	 => std_logic_vector(to_unsigned(90,8) ,
64414	 => std_logic_vector(to_unsigned(69,8) ,
64415	 => std_logic_vector(to_unsigned(108,8) ,
64416	 => std_logic_vector(to_unsigned(92,8) ,
64417	 => std_logic_vector(to_unsigned(51,8) ,
64418	 => std_logic_vector(to_unsigned(53,8) ,
64419	 => std_logic_vector(to_unsigned(77,8) ,
64420	 => std_logic_vector(to_unsigned(81,8) ,
64421	 => std_logic_vector(to_unsigned(82,8) ,
64422	 => std_logic_vector(to_unsigned(54,8) ,
64423	 => std_logic_vector(to_unsigned(54,8) ,
64424	 => std_logic_vector(to_unsigned(47,8) ,
64425	 => std_logic_vector(to_unsigned(41,8) ,
64426	 => std_logic_vector(to_unsigned(30,8) ,
64427	 => std_logic_vector(to_unsigned(17,8) ,
64428	 => std_logic_vector(to_unsigned(17,8) ,
64429	 => std_logic_vector(to_unsigned(29,8) ,
64430	 => std_logic_vector(to_unsigned(28,8) ,
64431	 => std_logic_vector(to_unsigned(62,8) ,
64432	 => std_logic_vector(to_unsigned(109,8) ,
64433	 => std_logic_vector(to_unsigned(91,8) ,
64434	 => std_logic_vector(to_unsigned(121,8) ,
64435	 => std_logic_vector(to_unsigned(128,8) ,
64436	 => std_logic_vector(to_unsigned(69,8) ,
64437	 => std_logic_vector(to_unsigned(84,8) ,
64438	 => std_logic_vector(to_unsigned(95,8) ,
64439	 => std_logic_vector(to_unsigned(95,8) ,
64440	 => std_logic_vector(to_unsigned(93,8) ,
64441	 => std_logic_vector(to_unsigned(86,8) ,
64442	 => std_logic_vector(to_unsigned(78,8) ,
64443	 => std_logic_vector(to_unsigned(93,8) ,
64444	 => std_logic_vector(to_unsigned(90,8) ,
64445	 => std_logic_vector(to_unsigned(92,8) ,
64446	 => std_logic_vector(to_unsigned(38,8) ,
64447	 => std_logic_vector(to_unsigned(17,8) ,
64448	 => std_logic_vector(to_unsigned(24,8) ,
64449	 => std_logic_vector(to_unsigned(18,8) ,
64450	 => std_logic_vector(to_unsigned(22,8) ,
64451	 => std_logic_vector(to_unsigned(23,8) ,
64452	 => std_logic_vector(to_unsigned(26,8) ,
64453	 => std_logic_vector(to_unsigned(58,8) ,
64454	 => std_logic_vector(to_unsigned(76,8) ,
64455	 => std_logic_vector(to_unsigned(82,8) ,
64456	 => std_logic_vector(to_unsigned(32,8) ,
64457	 => std_logic_vector(to_unsigned(29,8) ,
64458	 => std_logic_vector(to_unsigned(80,8) ,
64459	 => std_logic_vector(to_unsigned(78,8) ,
64460	 => std_logic_vector(to_unsigned(37,8) ,
64461	 => std_logic_vector(to_unsigned(10,8) ,
64462	 => std_logic_vector(to_unsigned(13,8) ,
64463	 => std_logic_vector(to_unsigned(14,8) ,
64464	 => std_logic_vector(to_unsigned(13,8) ,
64465	 => std_logic_vector(to_unsigned(16,8) ,
64466	 => std_logic_vector(to_unsigned(34,8) ,
64467	 => std_logic_vector(to_unsigned(13,8) ,
64468	 => std_logic_vector(to_unsigned(24,8) ,
64469	 => std_logic_vector(to_unsigned(107,8) ,
64470	 => std_logic_vector(to_unsigned(79,8) ,
64471	 => std_logic_vector(to_unsigned(65,8) ,
64472	 => std_logic_vector(to_unsigned(92,8) ,
64473	 => std_logic_vector(to_unsigned(69,8) ,
64474	 => std_logic_vector(to_unsigned(70,8) ,
64475	 => std_logic_vector(to_unsigned(95,8) ,
64476	 => std_logic_vector(to_unsigned(52,8) ,
64477	 => std_logic_vector(to_unsigned(16,8) ,
64478	 => std_logic_vector(to_unsigned(12,8) ,
64479	 => std_logic_vector(to_unsigned(7,8) ,
64480	 => std_logic_vector(to_unsigned(24,8) ,
64481	 => std_logic_vector(to_unsigned(42,8) ,
64482	 => std_logic_vector(to_unsigned(11,8) ,
64483	 => std_logic_vector(to_unsigned(16,8) ,
64484	 => std_logic_vector(to_unsigned(40,8) ,
64485	 => std_logic_vector(to_unsigned(32,8) ,
64486	 => std_logic_vector(to_unsigned(20,8) ,
64487	 => std_logic_vector(to_unsigned(17,8) ,
64488	 => std_logic_vector(to_unsigned(31,8) ,
64489	 => std_logic_vector(to_unsigned(57,8) ,
64490	 => std_logic_vector(to_unsigned(77,8) ,
64491	 => std_logic_vector(to_unsigned(76,8) ,
64492	 => std_logic_vector(to_unsigned(47,8) ,
64493	 => std_logic_vector(to_unsigned(48,8) ,
64494	 => std_logic_vector(to_unsigned(24,8) ,
64495	 => std_logic_vector(to_unsigned(25,8) ,
64496	 => std_logic_vector(to_unsigned(45,8) ,
64497	 => std_logic_vector(to_unsigned(27,8) ,
64498	 => std_logic_vector(to_unsigned(35,8) ,
64499	 => std_logic_vector(to_unsigned(69,8) ,
64500	 => std_logic_vector(to_unsigned(35,8) ,
64501	 => std_logic_vector(to_unsigned(10,8) ,
64502	 => std_logic_vector(to_unsigned(10,8) ,
64503	 => std_logic_vector(to_unsigned(13,8) ,
64504	 => std_logic_vector(to_unsigned(13,8) ,
64505	 => std_logic_vector(to_unsigned(24,8) ,
64506	 => std_logic_vector(to_unsigned(47,8) ,
64507	 => std_logic_vector(to_unsigned(37,8) ,
64508	 => std_logic_vector(to_unsigned(41,8) ,
64509	 => std_logic_vector(to_unsigned(32,8) ,
64510	 => std_logic_vector(to_unsigned(45,8) ,
64511	 => std_logic_vector(to_unsigned(57,8) ,
64512	 => std_logic_vector(to_unsigned(30,8) ,
64513	 => std_logic_vector(to_unsigned(28,8) ,
64514	 => std_logic_vector(to_unsigned(24,8) ,
64515	 => std_logic_vector(to_unsigned(42,8) ,
64516	 => std_logic_vector(to_unsigned(60,8) ,
64517	 => std_logic_vector(to_unsigned(16,8) ,
64518	 => std_logic_vector(to_unsigned(16,8) ,
64519	 => std_logic_vector(to_unsigned(13,8) ,
64520	 => std_logic_vector(to_unsigned(31,8) ,
64521	 => std_logic_vector(to_unsigned(58,8) ,
64522	 => std_logic_vector(to_unsigned(36,8) ,
64523	 => std_logic_vector(to_unsigned(24,8) ,
64524	 => std_logic_vector(to_unsigned(20,8) ,
64525	 => std_logic_vector(to_unsigned(28,8) ,
64526	 => std_logic_vector(to_unsigned(23,8) ,
64527	 => std_logic_vector(to_unsigned(24,8) ,
64528	 => std_logic_vector(to_unsigned(59,8) ,
64529	 => std_logic_vector(to_unsigned(35,8) ,
64530	 => std_logic_vector(to_unsigned(36,8) ,
64531	 => std_logic_vector(to_unsigned(32,8) ,
64532	 => std_logic_vector(to_unsigned(35,8) ,
64533	 => std_logic_vector(to_unsigned(35,8) ,
64534	 => std_logic_vector(to_unsigned(50,8) ,
64535	 => std_logic_vector(to_unsigned(63,8) ,
64536	 => std_logic_vector(to_unsigned(62,8) ,
64537	 => std_logic_vector(to_unsigned(66,8) ,
64538	 => std_logic_vector(to_unsigned(50,8) ,
64539	 => std_logic_vector(to_unsigned(44,8) ,
64540	 => std_logic_vector(to_unsigned(47,8) ,
64541	 => std_logic_vector(to_unsigned(84,8) ,
64542	 => std_logic_vector(to_unsigned(69,8) ,
64543	 => std_logic_vector(to_unsigned(48,8) ,
64544	 => std_logic_vector(to_unsigned(51,8) ,
64545	 => std_logic_vector(to_unsigned(41,8) ,
64546	 => std_logic_vector(to_unsigned(46,8) ,
64547	 => std_logic_vector(to_unsigned(37,8) ,
64548	 => std_logic_vector(to_unsigned(33,8) ,
64549	 => std_logic_vector(to_unsigned(28,8) ,
64550	 => std_logic_vector(to_unsigned(21,8) ,
64551	 => std_logic_vector(to_unsigned(22,8) ,
64552	 => std_logic_vector(to_unsigned(35,8) ,
64553	 => std_logic_vector(to_unsigned(37,8) ,
64554	 => std_logic_vector(to_unsigned(30,8) ,
64555	 => std_logic_vector(to_unsigned(36,8) ,
64556	 => std_logic_vector(to_unsigned(60,8) ,
64557	 => std_logic_vector(to_unsigned(76,8) ,
64558	 => std_logic_vector(to_unsigned(30,8) ,
64559	 => std_logic_vector(to_unsigned(13,8) ,
64560	 => std_logic_vector(to_unsigned(13,8) ,
64561	 => std_logic_vector(to_unsigned(29,8) ,
64562	 => std_logic_vector(to_unsigned(15,8) ,
64563	 => std_logic_vector(to_unsigned(12,8) ,
64564	 => std_logic_vector(to_unsigned(15,8) ,
64565	 => std_logic_vector(to_unsigned(16,8) ,
64566	 => std_logic_vector(to_unsigned(20,8) ,
64567	 => std_logic_vector(to_unsigned(31,8) ,
64568	 => std_logic_vector(to_unsigned(25,8) ,
64569	 => std_logic_vector(to_unsigned(19,8) ,
64570	 => std_logic_vector(to_unsigned(29,8) ,
64571	 => std_logic_vector(to_unsigned(40,8) ,
64572	 => std_logic_vector(to_unsigned(39,8) ,
64573	 => std_logic_vector(to_unsigned(37,8) ,
64574	 => std_logic_vector(to_unsigned(20,8) ,
64575	 => std_logic_vector(to_unsigned(29,8) ,
64576	 => std_logic_vector(to_unsigned(22,8) ,
64577	 => std_logic_vector(to_unsigned(14,8) ,
64578	 => std_logic_vector(to_unsigned(18,8) ,
64579	 => std_logic_vector(to_unsigned(28,8) ,
64580	 => std_logic_vector(to_unsigned(23,8) ,
64581	 => std_logic_vector(to_unsigned(16,8) ,
64582	 => std_logic_vector(to_unsigned(15,8) ,
64583	 => std_logic_vector(to_unsigned(19,8) ,
64584	 => std_logic_vector(to_unsigned(18,8) ,
64585	 => std_logic_vector(to_unsigned(16,8) ,
64586	 => std_logic_vector(to_unsigned(27,8) ,
64587	 => std_logic_vector(to_unsigned(33,8) ,
64588	 => std_logic_vector(to_unsigned(32,8) ,
64589	 => std_logic_vector(to_unsigned(36,8) ,
64590	 => std_logic_vector(to_unsigned(13,8) ,
64591	 => std_logic_vector(to_unsigned(0,8) ,
64592	 => std_logic_vector(to_unsigned(0,8) ,
64593	 => std_logic_vector(to_unsigned(29,8) ,
64594	 => std_logic_vector(to_unsigned(44,8) ,
64595	 => std_logic_vector(to_unsigned(17,8) ,
64596	 => std_logic_vector(to_unsigned(28,8) ,
64597	 => std_logic_vector(to_unsigned(34,8) ,
64598	 => std_logic_vector(to_unsigned(29,8) ,
64599	 => std_logic_vector(to_unsigned(32,8) ,
64600	 => std_logic_vector(to_unsigned(16,8) ,
64601	 => std_logic_vector(to_unsigned(16,8) ,
64602	 => std_logic_vector(to_unsigned(17,8) ,
64603	 => std_logic_vector(to_unsigned(8,8) ,
64604	 => std_logic_vector(to_unsigned(5,8) ,
64605	 => std_logic_vector(to_unsigned(1,8) ,
64606	 => std_logic_vector(to_unsigned(1,8) ,
64607	 => std_logic_vector(to_unsigned(9,8) ,
64608	 => std_logic_vector(to_unsigned(18,8) ,
64609	 => std_logic_vector(to_unsigned(13,8) ,
64610	 => std_logic_vector(to_unsigned(17,8) ,
64611	 => std_logic_vector(to_unsigned(52,8) ,
64612	 => std_logic_vector(to_unsigned(77,8) ,
64613	 => std_logic_vector(to_unsigned(11,8) ,
64614	 => std_logic_vector(to_unsigned(0,8) ,
64615	 => std_logic_vector(to_unsigned(0,8) ,
64616	 => std_logic_vector(to_unsigned(8,8) ,
64617	 => std_logic_vector(to_unsigned(47,8) ,
64618	 => std_logic_vector(to_unsigned(47,8) ,
64619	 => std_logic_vector(to_unsigned(20,8) ,
64620	 => std_logic_vector(to_unsigned(8,8) ,
64621	 => std_logic_vector(to_unsigned(14,8) ,
64622	 => std_logic_vector(to_unsigned(13,8) ,
64623	 => std_logic_vector(to_unsigned(12,8) ,
64624	 => std_logic_vector(to_unsigned(11,8) ,
64625	 => std_logic_vector(to_unsigned(20,8) ,
64626	 => std_logic_vector(to_unsigned(7,8) ,
64627	 => std_logic_vector(to_unsigned(10,8) ,
64628	 => std_logic_vector(to_unsigned(8,8) ,
64629	 => std_logic_vector(to_unsigned(8,8) ,
64630	 => std_logic_vector(to_unsigned(8,8) ,
64631	 => std_logic_vector(to_unsigned(7,8) ,
64632	 => std_logic_vector(to_unsigned(12,8) ,
64633	 => std_logic_vector(to_unsigned(18,8) ,
64634	 => std_logic_vector(to_unsigned(24,8) ,
64635	 => std_logic_vector(to_unsigned(25,8) ,
64636	 => std_logic_vector(to_unsigned(32,8) ,
64637	 => std_logic_vector(to_unsigned(32,8) ,
64638	 => std_logic_vector(to_unsigned(26,8) ,
64639	 => std_logic_vector(to_unsigned(13,8) ,
64640	 => std_logic_vector(to_unsigned(6,8) ,
64641	 => std_logic_vector(to_unsigned(111,8) ,
64642	 => std_logic_vector(to_unsigned(101,8) ,
64643	 => std_logic_vector(to_unsigned(97,8) ,
64644	 => std_logic_vector(to_unsigned(103,8) ,
64645	 => std_logic_vector(to_unsigned(77,8) ,
64646	 => std_logic_vector(to_unsigned(63,8) ,
64647	 => std_logic_vector(to_unsigned(73,8) ,
64648	 => std_logic_vector(to_unsigned(96,8) ,
64649	 => std_logic_vector(to_unsigned(91,8) ,
64650	 => std_logic_vector(to_unsigned(86,8) ,
64651	 => std_logic_vector(to_unsigned(80,8) ,
64652	 => std_logic_vector(to_unsigned(81,8) ,
64653	 => std_logic_vector(to_unsigned(81,8) ,
64654	 => std_logic_vector(to_unsigned(71,8) ,
64655	 => std_logic_vector(to_unsigned(61,8) ,
64656	 => std_logic_vector(to_unsigned(42,8) ,
64657	 => std_logic_vector(to_unsigned(40,8) ,
64658	 => std_logic_vector(to_unsigned(30,8) ,
64659	 => std_logic_vector(to_unsigned(35,8) ,
64660	 => std_logic_vector(to_unsigned(30,8) ,
64661	 => std_logic_vector(to_unsigned(15,8) ,
64662	 => std_logic_vector(to_unsigned(36,8) ,
64663	 => std_logic_vector(to_unsigned(51,8) ,
64664	 => std_logic_vector(to_unsigned(37,8) ,
64665	 => std_logic_vector(to_unsigned(39,8) ,
64666	 => std_logic_vector(to_unsigned(41,8) ,
64667	 => std_logic_vector(to_unsigned(39,8) ,
64668	 => std_logic_vector(to_unsigned(37,8) ,
64669	 => std_logic_vector(to_unsigned(29,8) ,
64670	 => std_logic_vector(to_unsigned(33,8) ,
64671	 => std_logic_vector(to_unsigned(40,8) ,
64672	 => std_logic_vector(to_unsigned(33,8) ,
64673	 => std_logic_vector(to_unsigned(25,8) ,
64674	 => std_logic_vector(to_unsigned(30,8) ,
64675	 => std_logic_vector(to_unsigned(36,8) ,
64676	 => std_logic_vector(to_unsigned(35,8) ,
64677	 => std_logic_vector(to_unsigned(29,8) ,
64678	 => std_logic_vector(to_unsigned(19,8) ,
64679	 => std_logic_vector(to_unsigned(21,8) ,
64680	 => std_logic_vector(to_unsigned(17,8) ,
64681	 => std_logic_vector(to_unsigned(19,8) ,
64682	 => std_logic_vector(to_unsigned(25,8) ,
64683	 => std_logic_vector(to_unsigned(37,8) ,
64684	 => std_logic_vector(to_unsigned(52,8) ,
64685	 => std_logic_vector(to_unsigned(51,8) ,
64686	 => std_logic_vector(to_unsigned(51,8) ,
64687	 => std_logic_vector(to_unsigned(56,8) ,
64688	 => std_logic_vector(to_unsigned(55,8) ,
64689	 => std_logic_vector(to_unsigned(42,8) ,
64690	 => std_logic_vector(to_unsigned(37,8) ,
64691	 => std_logic_vector(to_unsigned(29,8) ,
64692	 => std_logic_vector(to_unsigned(25,8) ,
64693	 => std_logic_vector(to_unsigned(39,8) ,
64694	 => std_logic_vector(to_unsigned(51,8) ,
64695	 => std_logic_vector(to_unsigned(51,8) ,
64696	 => std_logic_vector(to_unsigned(62,8) ,
64697	 => std_logic_vector(to_unsigned(58,8) ,
64698	 => std_logic_vector(to_unsigned(45,8) ,
64699	 => std_logic_vector(to_unsigned(50,8) ,
64700	 => std_logic_vector(to_unsigned(50,8) ,
64701	 => std_logic_vector(to_unsigned(40,8) ,
64702	 => std_logic_vector(to_unsigned(58,8) ,
64703	 => std_logic_vector(to_unsigned(66,8) ,
64704	 => std_logic_vector(to_unsigned(48,8) ,
64705	 => std_logic_vector(to_unsigned(58,8) ,
64706	 => std_logic_vector(to_unsigned(51,8) ,
64707	 => std_logic_vector(to_unsigned(61,8) ,
64708	 => std_logic_vector(to_unsigned(65,8) ,
64709	 => std_logic_vector(to_unsigned(62,8) ,
64710	 => std_logic_vector(to_unsigned(95,8) ,
64711	 => std_logic_vector(to_unsigned(97,8) ,
64712	 => std_logic_vector(to_unsigned(82,8) ,
64713	 => std_logic_vector(to_unsigned(105,8) ,
64714	 => std_logic_vector(to_unsigned(127,8) ,
64715	 => std_logic_vector(to_unsigned(121,8) ,
64716	 => std_logic_vector(to_unsigned(109,8) ,
64717	 => std_logic_vector(to_unsigned(105,8) ,
64718	 => std_logic_vector(to_unsigned(111,8) ,
64719	 => std_logic_vector(to_unsigned(67,8) ,
64720	 => std_logic_vector(to_unsigned(39,8) ,
64721	 => std_logic_vector(to_unsigned(41,8) ,
64722	 => std_logic_vector(to_unsigned(80,8) ,
64723	 => std_logic_vector(to_unsigned(112,8) ,
64724	 => std_logic_vector(to_unsigned(91,8) ,
64725	 => std_logic_vector(to_unsigned(74,8) ,
64726	 => std_logic_vector(to_unsigned(72,8) ,
64727	 => std_logic_vector(to_unsigned(72,8) ,
64728	 => std_logic_vector(to_unsigned(63,8) ,
64729	 => std_logic_vector(to_unsigned(44,8) ,
64730	 => std_logic_vector(to_unsigned(49,8) ,
64731	 => std_logic_vector(to_unsigned(53,8) ,
64732	 => std_logic_vector(to_unsigned(53,8) ,
64733	 => std_logic_vector(to_unsigned(58,8) ,
64734	 => std_logic_vector(to_unsigned(65,8) ,
64735	 => std_logic_vector(to_unsigned(74,8) ,
64736	 => std_logic_vector(to_unsigned(72,8) ,
64737	 => std_logic_vector(to_unsigned(51,8) ,
64738	 => std_logic_vector(to_unsigned(47,8) ,
64739	 => std_logic_vector(to_unsigned(52,8) ,
64740	 => std_logic_vector(to_unsigned(33,8) ,
64741	 => std_logic_vector(to_unsigned(41,8) ,
64742	 => std_logic_vector(to_unsigned(40,8) ,
64743	 => std_logic_vector(to_unsigned(54,8) ,
64744	 => std_logic_vector(to_unsigned(45,8) ,
64745	 => std_logic_vector(to_unsigned(39,8) ,
64746	 => std_logic_vector(to_unsigned(29,8) ,
64747	 => std_logic_vector(to_unsigned(18,8) ,
64748	 => std_logic_vector(to_unsigned(22,8) ,
64749	 => std_logic_vector(to_unsigned(45,8) ,
64750	 => std_logic_vector(to_unsigned(52,8) ,
64751	 => std_logic_vector(to_unsigned(58,8) ,
64752	 => std_logic_vector(to_unsigned(52,8) ,
64753	 => std_logic_vector(to_unsigned(37,8) ,
64754	 => std_logic_vector(to_unsigned(59,8) ,
64755	 => std_logic_vector(to_unsigned(68,8) ,
64756	 => std_logic_vector(to_unsigned(32,8) ,
64757	 => std_logic_vector(to_unsigned(41,8) ,
64758	 => std_logic_vector(to_unsigned(54,8) ,
64759	 => std_logic_vector(to_unsigned(67,8) ,
64760	 => std_logic_vector(to_unsigned(80,8) ,
64761	 => std_logic_vector(to_unsigned(45,8) ,
64762	 => std_logic_vector(to_unsigned(52,8) ,
64763	 => std_logic_vector(to_unsigned(103,8) ,
64764	 => std_logic_vector(to_unsigned(115,8) ,
64765	 => std_logic_vector(to_unsigned(96,8) ,
64766	 => std_logic_vector(to_unsigned(30,8) ,
64767	 => std_logic_vector(to_unsigned(20,8) ,
64768	 => std_logic_vector(to_unsigned(23,8) ,
64769	 => std_logic_vector(to_unsigned(15,8) ,
64770	 => std_logic_vector(to_unsigned(11,8) ,
64771	 => std_logic_vector(to_unsigned(17,8) ,
64772	 => std_logic_vector(to_unsigned(22,8) ,
64773	 => std_logic_vector(to_unsigned(34,8) ,
64774	 => std_logic_vector(to_unsigned(73,8) ,
64775	 => std_logic_vector(to_unsigned(85,8) ,
64776	 => std_logic_vector(to_unsigned(30,8) ,
64777	 => std_logic_vector(to_unsigned(51,8) ,
64778	 => std_logic_vector(to_unsigned(87,8) ,
64779	 => std_logic_vector(to_unsigned(79,8) ,
64780	 => std_logic_vector(to_unsigned(41,8) ,
64781	 => std_logic_vector(to_unsigned(8,8) ,
64782	 => std_logic_vector(to_unsigned(17,8) ,
64783	 => std_logic_vector(to_unsigned(24,8) ,
64784	 => std_logic_vector(to_unsigned(15,8) ,
64785	 => std_logic_vector(to_unsigned(22,8) ,
64786	 => std_logic_vector(to_unsigned(29,8) ,
64787	 => std_logic_vector(to_unsigned(15,8) ,
64788	 => std_logic_vector(to_unsigned(32,8) ,
64789	 => std_logic_vector(to_unsigned(93,8) ,
64790	 => std_logic_vector(to_unsigned(85,8) ,
64791	 => std_logic_vector(to_unsigned(79,8) ,
64792	 => std_logic_vector(to_unsigned(90,8) ,
64793	 => std_logic_vector(to_unsigned(55,8) ,
64794	 => std_logic_vector(to_unsigned(61,8) ,
64795	 => std_logic_vector(to_unsigned(95,8) ,
64796	 => std_logic_vector(to_unsigned(50,8) ,
64797	 => std_logic_vector(to_unsigned(19,8) ,
64798	 => std_logic_vector(to_unsigned(10,8) ,
64799	 => std_logic_vector(to_unsigned(4,8) ,
64800	 => std_logic_vector(to_unsigned(15,8) ,
64801	 => std_logic_vector(to_unsigned(22,8) ,
64802	 => std_logic_vector(to_unsigned(9,8) ,
64803	 => std_logic_vector(to_unsigned(18,8) ,
64804	 => std_logic_vector(to_unsigned(40,8) ,
64805	 => std_logic_vector(to_unsigned(35,8) ,
64806	 => std_logic_vector(to_unsigned(19,8) ,
64807	 => std_logic_vector(to_unsigned(19,8) ,
64808	 => std_logic_vector(to_unsigned(39,8) ,
64809	 => std_logic_vector(to_unsigned(63,8) ,
64810	 => std_logic_vector(to_unsigned(39,8) ,
64811	 => std_logic_vector(to_unsigned(33,8) ,
64812	 => std_logic_vector(to_unsigned(45,8) ,
64813	 => std_logic_vector(to_unsigned(23,8) ,
64814	 => std_logic_vector(to_unsigned(22,8) ,
64815	 => std_logic_vector(to_unsigned(31,8) ,
64816	 => std_logic_vector(to_unsigned(22,8) ,
64817	 => std_logic_vector(to_unsigned(34,8) ,
64818	 => std_logic_vector(to_unsigned(64,8) ,
64819	 => std_logic_vector(to_unsigned(43,8) ,
64820	 => std_logic_vector(to_unsigned(29,8) ,
64821	 => std_logic_vector(to_unsigned(13,8) ,
64822	 => std_logic_vector(to_unsigned(10,8) ,
64823	 => std_logic_vector(to_unsigned(16,8) ,
64824	 => std_logic_vector(to_unsigned(12,8) ,
64825	 => std_logic_vector(to_unsigned(16,8) ,
64826	 => std_logic_vector(to_unsigned(42,8) ,
64827	 => std_logic_vector(to_unsigned(53,8) ,
64828	 => std_logic_vector(to_unsigned(54,8) ,
64829	 => std_logic_vector(to_unsigned(59,8) ,
64830	 => std_logic_vector(to_unsigned(59,8) ,
64831	 => std_logic_vector(to_unsigned(57,8) ,
64832	 => std_logic_vector(to_unsigned(60,8) ,
64833	 => std_logic_vector(to_unsigned(50,8) ,
64834	 => std_logic_vector(to_unsigned(43,8) ,
64835	 => std_logic_vector(to_unsigned(47,8) ,
64836	 => std_logic_vector(to_unsigned(53,8) ,
64837	 => std_logic_vector(to_unsigned(28,8) ,
64838	 => std_logic_vector(to_unsigned(20,8) ,
64839	 => std_logic_vector(to_unsigned(8,8) ,
64840	 => std_logic_vector(to_unsigned(27,8) ,
64841	 => std_logic_vector(to_unsigned(52,8) ,
64842	 => std_logic_vector(to_unsigned(27,8) ,
64843	 => std_logic_vector(to_unsigned(12,8) ,
64844	 => std_logic_vector(to_unsigned(25,8) ,
64845	 => std_logic_vector(to_unsigned(46,8) ,
64846	 => std_logic_vector(to_unsigned(29,8) ,
64847	 => std_logic_vector(to_unsigned(18,8) ,
64848	 => std_logic_vector(to_unsigned(39,8) ,
64849	 => std_logic_vector(to_unsigned(25,8) ,
64850	 => std_logic_vector(to_unsigned(31,8) ,
64851	 => std_logic_vector(to_unsigned(29,8) ,
64852	 => std_logic_vector(to_unsigned(32,8) ,
64853	 => std_logic_vector(to_unsigned(37,8) ,
64854	 => std_logic_vector(to_unsigned(44,8) ,
64855	 => std_logic_vector(to_unsigned(46,8) ,
64856	 => std_logic_vector(to_unsigned(45,8) ,
64857	 => std_logic_vector(to_unsigned(52,8) ,
64858	 => std_logic_vector(to_unsigned(43,8) ,
64859	 => std_logic_vector(to_unsigned(26,8) ,
64860	 => std_logic_vector(to_unsigned(26,8) ,
64861	 => std_logic_vector(to_unsigned(57,8) ,
64862	 => std_logic_vector(to_unsigned(54,8) ,
64863	 => std_logic_vector(to_unsigned(65,8) ,
64864	 => std_logic_vector(to_unsigned(69,8) ,
64865	 => std_logic_vector(to_unsigned(49,8) ,
64866	 => std_logic_vector(to_unsigned(37,8) ,
64867	 => std_logic_vector(to_unsigned(37,8) ,
64868	 => std_logic_vector(to_unsigned(27,8) ,
64869	 => std_logic_vector(to_unsigned(22,8) ,
64870	 => std_logic_vector(to_unsigned(26,8) ,
64871	 => std_logic_vector(to_unsigned(30,8) ,
64872	 => std_logic_vector(to_unsigned(33,8) ,
64873	 => std_logic_vector(to_unsigned(41,8) ,
64874	 => std_logic_vector(to_unsigned(52,8) ,
64875	 => std_logic_vector(to_unsigned(73,8) ,
64876	 => std_logic_vector(to_unsigned(82,8) ,
64877	 => std_logic_vector(to_unsigned(122,8) ,
64878	 => std_logic_vector(to_unsigned(67,8) ,
64879	 => std_logic_vector(to_unsigned(23,8) ,
64880	 => std_logic_vector(to_unsigned(28,8) ,
64881	 => std_logic_vector(to_unsigned(39,8) ,
64882	 => std_logic_vector(to_unsigned(29,8) ,
64883	 => std_logic_vector(to_unsigned(23,8) ,
64884	 => std_logic_vector(to_unsigned(18,8) ,
64885	 => std_logic_vector(to_unsigned(14,8) ,
64886	 => std_logic_vector(to_unsigned(12,8) ,
64887	 => std_logic_vector(to_unsigned(16,8) ,
64888	 => std_logic_vector(to_unsigned(10,8) ,
64889	 => std_logic_vector(to_unsigned(10,8) ,
64890	 => std_logic_vector(to_unsigned(33,8) ,
64891	 => std_logic_vector(to_unsigned(43,8) ,
64892	 => std_logic_vector(to_unsigned(46,8) ,
64893	 => std_logic_vector(to_unsigned(46,8) ,
64894	 => std_logic_vector(to_unsigned(18,8) ,
64895	 => std_logic_vector(to_unsigned(12,8) ,
64896	 => std_logic_vector(to_unsigned(24,8) ,
64897	 => std_logic_vector(to_unsigned(23,8) ,
64898	 => std_logic_vector(to_unsigned(26,8) ,
64899	 => std_logic_vector(to_unsigned(23,8) ,
64900	 => std_logic_vector(to_unsigned(10,8) ,
64901	 => std_logic_vector(to_unsigned(14,8) ,
64902	 => std_logic_vector(to_unsigned(13,8) ,
64903	 => std_logic_vector(to_unsigned(13,8) ,
64904	 => std_logic_vector(to_unsigned(16,8) ,
64905	 => std_logic_vector(to_unsigned(17,8) ,
64906	 => std_logic_vector(to_unsigned(23,8) ,
64907	 => std_logic_vector(to_unsigned(22,8) ,
64908	 => std_logic_vector(to_unsigned(25,8) ,
64909	 => std_logic_vector(to_unsigned(24,8) ,
64910	 => std_logic_vector(to_unsigned(13,8) ,
64911	 => std_logic_vector(to_unsigned(1,8) ,
64912	 => std_logic_vector(to_unsigned(0,8) ,
64913	 => std_logic_vector(to_unsigned(12,8) ,
64914	 => std_logic_vector(to_unsigned(42,8) ,
64915	 => std_logic_vector(to_unsigned(24,8) ,
64916	 => std_logic_vector(to_unsigned(29,8) ,
64917	 => std_logic_vector(to_unsigned(33,8) ,
64918	 => std_logic_vector(to_unsigned(29,8) ,
64919	 => std_logic_vector(to_unsigned(20,8) ,
64920	 => std_logic_vector(to_unsigned(8,8) ,
64921	 => std_logic_vector(to_unsigned(13,8) ,
64922	 => std_logic_vector(to_unsigned(18,8) ,
64923	 => std_logic_vector(to_unsigned(12,8) ,
64924	 => std_logic_vector(to_unsigned(8,8) ,
64925	 => std_logic_vector(to_unsigned(1,8) ,
64926	 => std_logic_vector(to_unsigned(1,8) ,
64927	 => std_logic_vector(to_unsigned(7,8) ,
64928	 => std_logic_vector(to_unsigned(19,8) ,
64929	 => std_logic_vector(to_unsigned(11,8) ,
64930	 => std_logic_vector(to_unsigned(5,8) ,
64931	 => std_logic_vector(to_unsigned(12,8) ,
64932	 => std_logic_vector(to_unsigned(23,8) ,
64933	 => std_logic_vector(to_unsigned(12,8) ,
64934	 => std_logic_vector(to_unsigned(1,8) ,
64935	 => std_logic_vector(to_unsigned(0,8) ,
64936	 => std_logic_vector(to_unsigned(2,8) ,
64937	 => std_logic_vector(to_unsigned(27,8) ,
64938	 => std_logic_vector(to_unsigned(47,8) ,
64939	 => std_logic_vector(to_unsigned(18,8) ,
64940	 => std_logic_vector(to_unsigned(14,8) ,
64941	 => std_logic_vector(to_unsigned(15,8) ,
64942	 => std_logic_vector(to_unsigned(16,8) ,
64943	 => std_logic_vector(to_unsigned(35,8) ,
64944	 => std_logic_vector(to_unsigned(16,8) ,
64945	 => std_logic_vector(to_unsigned(12,8) ,
64946	 => std_logic_vector(to_unsigned(6,8) ,
64947	 => std_logic_vector(to_unsigned(9,8) ,
64948	 => std_logic_vector(to_unsigned(6,8) ,
64949	 => std_logic_vector(to_unsigned(6,8) ,
64950	 => std_logic_vector(to_unsigned(7,8) ,
64951	 => std_logic_vector(to_unsigned(4,8) ,
64952	 => std_logic_vector(to_unsigned(8,8) ,
64953	 => std_logic_vector(to_unsigned(4,8) ,
64954	 => std_logic_vector(to_unsigned(5,8) ,
64955	 => std_logic_vector(to_unsigned(6,8) ,
64956	 => std_logic_vector(to_unsigned(11,8) ,
64957	 => std_logic_vector(to_unsigned(13,8) ,
64958	 => std_logic_vector(to_unsigned(13,8) ,
64959	 => std_logic_vector(to_unsigned(9,8) ,
64960	 => std_logic_vector(to_unsigned(10,8) ,
64961	 => std_logic_vector(to_unsigned(107,8) ,
64962	 => std_logic_vector(to_unsigned(100,8) ,
64963	 => std_logic_vector(to_unsigned(97,8) ,
64964	 => std_logic_vector(to_unsigned(93,8) ,
64965	 => std_logic_vector(to_unsigned(96,8) ,
64966	 => std_logic_vector(to_unsigned(99,8) ,
64967	 => std_logic_vector(to_unsigned(96,8) ,
64968	 => std_logic_vector(to_unsigned(93,8) ,
64969	 => std_logic_vector(to_unsigned(90,8) ,
64970	 => std_logic_vector(to_unsigned(87,8) ,
64971	 => std_logic_vector(to_unsigned(81,8) ,
64972	 => std_logic_vector(to_unsigned(87,8) ,
64973	 => std_logic_vector(to_unsigned(69,8) ,
64974	 => std_logic_vector(to_unsigned(52,8) ,
64975	 => std_logic_vector(to_unsigned(72,8) ,
64976	 => std_logic_vector(to_unsigned(44,8) ,
64977	 => std_logic_vector(to_unsigned(44,8) ,
64978	 => std_logic_vector(to_unsigned(44,8) ,
64979	 => std_logic_vector(to_unsigned(33,8) ,
64980	 => std_logic_vector(to_unsigned(25,8) ,
64981	 => std_logic_vector(to_unsigned(29,8) ,
64982	 => std_logic_vector(to_unsigned(64,8) ,
64983	 => std_logic_vector(to_unsigned(50,8) ,
64984	 => std_logic_vector(to_unsigned(35,8) ,
64985	 => std_logic_vector(to_unsigned(40,8) ,
64986	 => std_logic_vector(to_unsigned(38,8) ,
64987	 => std_logic_vector(to_unsigned(45,8) ,
64988	 => std_logic_vector(to_unsigned(42,8) ,
64989	 => std_logic_vector(to_unsigned(37,8) ,
64990	 => std_logic_vector(to_unsigned(37,8) ,
64991	 => std_logic_vector(to_unsigned(30,8) ,
64992	 => std_logic_vector(to_unsigned(27,8) ,
64993	 => std_logic_vector(to_unsigned(34,8) ,
64994	 => std_logic_vector(to_unsigned(37,8) ,
64995	 => std_logic_vector(to_unsigned(36,8) ,
64996	 => std_logic_vector(to_unsigned(32,8) ,
64997	 => std_logic_vector(to_unsigned(33,8) ,
64998	 => std_logic_vector(to_unsigned(24,8) ,
64999	 => std_logic_vector(to_unsigned(19,8) ,
65000	 => std_logic_vector(to_unsigned(19,8) ,
65001	 => std_logic_vector(to_unsigned(26,8) ,
65002	 => std_logic_vector(to_unsigned(29,8) ,
65003	 => std_logic_vector(to_unsigned(35,8) ,
65004	 => std_logic_vector(to_unsigned(41,8) ,
65005	 => std_logic_vector(to_unsigned(41,8) ,
65006	 => std_logic_vector(to_unsigned(45,8) ,
65007	 => std_logic_vector(to_unsigned(52,8) ,
65008	 => std_logic_vector(to_unsigned(61,8) ,
65009	 => std_logic_vector(to_unsigned(44,8) ,
65010	 => std_logic_vector(to_unsigned(39,8) ,
65011	 => std_logic_vector(to_unsigned(41,8) ,
65012	 => std_logic_vector(to_unsigned(35,8) ,
65013	 => std_logic_vector(to_unsigned(37,8) ,
65014	 => std_logic_vector(to_unsigned(47,8) ,
65015	 => std_logic_vector(to_unsigned(47,8) ,
65016	 => std_logic_vector(to_unsigned(49,8) ,
65017	 => std_logic_vector(to_unsigned(54,8) ,
65018	 => std_logic_vector(to_unsigned(41,8) ,
65019	 => std_logic_vector(to_unsigned(42,8) ,
65020	 => std_logic_vector(to_unsigned(84,8) ,
65021	 => std_logic_vector(to_unsigned(77,8) ,
65022	 => std_logic_vector(to_unsigned(48,8) ,
65023	 => std_logic_vector(to_unsigned(62,8) ,
65024	 => std_logic_vector(to_unsigned(62,8) ,
65025	 => std_logic_vector(to_unsigned(72,8) ,
65026	 => std_logic_vector(to_unsigned(65,8) ,
65027	 => std_logic_vector(to_unsigned(64,8) ,
65028	 => std_logic_vector(to_unsigned(59,8) ,
65029	 => std_logic_vector(to_unsigned(50,8) ,
65030	 => std_logic_vector(to_unsigned(68,8) ,
65031	 => std_logic_vector(to_unsigned(66,8) ,
65032	 => std_logic_vector(to_unsigned(57,8) ,
65033	 => std_logic_vector(to_unsigned(104,8) ,
65034	 => std_logic_vector(to_unsigned(138,8) ,
65035	 => std_logic_vector(to_unsigned(130,8) ,
65036	 => std_logic_vector(to_unsigned(108,8) ,
65037	 => std_logic_vector(to_unsigned(90,8) ,
65038	 => std_logic_vector(to_unsigned(109,8) ,
65039	 => std_logic_vector(to_unsigned(77,8) ,
65040	 => std_logic_vector(to_unsigned(32,8) ,
65041	 => std_logic_vector(to_unsigned(22,8) ,
65042	 => std_logic_vector(to_unsigned(62,8) ,
65043	 => std_logic_vector(to_unsigned(147,8) ,
65044	 => std_logic_vector(to_unsigned(96,8) ,
65045	 => std_logic_vector(to_unsigned(32,8) ,
65046	 => std_logic_vector(to_unsigned(44,8) ,
65047	 => std_logic_vector(to_unsigned(58,8) ,
65048	 => std_logic_vector(to_unsigned(53,8) ,
65049	 => std_logic_vector(to_unsigned(70,8) ,
65050	 => std_logic_vector(to_unsigned(56,8) ,
65051	 => std_logic_vector(to_unsigned(38,8) ,
65052	 => std_logic_vector(to_unsigned(47,8) ,
65053	 => std_logic_vector(to_unsigned(91,8) ,
65054	 => std_logic_vector(to_unsigned(68,8) ,
65055	 => std_logic_vector(to_unsigned(66,8) ,
65056	 => std_logic_vector(to_unsigned(71,8) ,
65057	 => std_logic_vector(to_unsigned(60,8) ,
65058	 => std_logic_vector(to_unsigned(64,8) ,
65059	 => std_logic_vector(to_unsigned(60,8) ,
65060	 => std_logic_vector(to_unsigned(60,8) ,
65061	 => std_logic_vector(to_unsigned(58,8) ,
65062	 => std_logic_vector(to_unsigned(47,8) ,
65063	 => std_logic_vector(to_unsigned(44,8) ,
65064	 => std_logic_vector(to_unsigned(44,8) ,
65065	 => std_logic_vector(to_unsigned(33,8) ,
65066	 => std_logic_vector(to_unsigned(28,8) ,
65067	 => std_logic_vector(to_unsigned(21,8) ,
65068	 => std_logic_vector(to_unsigned(26,8) ,
65069	 => std_logic_vector(to_unsigned(61,8) ,
65070	 => std_logic_vector(to_unsigned(82,8) ,
65071	 => std_logic_vector(to_unsigned(58,8) ,
65072	 => std_logic_vector(to_unsigned(50,8) ,
65073	 => std_logic_vector(to_unsigned(49,8) ,
65074	 => std_logic_vector(to_unsigned(42,8) ,
65075	 => std_logic_vector(to_unsigned(41,8) ,
65076	 => std_logic_vector(to_unsigned(34,8) ,
65077	 => std_logic_vector(to_unsigned(26,8) ,
65078	 => std_logic_vector(to_unsigned(23,8) ,
65079	 => std_logic_vector(to_unsigned(30,8) ,
65080	 => std_logic_vector(to_unsigned(34,8) ,
65081	 => std_logic_vector(to_unsigned(30,8) ,
65082	 => std_logic_vector(to_unsigned(51,8) ,
65083	 => std_logic_vector(to_unsigned(60,8) ,
65084	 => std_logic_vector(to_unsigned(63,8) ,
65085	 => std_logic_vector(to_unsigned(41,8) ,
65086	 => std_logic_vector(to_unsigned(24,8) ,
65087	 => std_logic_vector(to_unsigned(18,8) ,
65088	 => std_logic_vector(to_unsigned(20,8) ,
65089	 => std_logic_vector(to_unsigned(69,8) ,
65090	 => std_logic_vector(to_unsigned(61,8) ,
65091	 => std_logic_vector(to_unsigned(80,8) ,
65092	 => std_logic_vector(to_unsigned(112,8) ,
65093	 => std_logic_vector(to_unsigned(82,8) ,
65094	 => std_logic_vector(to_unsigned(67,8) ,
65095	 => std_logic_vector(to_unsigned(45,8) ,
65096	 => std_logic_vector(to_unsigned(51,8) ,
65097	 => std_logic_vector(to_unsigned(58,8) ,
65098	 => std_logic_vector(to_unsigned(80,8) ,
65099	 => std_logic_vector(to_unsigned(93,8) ,
65100	 => std_logic_vector(to_unsigned(58,8) ,
65101	 => std_logic_vector(to_unsigned(12,8) ,
65102	 => std_logic_vector(to_unsigned(20,8) ,
65103	 => std_logic_vector(to_unsigned(29,8) ,
65104	 => std_logic_vector(to_unsigned(14,8) ,
65105	 => std_logic_vector(to_unsigned(16,8) ,
65106	 => std_logic_vector(to_unsigned(24,8) ,
65107	 => std_logic_vector(to_unsigned(14,8) ,
65108	 => std_logic_vector(to_unsigned(26,8) ,
65109	 => std_logic_vector(to_unsigned(85,8) ,
65110	 => std_logic_vector(to_unsigned(108,8) ,
65111	 => std_logic_vector(to_unsigned(104,8) ,
65112	 => std_logic_vector(to_unsigned(80,8) ,
65113	 => std_logic_vector(to_unsigned(97,8) ,
65114	 => std_logic_vector(to_unsigned(88,8) ,
65115	 => std_logic_vector(to_unsigned(85,8) ,
65116	 => std_logic_vector(to_unsigned(43,8) ,
65117	 => std_logic_vector(to_unsigned(13,8) ,
65118	 => std_logic_vector(to_unsigned(9,8) ,
65119	 => std_logic_vector(to_unsigned(5,8) ,
65120	 => std_logic_vector(to_unsigned(16,8) ,
65121	 => std_logic_vector(to_unsigned(29,8) ,
65122	 => std_logic_vector(to_unsigned(21,8) ,
65123	 => std_logic_vector(to_unsigned(22,8) ,
65124	 => std_logic_vector(to_unsigned(36,8) ,
65125	 => std_logic_vector(to_unsigned(23,8) ,
65126	 => std_logic_vector(to_unsigned(11,8) ,
65127	 => std_logic_vector(to_unsigned(8,8) ,
65128	 => std_logic_vector(to_unsigned(18,8) ,
65129	 => std_logic_vector(to_unsigned(58,8) ,
65130	 => std_logic_vector(to_unsigned(40,8) ,
65131	 => std_logic_vector(to_unsigned(29,8) ,
65132	 => std_logic_vector(to_unsigned(23,8) ,
65133	 => std_logic_vector(to_unsigned(20,8) ,
65134	 => std_logic_vector(to_unsigned(36,8) ,
65135	 => std_logic_vector(to_unsigned(26,8) ,
65136	 => std_logic_vector(to_unsigned(33,8) ,
65137	 => std_logic_vector(to_unsigned(63,8) ,
65138	 => std_logic_vector(to_unsigned(41,8) ,
65139	 => std_logic_vector(to_unsigned(32,8) ,
65140	 => std_logic_vector(to_unsigned(34,8) ,
65141	 => std_logic_vector(to_unsigned(12,8) ,
65142	 => std_logic_vector(to_unsigned(9,8) ,
65143	 => std_logic_vector(to_unsigned(11,8) ,
65144	 => std_logic_vector(to_unsigned(11,8) ,
65145	 => std_logic_vector(to_unsigned(24,8) ,
65146	 => std_logic_vector(to_unsigned(44,8) ,
65147	 => std_logic_vector(to_unsigned(25,8) ,
65148	 => std_logic_vector(to_unsigned(22,8) ,
65149	 => std_logic_vector(to_unsigned(32,8) ,
65150	 => std_logic_vector(to_unsigned(49,8) ,
65151	 => std_logic_vector(to_unsigned(49,8) ,
65152	 => std_logic_vector(to_unsigned(58,8) ,
65153	 => std_logic_vector(to_unsigned(63,8) ,
65154	 => std_logic_vector(to_unsigned(62,8) ,
65155	 => std_logic_vector(to_unsigned(54,8) ,
65156	 => std_logic_vector(to_unsigned(53,8) ,
65157	 => std_logic_vector(to_unsigned(50,8) ,
65158	 => std_logic_vector(to_unsigned(50,8) ,
65159	 => std_logic_vector(to_unsigned(37,8) ,
65160	 => std_logic_vector(to_unsigned(45,8) ,
65161	 => std_logic_vector(to_unsigned(43,8) ,
65162	 => std_logic_vector(to_unsigned(17,8) ,
65163	 => std_logic_vector(to_unsigned(10,8) ,
65164	 => std_logic_vector(to_unsigned(29,8) ,
65165	 => std_logic_vector(to_unsigned(53,8) ,
65166	 => std_logic_vector(to_unsigned(30,8) ,
65167	 => std_logic_vector(to_unsigned(13,8) ,
65168	 => std_logic_vector(to_unsigned(37,8) ,
65169	 => std_logic_vector(to_unsigned(19,8) ,
65170	 => std_logic_vector(to_unsigned(25,8) ,
65171	 => std_logic_vector(to_unsigned(23,8) ,
65172	 => std_logic_vector(to_unsigned(24,8) ,
65173	 => std_logic_vector(to_unsigned(34,8) ,
65174	 => std_logic_vector(to_unsigned(39,8) ,
65175	 => std_logic_vector(to_unsigned(42,8) ,
65176	 => std_logic_vector(to_unsigned(36,8) ,
65177	 => std_logic_vector(to_unsigned(37,8) ,
65178	 => std_logic_vector(to_unsigned(31,8) ,
65179	 => std_logic_vector(to_unsigned(22,8) ,
65180	 => std_logic_vector(to_unsigned(24,8) ,
65181	 => std_logic_vector(to_unsigned(25,8) ,
65182	 => std_logic_vector(to_unsigned(22,8) ,
65183	 => std_logic_vector(to_unsigned(58,8) ,
65184	 => std_logic_vector(to_unsigned(61,8) ,
65185	 => std_logic_vector(to_unsigned(45,8) ,
65186	 => std_logic_vector(to_unsigned(44,8) ,
65187	 => std_logic_vector(to_unsigned(30,8) ,
65188	 => std_logic_vector(to_unsigned(25,8) ,
65189	 => std_logic_vector(to_unsigned(72,8) ,
65190	 => std_logic_vector(to_unsigned(131,8) ,
65191	 => std_logic_vector(to_unsigned(93,8) ,
65192	 => std_logic_vector(to_unsigned(25,8) ,
65193	 => std_logic_vector(to_unsigned(25,8) ,
65194	 => std_logic_vector(to_unsigned(37,8) ,
65195	 => std_logic_vector(to_unsigned(44,8) ,
65196	 => std_logic_vector(to_unsigned(36,8) ,
65197	 => std_logic_vector(to_unsigned(88,8) ,
65198	 => std_logic_vector(to_unsigned(63,8) ,
65199	 => std_logic_vector(to_unsigned(8,8) ,
65200	 => std_logic_vector(to_unsigned(13,8) ,
65201	 => std_logic_vector(to_unsigned(40,8) ,
65202	 => std_logic_vector(to_unsigned(41,8) ,
65203	 => std_logic_vector(to_unsigned(48,8) ,
65204	 => std_logic_vector(to_unsigned(42,8) ,
65205	 => std_logic_vector(to_unsigned(39,8) ,
65206	 => std_logic_vector(to_unsigned(26,8) ,
65207	 => std_logic_vector(to_unsigned(11,8) ,
65208	 => std_logic_vector(to_unsigned(16,8) ,
65209	 => std_logic_vector(to_unsigned(26,8) ,
65210	 => std_logic_vector(to_unsigned(42,8) ,
65211	 => std_logic_vector(to_unsigned(24,8) ,
65212	 => std_logic_vector(to_unsigned(25,8) ,
65213	 => std_logic_vector(to_unsigned(49,8) ,
65214	 => std_logic_vector(to_unsigned(35,8) ,
65215	 => std_logic_vector(to_unsigned(19,8) ,
65216	 => std_logic_vector(to_unsigned(27,8) ,
65217	 => std_logic_vector(to_unsigned(31,8) ,
65218	 => std_logic_vector(to_unsigned(34,8) ,
65219	 => std_logic_vector(to_unsigned(27,8) ,
65220	 => std_logic_vector(to_unsigned(18,8) ,
65221	 => std_logic_vector(to_unsigned(16,8) ,
65222	 => std_logic_vector(to_unsigned(20,8) ,
65223	 => std_logic_vector(to_unsigned(24,8) ,
65224	 => std_logic_vector(to_unsigned(26,8) ,
65225	 => std_logic_vector(to_unsigned(24,8) ,
65226	 => std_logic_vector(to_unsigned(23,8) ,
65227	 => std_logic_vector(to_unsigned(20,8) ,
65228	 => std_logic_vector(to_unsigned(25,8) ,
65229	 => std_logic_vector(to_unsigned(19,8) ,
65230	 => std_logic_vector(to_unsigned(10,8) ,
65231	 => std_logic_vector(to_unsigned(2,8) ,
65232	 => std_logic_vector(to_unsigned(0,8) ,
65233	 => std_logic_vector(to_unsigned(3,8) ,
65234	 => std_logic_vector(to_unsigned(17,8) ,
65235	 => std_logic_vector(to_unsigned(24,8) ,
65236	 => std_logic_vector(to_unsigned(29,8) ,
65237	 => std_logic_vector(to_unsigned(30,8) ,
65238	 => std_logic_vector(to_unsigned(29,8) ,
65239	 => std_logic_vector(to_unsigned(24,8) ,
65240	 => std_logic_vector(to_unsigned(19,8) ,
65241	 => std_logic_vector(to_unsigned(24,8) ,
65242	 => std_logic_vector(to_unsigned(19,8) ,
65243	 => std_logic_vector(to_unsigned(18,8) ,
65244	 => std_logic_vector(to_unsigned(12,8) ,
65245	 => std_logic_vector(to_unsigned(0,8) ,
65246	 => std_logic_vector(to_unsigned(0,8) ,
65247	 => std_logic_vector(to_unsigned(4,8) ,
65248	 => std_logic_vector(to_unsigned(10,8) ,
65249	 => std_logic_vector(to_unsigned(14,8) ,
65250	 => std_logic_vector(to_unsigned(12,8) ,
65251	 => std_logic_vector(to_unsigned(12,8) ,
65252	 => std_logic_vector(to_unsigned(17,8) ,
65253	 => std_logic_vector(to_unsigned(17,8) ,
65254	 => std_logic_vector(to_unsigned(5,8) ,
65255	 => std_logic_vector(to_unsigned(1,8) ,
65256	 => std_logic_vector(to_unsigned(0,8) ,
65257	 => std_logic_vector(to_unsigned(5,8) ,
65258	 => std_logic_vector(to_unsigned(29,8) ,
65259	 => std_logic_vector(to_unsigned(23,8) ,
65260	 => std_logic_vector(to_unsigned(21,8) ,
65261	 => std_logic_vector(to_unsigned(24,8) ,
65262	 => std_logic_vector(to_unsigned(25,8) ,
65263	 => std_logic_vector(to_unsigned(33,8) ,
65264	 => std_logic_vector(to_unsigned(18,8) ,
65265	 => std_logic_vector(to_unsigned(15,8) ,
65266	 => std_logic_vector(to_unsigned(14,8) ,
65267	 => std_logic_vector(to_unsigned(11,8) ,
65268	 => std_logic_vector(to_unsigned(8,8) ,
65269	 => std_logic_vector(to_unsigned(12,8) ,
65270	 => std_logic_vector(to_unsigned(27,8) ,
65271	 => std_logic_vector(to_unsigned(8,8) ,
65272	 => std_logic_vector(to_unsigned(10,8) ,
65273	 => std_logic_vector(to_unsigned(9,8) ,
65274	 => std_logic_vector(to_unsigned(10,8) ,
65275	 => std_logic_vector(to_unsigned(8,8) ,
65276	 => std_logic_vector(to_unsigned(8,8) ,
65277	 => std_logic_vector(to_unsigned(5,8) ,
65278	 => std_logic_vector(to_unsigned(15,8) ,
65279	 => std_logic_vector(to_unsigned(19,8) ,
65280	 => std_logic_vector(to_unsigned(6,8) ,
65281	 => std_logic_vector(to_unsigned(104,8) ,
65282	 => std_logic_vector(to_unsigned(95,8) ,
65283	 => std_logic_vector(to_unsigned(95,8) ,
65284	 => std_logic_vector(to_unsigned(84,8) ,
65285	 => std_logic_vector(to_unsigned(105,8) ,
65286	 => std_logic_vector(to_unsigned(108,8) ,
65287	 => std_logic_vector(to_unsigned(91,8) ,
65288	 => std_logic_vector(to_unsigned(95,8) ,
65289	 => std_logic_vector(to_unsigned(97,8) ,
65290	 => std_logic_vector(to_unsigned(88,8) ,
65291	 => std_logic_vector(to_unsigned(84,8) ,
65292	 => std_logic_vector(to_unsigned(86,8) ,
65293	 => std_logic_vector(to_unsigned(54,8) ,
65294	 => std_logic_vector(to_unsigned(43,8) ,
65295	 => std_logic_vector(to_unsigned(72,8) ,
65296	 => std_logic_vector(to_unsigned(68,8) ,
65297	 => std_logic_vector(to_unsigned(73,8) ,
65298	 => std_logic_vector(to_unsigned(81,8) ,
65299	 => std_logic_vector(to_unsigned(58,8) ,
65300	 => std_logic_vector(to_unsigned(51,8) ,
65301	 => std_logic_vector(to_unsigned(64,8) ,
65302	 => std_logic_vector(to_unsigned(95,8) ,
65303	 => std_logic_vector(to_unsigned(72,8) ,
65304	 => std_logic_vector(to_unsigned(35,8) ,
65305	 => std_logic_vector(to_unsigned(35,8) ,
65306	 => std_logic_vector(to_unsigned(41,8) ,
65307	 => std_logic_vector(to_unsigned(45,8) ,
65308	 => std_logic_vector(to_unsigned(42,8) ,
65309	 => std_logic_vector(to_unsigned(37,8) ,
65310	 => std_logic_vector(to_unsigned(31,8) ,
65311	 => std_logic_vector(to_unsigned(31,8) ,
65312	 => std_logic_vector(to_unsigned(32,8) ,
65313	 => std_logic_vector(to_unsigned(36,8) ,
65314	 => std_logic_vector(to_unsigned(32,8) ,
65315	 => std_logic_vector(to_unsigned(30,8) ,
65316	 => std_logic_vector(to_unsigned(29,8) ,
65317	 => std_logic_vector(to_unsigned(35,8) ,
65318	 => std_logic_vector(to_unsigned(27,8) ,
65319	 => std_logic_vector(to_unsigned(13,8) ,
65320	 => std_logic_vector(to_unsigned(23,8) ,
65321	 => std_logic_vector(to_unsigned(32,8) ,
65322	 => std_logic_vector(to_unsigned(24,8) ,
65323	 => std_logic_vector(to_unsigned(27,8) ,
65324	 => std_logic_vector(to_unsigned(31,8) ,
65325	 => std_logic_vector(to_unsigned(37,8) ,
65326	 => std_logic_vector(to_unsigned(40,8) ,
65327	 => std_logic_vector(to_unsigned(45,8) ,
65328	 => std_logic_vector(to_unsigned(56,8) ,
65329	 => std_logic_vector(to_unsigned(43,8) ,
65330	 => std_logic_vector(to_unsigned(35,8) ,
65331	 => std_logic_vector(to_unsigned(48,8) ,
65332	 => std_logic_vector(to_unsigned(32,8) ,
65333	 => std_logic_vector(to_unsigned(20,8) ,
65334	 => std_logic_vector(to_unsigned(46,8) ,
65335	 => std_logic_vector(to_unsigned(46,8) ,
65336	 => std_logic_vector(to_unsigned(47,8) ,
65337	 => std_logic_vector(to_unsigned(44,8) ,
65338	 => std_logic_vector(to_unsigned(49,8) ,
65339	 => std_logic_vector(to_unsigned(65,8) ,
65340	 => std_logic_vector(to_unsigned(93,8) ,
65341	 => std_logic_vector(to_unsigned(85,8) ,
65342	 => std_logic_vector(to_unsigned(67,8) ,
65343	 => std_logic_vector(to_unsigned(71,8) ,
65344	 => std_logic_vector(to_unsigned(93,8) ,
65345	 => std_logic_vector(to_unsigned(95,8) ,
65346	 => std_logic_vector(to_unsigned(92,8) ,
65347	 => std_logic_vector(to_unsigned(96,8) ,
65348	 => std_logic_vector(to_unsigned(93,8) ,
65349	 => std_logic_vector(to_unsigned(92,8) ,
65350	 => std_logic_vector(to_unsigned(86,8) ,
65351	 => std_logic_vector(to_unsigned(78,8) ,
65352	 => std_logic_vector(to_unsigned(88,8) ,
65353	 => std_logic_vector(to_unsigned(107,8) ,
65354	 => std_logic_vector(to_unsigned(121,8) ,
65355	 => std_logic_vector(to_unsigned(121,8) ,
65356	 => std_logic_vector(to_unsigned(93,8) ,
65357	 => std_logic_vector(to_unsigned(86,8) ,
65358	 => std_logic_vector(to_unsigned(108,8) ,
65359	 => std_logic_vector(to_unsigned(101,8) ,
65360	 => std_logic_vector(to_unsigned(78,8) ,
65361	 => std_logic_vector(to_unsigned(62,8) ,
65362	 => std_logic_vector(to_unsigned(79,8) ,
65363	 => std_logic_vector(to_unsigned(125,8) ,
65364	 => std_logic_vector(to_unsigned(96,8) ,
65365	 => std_logic_vector(to_unsigned(30,8) ,
65366	 => std_logic_vector(to_unsigned(41,8) ,
65367	 => std_logic_vector(to_unsigned(60,8) ,
65368	 => std_logic_vector(to_unsigned(79,8) ,
65369	 => std_logic_vector(to_unsigned(58,8) ,
65370	 => std_logic_vector(to_unsigned(24,8) ,
65371	 => std_logic_vector(to_unsigned(39,8) ,
65372	 => std_logic_vector(to_unsigned(71,8) ,
65373	 => std_logic_vector(to_unsigned(86,8) ,
65374	 => std_logic_vector(to_unsigned(58,8) ,
65375	 => std_logic_vector(to_unsigned(81,8) ,
65376	 => std_logic_vector(to_unsigned(79,8) ,
65377	 => std_logic_vector(to_unsigned(41,8) ,
65378	 => std_logic_vector(to_unsigned(31,8) ,
65379	 => std_logic_vector(to_unsigned(47,8) ,
65380	 => std_logic_vector(to_unsigned(37,8) ,
65381	 => std_logic_vector(to_unsigned(42,8) ,
65382	 => std_logic_vector(to_unsigned(43,8) ,
65383	 => std_logic_vector(to_unsigned(37,8) ,
65384	 => std_logic_vector(to_unsigned(32,8) ,
65385	 => std_logic_vector(to_unsigned(28,8) ,
65386	 => std_logic_vector(to_unsigned(25,8) ,
65387	 => std_logic_vector(to_unsigned(22,8) ,
65388	 => std_logic_vector(to_unsigned(23,8) ,
65389	 => std_logic_vector(to_unsigned(56,8) ,
65390	 => std_logic_vector(to_unsigned(112,8) ,
65391	 => std_logic_vector(to_unsigned(69,8) ,
65392	 => std_logic_vector(to_unsigned(54,8) ,
65393	 => std_logic_vector(to_unsigned(108,8) ,
65394	 => std_logic_vector(to_unsigned(90,8) ,
65395	 => std_logic_vector(to_unsigned(57,8) ,
65396	 => std_logic_vector(to_unsigned(43,8) ,
65397	 => std_logic_vector(to_unsigned(43,8) ,
65398	 => std_logic_vector(to_unsigned(42,8) ,
65399	 => std_logic_vector(to_unsigned(40,8) ,
65400	 => std_logic_vector(to_unsigned(35,8) ,
65401	 => std_logic_vector(to_unsigned(47,8) ,
65402	 => std_logic_vector(to_unsigned(41,8) ,
65403	 => std_logic_vector(to_unsigned(26,8) ,
65404	 => std_logic_vector(to_unsigned(16,8) ,
65405	 => std_logic_vector(to_unsigned(16,8) ,
65406	 => std_logic_vector(to_unsigned(25,8) ,
65407	 => std_logic_vector(to_unsigned(17,8) ,
65408	 => std_logic_vector(to_unsigned(32,8) ,
65409	 => std_logic_vector(to_unsigned(146,8) ,
65410	 => std_logic_vector(to_unsigned(136,8) ,
65411	 => std_logic_vector(to_unsigned(141,8) ,
65412	 => std_logic_vector(to_unsigned(177,8) ,
65413	 => std_logic_vector(to_unsigned(103,8) ,
65414	 => std_logic_vector(to_unsigned(48,8) ,
65415	 => std_logic_vector(to_unsigned(32,8) ,
65416	 => std_logic_vector(to_unsigned(40,8) ,
65417	 => std_logic_vector(to_unsigned(28,8) ,
65418	 => std_logic_vector(to_unsigned(64,8) ,
65419	 => std_logic_vector(to_unsigned(67,8) ,
65420	 => std_logic_vector(to_unsigned(24,8) ,
65421	 => std_logic_vector(to_unsigned(19,8) ,
65422	 => std_logic_vector(to_unsigned(22,8) ,
65423	 => std_logic_vector(to_unsigned(24,8) ,
65424	 => std_logic_vector(to_unsigned(12,8) ,
65425	 => std_logic_vector(to_unsigned(10,8) ,
65426	 => std_logic_vector(to_unsigned(20,8) ,
65427	 => std_logic_vector(to_unsigned(20,8) ,
65428	 => std_logic_vector(to_unsigned(30,8) ,
65429	 => std_logic_vector(to_unsigned(88,8) ,
65430	 => std_logic_vector(to_unsigned(93,8) ,
65431	 => std_logic_vector(to_unsigned(81,8) ,
65432	 => std_logic_vector(to_unsigned(72,8) ,
65433	 => std_logic_vector(to_unsigned(119,8) ,
65434	 => std_logic_vector(to_unsigned(90,8) ,
65435	 => std_logic_vector(to_unsigned(72,8) ,
65436	 => std_logic_vector(to_unsigned(42,8) ,
65437	 => std_logic_vector(to_unsigned(12,8) ,
65438	 => std_logic_vector(to_unsigned(8,8) ,
65439	 => std_logic_vector(to_unsigned(4,8) ,
65440	 => std_logic_vector(to_unsigned(15,8) ,
65441	 => std_logic_vector(to_unsigned(40,8) ,
65442	 => std_logic_vector(to_unsigned(24,8) ,
65443	 => std_logic_vector(to_unsigned(31,8) ,
65444	 => std_logic_vector(to_unsigned(36,8) ,
65445	 => std_logic_vector(to_unsigned(25,8) ,
65446	 => std_logic_vector(to_unsigned(18,8) ,
65447	 => std_logic_vector(to_unsigned(17,8) ,
65448	 => std_logic_vector(to_unsigned(27,8) ,
65449	 => std_logic_vector(to_unsigned(50,8) ,
65450	 => std_logic_vector(to_unsigned(37,8) ,
65451	 => std_logic_vector(to_unsigned(40,8) ,
65452	 => std_logic_vector(to_unsigned(40,8) ,
65453	 => std_logic_vector(to_unsigned(29,8) ,
65454	 => std_logic_vector(to_unsigned(22,8) ,
65455	 => std_logic_vector(to_unsigned(29,8) ,
65456	 => std_logic_vector(to_unsigned(56,8) ,
65457	 => std_logic_vector(to_unsigned(27,8) ,
65458	 => std_logic_vector(to_unsigned(24,8) ,
65459	 => std_logic_vector(to_unsigned(38,8) ,
65460	 => std_logic_vector(to_unsigned(18,8) ,
65461	 => std_logic_vector(to_unsigned(8,8) ,
65462	 => std_logic_vector(to_unsigned(7,8) ,
65463	 => std_logic_vector(to_unsigned(8,8) ,
65464	 => std_logic_vector(to_unsigned(10,8) ,
65465	 => std_logic_vector(to_unsigned(15,8) ,
65466	 => std_logic_vector(to_unsigned(41,8) ,
65467	 => std_logic_vector(to_unsigned(41,8) ,
65468	 => std_logic_vector(to_unsigned(36,8) ,
65469	 => std_logic_vector(to_unsigned(35,8) ,
65470	 => std_logic_vector(to_unsigned(44,8) ,
65471	 => std_logic_vector(to_unsigned(51,8) ,
65472	 => std_logic_vector(to_unsigned(32,8) ,
65473	 => std_logic_vector(to_unsigned(23,8) ,
65474	 => std_logic_vector(to_unsigned(35,8) ,
65475	 => std_logic_vector(to_unsigned(52,8) ,
65476	 => std_logic_vector(to_unsigned(47,8) ,
65477	 => std_logic_vector(to_unsigned(45,8) ,
65478	 => std_logic_vector(to_unsigned(43,8) ,
65479	 => std_logic_vector(to_unsigned(53,8) ,
65480	 => std_logic_vector(to_unsigned(51,8) ,
65481	 => std_logic_vector(to_unsigned(30,8) ,
65482	 => std_logic_vector(to_unsigned(18,8) ,
65483	 => std_logic_vector(to_unsigned(20,8) ,
65484	 => std_logic_vector(to_unsigned(18,8) ,
65485	 => std_logic_vector(to_unsigned(23,8) ,
65486	 => std_logic_vector(to_unsigned(17,8) ,
65487	 => std_logic_vector(to_unsigned(14,8) ,
65488	 => std_logic_vector(to_unsigned(35,8) ,
65489	 => std_logic_vector(to_unsigned(19,8) ,
65490	 => std_logic_vector(to_unsigned(23,8) ,
65491	 => std_logic_vector(to_unsigned(20,8) ,
65492	 => std_logic_vector(to_unsigned(27,8) ,
65493	 => std_logic_vector(to_unsigned(37,8) ,
65494	 => std_logic_vector(to_unsigned(37,8) ,
65495	 => std_logic_vector(to_unsigned(37,8) ,
65496	 => std_logic_vector(to_unsigned(47,8) ,
65497	 => std_logic_vector(to_unsigned(46,8) ,
65498	 => std_logic_vector(to_unsigned(38,8) ,
65499	 => std_logic_vector(to_unsigned(23,8) ,
65500	 => std_logic_vector(to_unsigned(17,8) ,
65501	 => std_logic_vector(to_unsigned(21,8) ,
65502	 => std_logic_vector(to_unsigned(20,8) ,
65503	 => std_logic_vector(to_unsigned(41,8) ,
65504	 => std_logic_vector(to_unsigned(44,8) ,
65505	 => std_logic_vector(to_unsigned(41,8) ,
65506	 => std_logic_vector(to_unsigned(46,8) ,
65507	 => std_logic_vector(to_unsigned(29,8) ,
65508	 => std_logic_vector(to_unsigned(25,8) ,
65509	 => std_logic_vector(to_unsigned(19,8) ,
65510	 => std_logic_vector(to_unsigned(51,8) ,
65511	 => std_logic_vector(to_unsigned(86,8) ,
65512	 => std_logic_vector(to_unsigned(37,8) ,
65513	 => std_logic_vector(to_unsigned(20,8) ,
65514	 => std_logic_vector(to_unsigned(20,8) ,
65515	 => std_logic_vector(to_unsigned(33,8) ,
65516	 => std_logic_vector(to_unsigned(45,8) ,
65517	 => std_logic_vector(to_unsigned(88,8) ,
65518	 => std_logic_vector(to_unsigned(63,8) ,
65519	 => std_logic_vector(to_unsigned(17,8) ,
65520	 => std_logic_vector(to_unsigned(49,8) ,
65521	 => std_logic_vector(to_unsigned(63,8) ,
65522	 => std_logic_vector(to_unsigned(57,8) ,
65523	 => std_logic_vector(to_unsigned(72,8) ,
65524	 => std_logic_vector(to_unsigned(51,8) ,
65525	 => std_logic_vector(to_unsigned(52,8) ,
65526	 => std_logic_vector(to_unsigned(31,8) ,
65527	 => std_logic_vector(to_unsigned(9,8) ,
65528	 => std_logic_vector(to_unsigned(35,8) ,
65529	 => std_logic_vector(to_unsigned(71,8) ,
65530	 => std_logic_vector(to_unsigned(63,8) ,
65531	 => std_logic_vector(to_unsigned(15,8) ,
65532	 => std_logic_vector(to_unsigned(12,8) ,
65533	 => std_logic_vector(to_unsigned(16,8) ,
65534	 => std_logic_vector(to_unsigned(15,8) ,
65535	 => std_logic_vector(to_unsigned(16,8) ,
65536	 => std_logic_vector(to_unsigned(20,8) ,
65537	 => std_logic_vector(to_unsigned(25,8) ,
65538	 => std_logic_vector(to_unsigned(23,8) ,
65539	 => std_logic_vector(to_unsigned(25,8) ,
65540	 => std_logic_vector(to_unsigned(24,8) ,
65541	 => std_logic_vector(to_unsigned(20,8) ,
65542	 => std_logic_vector(to_unsigned(29,8) ,
65543	 => std_logic_vector(to_unsigned(31,8) ,
65544	 => std_logic_vector(to_unsigned(20,8) ,
65545	 => std_logic_vector(to_unsigned(16,8) ,
65546	 => std_logic_vector(to_unsigned(32,8) ,
65547	 => std_logic_vector(to_unsigned(37,8) ,
65548	 => std_logic_vector(to_unsigned(36,8) ,
65549	 => std_logic_vector(to_unsigned(19,8) ,
65550	 => std_logic_vector(to_unsigned(27,8) ,
65551	 => std_logic_vector(to_unsigned(8,8) ,
65552	 => std_logic_vector(to_unsigned(0,8) ,
65553	 => std_logic_vector(to_unsigned(2,8) ,
65554	 => std_logic_vector(to_unsigned(17,8) ,
65555	 => std_logic_vector(to_unsigned(22,8) ,
65556	 => std_logic_vector(to_unsigned(25,8) ,
65557	 => std_logic_vector(to_unsigned(25,8) ,
65558	 => std_logic_vector(to_unsigned(29,8) ,
65559	 => std_logic_vector(to_unsigned(31,8) ,
65560	 => std_logic_vector(to_unsigned(20,8) ,
65561	 => std_logic_vector(to_unsigned(28,8) ,
65562	 => std_logic_vector(to_unsigned(30,8) ,
65563	 => std_logic_vector(to_unsigned(24,8) ,
65564	 => std_logic_vector(to_unsigned(13,8) ,
65565	 => std_logic_vector(to_unsigned(1,8) ,
65566	 => std_logic_vector(to_unsigned(0,8) ,
65567	 => std_logic_vector(to_unsigned(5,8) ,
65568	 => std_logic_vector(to_unsigned(10,8) ,
65569	 => std_logic_vector(to_unsigned(13,8) ,
65570	 => std_logic_vector(to_unsigned(29,8) ,
65571	 => std_logic_vector(to_unsigned(35,8) ,
65572	 => std_logic_vector(to_unsigned(30,8) ,
65573	 => std_logic_vector(to_unsigned(22,8) ,
65574	 => std_logic_vector(to_unsigned(12,8) ,
65575	 => std_logic_vector(to_unsigned(1,8) ,
65576	 => std_logic_vector(to_unsigned(0,8) ,
65577	 => std_logic_vector(to_unsigned(1,8) ,
65578	 => std_logic_vector(to_unsigned(14,8) ,
65579	 => std_logic_vector(to_unsigned(23,8) ,
65580	 => std_logic_vector(to_unsigned(24,8) ,
65581	 => std_logic_vector(to_unsigned(23,8) ,
65582	 => std_logic_vector(to_unsigned(14,8) ,
65583	 => std_logic_vector(to_unsigned(12,8) ,
65584	 => std_logic_vector(to_unsigned(17,8) ,
65585	 => std_logic_vector(to_unsigned(31,8) ,
65586	 => std_logic_vector(to_unsigned(27,8) ,
65587	 => std_logic_vector(to_unsigned(22,8) ,
65588	 => std_logic_vector(to_unsigned(21,8) ,
65589	 => std_logic_vector(to_unsigned(19,8) ,
65590	 => std_logic_vector(to_unsigned(25,8) ,
65591	 => std_logic_vector(to_unsigned(21,8) ,
65592	 => std_logic_vector(to_unsigned(20,8) ,
65593	 => std_logic_vector(to_unsigned(18,8) ,
65594	 => std_logic_vector(to_unsigned(17,8) ,
65595	 => std_logic_vector(to_unsigned(15,8) ,
65596	 => std_logic_vector(to_unsigned(17,8) ,
65597	 => std_logic_vector(to_unsigned(16,8) ,
65598	 => std_logic_vector(to_unsigned(22,8) ,
65599	 => std_logic_vector(to_unsigned(21,8) ,
65600	 => std_logic_vector(to_unsigned(2,8) ,
65601	 => std_logic_vector(to_unsigned(116,8) ,
65602	 => std_logic_vector(to_unsigned(92,8) ,
65603	 => std_logic_vector(to_unsigned(97,8) ,
65604	 => std_logic_vector(to_unsigned(80,8) ,
65605	 => std_logic_vector(to_unsigned(101,8) ,
65606	 => std_logic_vector(to_unsigned(114,8) ,
65607	 => std_logic_vector(to_unsigned(96,8) ,
65608	 => std_logic_vector(to_unsigned(100,8) ,
65609	 => std_logic_vector(to_unsigned(99,8) ,
65610	 => std_logic_vector(to_unsigned(96,8) ,
65611	 => std_logic_vector(to_unsigned(88,8) ,
65612	 => std_logic_vector(to_unsigned(59,8) ,
65613	 => std_logic_vector(to_unsigned(39,8) ,
65614	 => std_logic_vector(to_unsigned(33,8) ,
65615	 => std_logic_vector(to_unsigned(49,8) ,
65616	 => std_logic_vector(to_unsigned(73,8) ,
65617	 => std_logic_vector(to_unsigned(70,8) ,
65618	 => std_logic_vector(to_unsigned(66,8) ,
65619	 => std_logic_vector(to_unsigned(77,8) ,
65620	 => std_logic_vector(to_unsigned(88,8) ,
65621	 => std_logic_vector(to_unsigned(100,8) ,
65622	 => std_logic_vector(to_unsigned(108,8) ,
65623	 => std_logic_vector(to_unsigned(76,8) ,
65624	 => std_logic_vector(to_unsigned(36,8) ,
65625	 => std_logic_vector(to_unsigned(40,8) ,
65626	 => std_logic_vector(to_unsigned(38,8) ,
65627	 => std_logic_vector(to_unsigned(37,8) ,
65628	 => std_logic_vector(to_unsigned(33,8) ,
65629	 => std_logic_vector(to_unsigned(32,8) ,
65630	 => std_logic_vector(to_unsigned(37,8) ,
65631	 => std_logic_vector(to_unsigned(37,8) ,
65632	 => std_logic_vector(to_unsigned(33,8) ,
65633	 => std_logic_vector(to_unsigned(30,8) ,
65634	 => std_logic_vector(to_unsigned(31,8) ,
65635	 => std_logic_vector(to_unsigned(35,8) ,
65636	 => std_logic_vector(to_unsigned(33,8) ,
65637	 => std_logic_vector(to_unsigned(32,8) ,
65638	 => std_logic_vector(to_unsigned(24,8) ,
65639	 => std_logic_vector(to_unsigned(16,8) ,
65640	 => std_logic_vector(to_unsigned(24,8) ,
65641	 => std_logic_vector(to_unsigned(27,8) ,
65642	 => std_logic_vector(to_unsigned(24,8) ,
65643	 => std_logic_vector(to_unsigned(29,8) ,
65644	 => std_logic_vector(to_unsigned(37,8) ,
65645	 => std_logic_vector(to_unsigned(41,8) ,
65646	 => std_logic_vector(to_unsigned(41,8) ,
65647	 => std_logic_vector(to_unsigned(52,8) ,
65648	 => std_logic_vector(to_unsigned(52,8) ,
65649	 => std_logic_vector(to_unsigned(39,8) ,
65650	 => std_logic_vector(to_unsigned(41,8) ,
65651	 => std_logic_vector(to_unsigned(47,8) ,
65652	 => std_logic_vector(to_unsigned(48,8) ,
65653	 => std_logic_vector(to_unsigned(26,8) ,
65654	 => std_logic_vector(to_unsigned(37,8) ,
65655	 => std_logic_vector(to_unsigned(39,8) ,
65656	 => std_logic_vector(to_unsigned(42,8) ,
65657	 => std_logic_vector(to_unsigned(55,8) ,
65658	 => std_logic_vector(to_unsigned(79,8) ,
65659	 => std_logic_vector(to_unsigned(95,8) ,
65660	 => std_logic_vector(to_unsigned(88,8) ,
65661	 => std_logic_vector(to_unsigned(78,8) ,
65662	 => std_logic_vector(to_unsigned(91,8) ,
65663	 => std_logic_vector(to_unsigned(91,8) ,
65664	 => std_logic_vector(to_unsigned(86,8) ,
65665	 => std_logic_vector(to_unsigned(90,8) ,
65666	 => std_logic_vector(to_unsigned(90,8) ,
65667	 => std_logic_vector(to_unsigned(101,8) ,
65668	 => std_logic_vector(to_unsigned(109,8) ,
65669	 => std_logic_vector(to_unsigned(109,8) ,
65670	 => std_logic_vector(to_unsigned(114,8) ,
65671	 => std_logic_vector(to_unsigned(101,8) ,
65672	 => std_logic_vector(to_unsigned(104,8) ,
65673	 => std_logic_vector(to_unsigned(103,8) ,
65674	 => std_logic_vector(to_unsigned(109,8) ,
65675	 => std_logic_vector(to_unsigned(104,8) ,
65676	 => std_logic_vector(to_unsigned(92,8) ,
65677	 => std_logic_vector(to_unsigned(88,8) ,
65678	 => std_logic_vector(to_unsigned(96,8) ,
65679	 => std_logic_vector(to_unsigned(96,8) ,
65680	 => std_logic_vector(to_unsigned(99,8) ,
65681	 => std_logic_vector(to_unsigned(109,8) ,
65682	 => std_logic_vector(to_unsigned(105,8) ,
65683	 => std_logic_vector(to_unsigned(95,8) ,
65684	 => std_logic_vector(to_unsigned(85,8) ,
65685	 => std_logic_vector(to_unsigned(57,8) ,
65686	 => std_logic_vector(to_unsigned(65,8) ,
65687	 => std_logic_vector(to_unsigned(77,8) ,
65688	 => std_logic_vector(to_unsigned(59,8) ,
65689	 => std_logic_vector(to_unsigned(25,8) ,
65690	 => std_logic_vector(to_unsigned(18,8) ,
65691	 => std_logic_vector(to_unsigned(40,8) ,
65692	 => std_logic_vector(to_unsigned(51,8) ,
65693	 => std_logic_vector(to_unsigned(55,8) ,
65694	 => std_logic_vector(to_unsigned(54,8) ,
65695	 => std_logic_vector(to_unsigned(57,8) ,
65696	 => std_logic_vector(to_unsigned(55,8) ,
65697	 => std_logic_vector(to_unsigned(49,8) ,
65698	 => std_logic_vector(to_unsigned(47,8) ,
65699	 => std_logic_vector(to_unsigned(47,8) ,
65700	 => std_logic_vector(to_unsigned(31,8) ,
65701	 => std_logic_vector(to_unsigned(40,8) ,
65702	 => std_logic_vector(to_unsigned(43,8) ,
65703	 => std_logic_vector(to_unsigned(35,8) ,
65704	 => std_logic_vector(to_unsigned(30,8) ,
65705	 => std_logic_vector(to_unsigned(30,8) ,
65706	 => std_logic_vector(to_unsigned(24,8) ,
65707	 => std_logic_vector(to_unsigned(15,8) ,
65708	 => std_logic_vector(to_unsigned(20,8) ,
65709	 => std_logic_vector(to_unsigned(39,8) ,
65710	 => std_logic_vector(to_unsigned(37,8) ,
65711	 => std_logic_vector(to_unsigned(37,8) ,
65712	 => std_logic_vector(to_unsigned(57,8) ,
65713	 => std_logic_vector(to_unsigned(131,8) ,
65714	 => std_logic_vector(to_unsigned(125,8) ,
65715	 => std_logic_vector(to_unsigned(57,8) ,
65716	 => std_logic_vector(to_unsigned(31,8) ,
65717	 => std_logic_vector(to_unsigned(37,8) ,
65718	 => std_logic_vector(to_unsigned(48,8) ,
65719	 => std_logic_vector(to_unsigned(32,8) ,
65720	 => std_logic_vector(to_unsigned(49,8) ,
65721	 => std_logic_vector(to_unsigned(55,8) ,
65722	 => std_logic_vector(to_unsigned(48,8) ,
65723	 => std_logic_vector(to_unsigned(46,8) ,
65724	 => std_logic_vector(to_unsigned(47,8) ,
65725	 => std_logic_vector(to_unsigned(38,8) ,
65726	 => std_logic_vector(to_unsigned(37,8) ,
65727	 => std_logic_vector(to_unsigned(41,8) ,
65728	 => std_logic_vector(to_unsigned(25,8) ,
65729	 => std_logic_vector(to_unsigned(49,8) ,
65730	 => std_logic_vector(to_unsigned(51,8) ,
65731	 => std_logic_vector(to_unsigned(68,8) ,
65732	 => std_logic_vector(to_unsigned(104,8) ,
65733	 => std_logic_vector(to_unsigned(59,8) ,
65734	 => std_logic_vector(to_unsigned(30,8) ,
65735	 => std_logic_vector(to_unsigned(34,8) ,
65736	 => std_logic_vector(to_unsigned(35,8) ,
65737	 => std_logic_vector(to_unsigned(41,8) ,
65738	 => std_logic_vector(to_unsigned(73,8) ,
65739	 => std_logic_vector(to_unsigned(50,8) ,
65740	 => std_logic_vector(to_unsigned(22,8) ,
65741	 => std_logic_vector(to_unsigned(25,8) ,
65742	 => std_logic_vector(to_unsigned(22,8) ,
65743	 => std_logic_vector(to_unsigned(23,8) ,
65744	 => std_logic_vector(to_unsigned(13,8) ,
65745	 => std_logic_vector(to_unsigned(14,8) ,
65746	 => std_logic_vector(to_unsigned(15,8) ,
65747	 => std_logic_vector(to_unsigned(9,8) ,
65748	 => std_logic_vector(to_unsigned(25,8) ,
65749	 => std_logic_vector(to_unsigned(92,8) ,
65750	 => std_logic_vector(to_unsigned(68,8) ,
65751	 => std_logic_vector(to_unsigned(59,8) ,
65752	 => std_logic_vector(to_unsigned(78,8) ,
65753	 => std_logic_vector(to_unsigned(77,8) ,
65754	 => std_logic_vector(to_unsigned(70,8) ,
65755	 => std_logic_vector(to_unsigned(76,8) ,
65756	 => std_logic_vector(to_unsigned(44,8) ,
65757	 => std_logic_vector(to_unsigned(13,8) ,
65758	 => std_logic_vector(to_unsigned(8,8) ,
65759	 => std_logic_vector(to_unsigned(4,8) ,
65760	 => std_logic_vector(to_unsigned(13,8) ,
65761	 => std_logic_vector(to_unsigned(23,8) ,
65762	 => std_logic_vector(to_unsigned(13,8) ,
65763	 => std_logic_vector(to_unsigned(19,8) ,
65764	 => std_logic_vector(to_unsigned(34,8) ,
65765	 => std_logic_vector(to_unsigned(30,8) ,
65766	 => std_logic_vector(to_unsigned(18,8) ,
65767	 => std_logic_vector(to_unsigned(17,8) ,
65768	 => std_logic_vector(to_unsigned(30,8) ,
65769	 => std_logic_vector(to_unsigned(59,8) ,
65770	 => std_logic_vector(to_unsigned(33,8) ,
65771	 => std_logic_vector(to_unsigned(27,8) ,
65772	 => std_logic_vector(to_unsigned(54,8) ,
65773	 => std_logic_vector(to_unsigned(27,8) ,
65774	 => std_logic_vector(to_unsigned(21,8) ,
65775	 => std_logic_vector(to_unsigned(62,8) ,
65776	 => std_logic_vector(to_unsigned(44,8) ,
65777	 => std_logic_vector(to_unsigned(25,8) ,
65778	 => std_logic_vector(to_unsigned(32,8) ,
65779	 => std_logic_vector(to_unsigned(26,8) ,
65780	 => std_logic_vector(to_unsigned(23,8) ,
65781	 => std_logic_vector(to_unsigned(9,8) ,
65782	 => std_logic_vector(to_unsigned(7,8) ,
65783	 => std_logic_vector(to_unsigned(10,8) ,
65784	 => std_logic_vector(to_unsigned(10,8) ,
65785	 => std_logic_vector(to_unsigned(14,8) ,
65786	 => std_logic_vector(to_unsigned(37,8) ,
65787	 => std_logic_vector(to_unsigned(62,8) ,
65788	 => std_logic_vector(to_unsigned(76,8) ,
65789	 => std_logic_vector(to_unsigned(72,8) ,
65790	 => std_logic_vector(to_unsigned(51,8) ,
65791	 => std_logic_vector(to_unsigned(55,8) ,
65792	 => std_logic_vector(to_unsigned(50,8) ,
65793	 => std_logic_vector(to_unsigned(34,8) ,
65794	 => std_logic_vector(to_unsigned(37,8) ,
65795	 => std_logic_vector(to_unsigned(53,8) ,
65796	 => std_logic_vector(to_unsigned(52,8) ,
65797	 => std_logic_vector(to_unsigned(29,8) ,
65798	 => std_logic_vector(to_unsigned(15,8) ,
65799	 => std_logic_vector(to_unsigned(22,8) ,
65800	 => std_logic_vector(to_unsigned(38,8) ,
65801	 => std_logic_vector(to_unsigned(40,8) ,
65802	 => std_logic_vector(to_unsigned(32,8) ,
65803	 => std_logic_vector(to_unsigned(16,8) ,
65804	 => std_logic_vector(to_unsigned(16,8) ,
65805	 => std_logic_vector(to_unsigned(22,8) ,
65806	 => std_logic_vector(to_unsigned(16,8) ,
65807	 => std_logic_vector(to_unsigned(13,8) ,
65808	 => std_logic_vector(to_unsigned(37,8) ,
65809	 => std_logic_vector(to_unsigned(41,8) ,
65810	 => std_logic_vector(to_unsigned(35,8) ,
65811	 => std_logic_vector(to_unsigned(24,8) ,
65812	 => std_logic_vector(to_unsigned(32,8) ,
65813	 => std_logic_vector(to_unsigned(43,8) ,
65814	 => std_logic_vector(to_unsigned(20,8) ,
65815	 => std_logic_vector(to_unsigned(12,8) ,
65816	 => std_logic_vector(to_unsigned(29,8) ,
65817	 => std_logic_vector(to_unsigned(37,8) ,
65818	 => std_logic_vector(to_unsigned(45,8) ,
65819	 => std_logic_vector(to_unsigned(19,8) ,
65820	 => std_logic_vector(to_unsigned(5,8) ,
65821	 => std_logic_vector(to_unsigned(6,8) ,
65822	 => std_logic_vector(to_unsigned(5,8) ,
65823	 => std_logic_vector(to_unsigned(36,8) ,
65824	 => std_logic_vector(to_unsigned(52,8) ,
65825	 => std_logic_vector(to_unsigned(44,8) ,
65826	 => std_logic_vector(to_unsigned(36,8) ,
65827	 => std_logic_vector(to_unsigned(39,8) ,
65828	 => std_logic_vector(to_unsigned(31,8) ,
65829	 => std_logic_vector(to_unsigned(12,8) ,
65830	 => std_logic_vector(to_unsigned(37,8) ,
65831	 => std_logic_vector(to_unsigned(73,8) ,
65832	 => std_logic_vector(to_unsigned(25,8) ,
65833	 => std_logic_vector(to_unsigned(12,8) ,
65834	 => std_logic_vector(to_unsigned(17,8) ,
65835	 => std_logic_vector(to_unsigned(52,8) ,
65836	 => std_logic_vector(to_unsigned(82,8) ,
65837	 => std_logic_vector(to_unsigned(73,8) ,
65838	 => std_logic_vector(to_unsigned(33,8) ,
65839	 => std_logic_vector(to_unsigned(36,8) ,
65840	 => std_logic_vector(to_unsigned(101,8) ,
65841	 => std_logic_vector(to_unsigned(69,8) ,
65842	 => std_logic_vector(to_unsigned(107,8) ,
65843	 => std_logic_vector(to_unsigned(151,8) ,
65844	 => std_logic_vector(to_unsigned(116,8) ,
65845	 => std_logic_vector(to_unsigned(48,8) ,
65846	 => std_logic_vector(to_unsigned(24,8) ,
65847	 => std_logic_vector(to_unsigned(16,8) ,
65848	 => std_logic_vector(to_unsigned(49,8) ,
65849	 => std_logic_vector(to_unsigned(85,8) ,
65850	 => std_logic_vector(to_unsigned(55,8) ,
65851	 => std_logic_vector(to_unsigned(22,8) ,
65852	 => std_logic_vector(to_unsigned(16,8) ,
65853	 => std_logic_vector(to_unsigned(13,8) ,
65854	 => std_logic_vector(to_unsigned(13,8) ,
65855	 => std_logic_vector(to_unsigned(10,8) ,
65856	 => std_logic_vector(to_unsigned(12,8) ,
65857	 => std_logic_vector(to_unsigned(10,8) ,
65858	 => std_logic_vector(to_unsigned(16,8) ,
65859	 => std_logic_vector(to_unsigned(14,8) ,
65860	 => std_logic_vector(to_unsigned(10,8) ,
65861	 => std_logic_vector(to_unsigned(18,8) ,
65862	 => std_logic_vector(to_unsigned(26,8) ,
65863	 => std_logic_vector(to_unsigned(29,8) ,
65864	 => std_logic_vector(to_unsigned(19,8) ,
65865	 => std_logic_vector(to_unsigned(25,8) ,
65866	 => std_logic_vector(to_unsigned(41,8) ,
65867	 => std_logic_vector(to_unsigned(38,8) ,
65868	 => std_logic_vector(to_unsigned(32,8) ,
65869	 => std_logic_vector(to_unsigned(17,8) ,
65870	 => std_logic_vector(to_unsigned(41,8) ,
65871	 => std_logic_vector(to_unsigned(22,8) ,
65872	 => std_logic_vector(to_unsigned(0,8) ,
65873	 => std_logic_vector(to_unsigned(1,8) ,
65874	 => std_logic_vector(to_unsigned(15,8) ,
65875	 => std_logic_vector(to_unsigned(30,8) ,
65876	 => std_logic_vector(to_unsigned(27,8) ,
65877	 => std_logic_vector(to_unsigned(29,8) ,
65878	 => std_logic_vector(to_unsigned(26,8) ,
65879	 => std_logic_vector(to_unsigned(17,8) ,
65880	 => std_logic_vector(to_unsigned(12,8) ,
65881	 => std_logic_vector(to_unsigned(17,8) ,
65882	 => std_logic_vector(to_unsigned(17,8) ,
65883	 => std_logic_vector(to_unsigned(12,8) ,
65884	 => std_logic_vector(to_unsigned(13,8) ,
65885	 => std_logic_vector(to_unsigned(1,8) ,
65886	 => std_logic_vector(to_unsigned(0,8) ,
65887	 => std_logic_vector(to_unsigned(4,8) ,
65888	 => std_logic_vector(to_unsigned(22,8) ,
65889	 => std_logic_vector(to_unsigned(16,8) ,
65890	 => std_logic_vector(to_unsigned(19,8) ,
65891	 => std_logic_vector(to_unsigned(21,8) ,
65892	 => std_logic_vector(to_unsigned(25,8) ,
65893	 => std_logic_vector(to_unsigned(26,8) ,
65894	 => std_logic_vector(to_unsigned(13,8) ,
65895	 => std_logic_vector(to_unsigned(8,8) ,
65896	 => std_logic_vector(to_unsigned(1,8) ,
65897	 => std_logic_vector(to_unsigned(0,8) ,
65898	 => std_logic_vector(to_unsigned(6,8) ,
65899	 => std_logic_vector(to_unsigned(32,8) ,
65900	 => std_logic_vector(to_unsigned(26,8) ,
65901	 => std_logic_vector(to_unsigned(23,8) ,
65902	 => std_logic_vector(to_unsigned(20,8) ,
65903	 => std_logic_vector(to_unsigned(29,8) ,
65904	 => std_logic_vector(to_unsigned(26,8) ,
65905	 => std_logic_vector(to_unsigned(27,8) ,
65906	 => std_logic_vector(to_unsigned(30,8) ,
65907	 => std_logic_vector(to_unsigned(27,8) ,
65908	 => std_logic_vector(to_unsigned(23,8) ,
65909	 => std_logic_vector(to_unsigned(12,8) ,
65910	 => std_logic_vector(to_unsigned(20,8) ,
65911	 => std_logic_vector(to_unsigned(33,8) ,
65912	 => std_logic_vector(to_unsigned(35,8) ,
65913	 => std_logic_vector(to_unsigned(34,8) ,
65914	 => std_logic_vector(to_unsigned(26,8) ,
65915	 => std_logic_vector(to_unsigned(24,8) ,
65916	 => std_logic_vector(to_unsigned(22,8) ,
65917	 => std_logic_vector(to_unsigned(43,8) ,
65918	 => std_logic_vector(to_unsigned(61,8) ,
65919	 => std_logic_vector(to_unsigned(48,8) ,
65920	 => std_logic_vector(to_unsigned(29,8) ,
65921	 => std_logic_vector(to_unsigned(124,8) ,
65922	 => std_logic_vector(to_unsigned(124,8) ,
65923	 => std_logic_vector(to_unsigned(122,8) ,
65924	 => std_logic_vector(to_unsigned(99,8) ,
65925	 => std_logic_vector(to_unsigned(107,8) ,
65926	 => std_logic_vector(to_unsigned(111,8) ,
65927	 => std_logic_vector(to_unsigned(101,8) ,
65928	 => std_logic_vector(to_unsigned(97,8) ,
65929	 => std_logic_vector(to_unsigned(95,8) ,
65930	 => std_logic_vector(to_unsigned(101,8) ,
65931	 => std_logic_vector(to_unsigned(82,8) ,
65932	 => std_logic_vector(to_unsigned(45,8) ,
65933	 => std_logic_vector(to_unsigned(37,8) ,
65934	 => std_logic_vector(to_unsigned(24,8) ,
65935	 => std_logic_vector(to_unsigned(38,8) ,
65936	 => std_logic_vector(to_unsigned(72,8) ,
65937	 => std_logic_vector(to_unsigned(73,8) ,
65938	 => std_logic_vector(to_unsigned(69,8) ,
65939	 => std_logic_vector(to_unsigned(55,8) ,
65940	 => std_logic_vector(to_unsigned(84,8) ,
65941	 => std_logic_vector(to_unsigned(128,8) ,
65942	 => std_logic_vector(to_unsigned(128,8) ,
65943	 => std_logic_vector(to_unsigned(90,8) ,
65944	 => std_logic_vector(to_unsigned(46,8) ,
65945	 => std_logic_vector(to_unsigned(48,8) ,
65946	 => std_logic_vector(to_unsigned(37,8) ,
65947	 => std_logic_vector(to_unsigned(32,8) ,
65948	 => std_logic_vector(to_unsigned(35,8) ,
65949	 => std_logic_vector(to_unsigned(35,8) ,
65950	 => std_logic_vector(to_unsigned(39,8) ,
65951	 => std_logic_vector(to_unsigned(33,8) ,
65952	 => std_logic_vector(to_unsigned(30,8) ,
65953	 => std_logic_vector(to_unsigned(32,8) ,
65954	 => std_logic_vector(to_unsigned(34,8) ,
65955	 => std_logic_vector(to_unsigned(32,8) ,
65956	 => std_logic_vector(to_unsigned(27,8) ,
65957	 => std_logic_vector(to_unsigned(28,8) ,
65958	 => std_logic_vector(to_unsigned(22,8) ,
65959	 => std_logic_vector(to_unsigned(18,8) ,
65960	 => std_logic_vector(to_unsigned(19,8) ,
65961	 => std_logic_vector(to_unsigned(18,8) ,
65962	 => std_logic_vector(to_unsigned(21,8) ,
65963	 => std_logic_vector(to_unsigned(24,8) ,
65964	 => std_logic_vector(to_unsigned(30,8) ,
65965	 => std_logic_vector(to_unsigned(35,8) ,
65966	 => std_logic_vector(to_unsigned(37,8) ,
65967	 => std_logic_vector(to_unsigned(43,8) ,
65968	 => std_logic_vector(to_unsigned(44,8) ,
65969	 => std_logic_vector(to_unsigned(37,8) ,
65970	 => std_logic_vector(to_unsigned(35,8) ,
65971	 => std_logic_vector(to_unsigned(40,8) ,
65972	 => std_logic_vector(to_unsigned(45,8) ,
65973	 => std_logic_vector(to_unsigned(31,8) ,
65974	 => std_logic_vector(to_unsigned(37,8) ,
65975	 => std_logic_vector(to_unsigned(37,8) ,
65976	 => std_logic_vector(to_unsigned(54,8) ,
65977	 => std_logic_vector(to_unsigned(88,8) ,
65978	 => std_logic_vector(to_unsigned(82,8) ,
65979	 => std_logic_vector(to_unsigned(82,8) ,
65980	 => std_logic_vector(to_unsigned(88,8) ,
65981	 => std_logic_vector(to_unsigned(87,8) ,
65982	 => std_logic_vector(to_unsigned(74,8) ,
65983	 => std_logic_vector(to_unsigned(78,8) ,
65984	 => std_logic_vector(to_unsigned(81,8) ,
65985	 => std_logic_vector(to_unsigned(85,8) ,
65986	 => std_logic_vector(to_unsigned(86,8) ,
65987	 => std_logic_vector(to_unsigned(92,8) ,
65988	 => std_logic_vector(to_unsigned(93,8) ,
65989	 => std_logic_vector(to_unsigned(78,8) ,
65990	 => std_logic_vector(to_unsigned(86,8) ,
65991	 => std_logic_vector(to_unsigned(100,8) ,
65992	 => std_logic_vector(to_unsigned(112,8) ,
65993	 => std_logic_vector(to_unsigned(111,8) ,
65994	 => std_logic_vector(to_unsigned(108,8) ,
65995	 => std_logic_vector(to_unsigned(99,8) ,
65996	 => std_logic_vector(to_unsigned(88,8) ,
65997	 => std_logic_vector(to_unsigned(87,8) ,
65998	 => std_logic_vector(to_unsigned(104,8) ,
65999	 => std_logic_vector(to_unsigned(71,8) ,
66000	 => std_logic_vector(to_unsigned(33,8) ,
66001	 => std_logic_vector(to_unsigned(56,8) ,
66002	 => std_logic_vector(to_unsigned(81,8) ,
66003	 => std_logic_vector(to_unsigned(71,8) ,
66004	 => std_logic_vector(to_unsigned(74,8) ,
66005	 => std_logic_vector(to_unsigned(77,8) ,
66006	 => std_logic_vector(to_unsigned(71,8) ,
66007	 => std_logic_vector(to_unsigned(57,8) ,
66008	 => std_logic_vector(to_unsigned(40,8) ,
66009	 => std_logic_vector(to_unsigned(35,8) ,
66010	 => std_logic_vector(to_unsigned(31,8) ,
66011	 => std_logic_vector(to_unsigned(40,8) ,
66012	 => std_logic_vector(to_unsigned(52,8) ,
66013	 => std_logic_vector(to_unsigned(57,8) ,
66014	 => std_logic_vector(to_unsigned(54,8) ,
66015	 => std_logic_vector(to_unsigned(63,8) ,
66016	 => std_logic_vector(to_unsigned(76,8) ,
66017	 => std_logic_vector(to_unsigned(66,8) ,
66018	 => std_logic_vector(to_unsigned(76,8) ,
66019	 => std_logic_vector(to_unsigned(58,8) ,
66020	 => std_logic_vector(to_unsigned(57,8) ,
66021	 => std_logic_vector(to_unsigned(50,8) ,
66022	 => std_logic_vector(to_unsigned(41,8) ,
66023	 => std_logic_vector(to_unsigned(29,8) ,
66024	 => std_logic_vector(to_unsigned(24,8) ,
66025	 => std_logic_vector(to_unsigned(27,8) ,
66026	 => std_logic_vector(to_unsigned(25,8) ,
66027	 => std_logic_vector(to_unsigned(18,8) ,
66028	 => std_logic_vector(to_unsigned(21,8) ,
66029	 => std_logic_vector(to_unsigned(54,8) ,
66030	 => std_logic_vector(to_unsigned(73,8) ,
66031	 => std_logic_vector(to_unsigned(60,8) ,
66032	 => std_logic_vector(to_unsigned(51,8) ,
66033	 => std_logic_vector(to_unsigned(48,8) ,
66034	 => std_logic_vector(to_unsigned(41,8) ,
66035	 => std_logic_vector(to_unsigned(40,8) ,
66036	 => std_logic_vector(to_unsigned(40,8) ,
66037	 => std_logic_vector(to_unsigned(42,8) ,
66038	 => std_logic_vector(to_unsigned(40,8) ,
66039	 => std_logic_vector(to_unsigned(19,8) ,
66040	 => std_logic_vector(to_unsigned(41,8) ,
66041	 => std_logic_vector(to_unsigned(57,8) ,
66042	 => std_logic_vector(to_unsigned(33,8) ,
66043	 => std_logic_vector(to_unsigned(31,8) ,
66044	 => std_logic_vector(to_unsigned(46,8) ,
66045	 => std_logic_vector(to_unsigned(37,8) ,
66046	 => std_logic_vector(to_unsigned(41,8) ,
66047	 => std_logic_vector(to_unsigned(43,8) ,
66048	 => std_logic_vector(to_unsigned(18,8) ,
66049	 => std_logic_vector(to_unsigned(24,8) ,
66050	 => std_logic_vector(to_unsigned(26,8) ,
66051	 => std_logic_vector(to_unsigned(33,8) ,
66052	 => std_logic_vector(to_unsigned(46,8) ,
66053	 => std_logic_vector(to_unsigned(37,8) ,
66054	 => std_logic_vector(to_unsigned(38,8) ,
66055	 => std_logic_vector(to_unsigned(37,8) ,
66056	 => std_logic_vector(to_unsigned(37,8) ,
66057	 => std_logic_vector(to_unsigned(40,8) ,
66058	 => std_logic_vector(to_unsigned(58,8) ,
66059	 => std_logic_vector(to_unsigned(37,8) ,
66060	 => std_logic_vector(to_unsigned(36,8) ,
66061	 => std_logic_vector(to_unsigned(25,8) ,
66062	 => std_logic_vector(to_unsigned(15,8) ,
66063	 => std_logic_vector(to_unsigned(31,8) ,
66064	 => std_logic_vector(to_unsigned(26,8) ,
66065	 => std_logic_vector(to_unsigned(18,8) ,
66066	 => std_logic_vector(to_unsigned(23,8) ,
66067	 => std_logic_vector(to_unsigned(18,8) ,
66068	 => std_logic_vector(to_unsigned(29,8) ,
66069	 => std_logic_vector(to_unsigned(101,8) ,
66070	 => std_logic_vector(to_unsigned(61,8) ,
66071	 => std_logic_vector(to_unsigned(22,8) ,
66072	 => std_logic_vector(to_unsigned(85,8) ,
66073	 => std_logic_vector(to_unsigned(44,8) ,
66074	 => std_logic_vector(to_unsigned(37,8) ,
66075	 => std_logic_vector(to_unsigned(85,8) ,
66076	 => std_logic_vector(to_unsigned(45,8) ,
66077	 => std_logic_vector(to_unsigned(10,8) ,
66078	 => std_logic_vector(to_unsigned(8,8) ,
66079	 => std_logic_vector(to_unsigned(5,8) ,
66080	 => std_logic_vector(to_unsigned(15,8) ,
66081	 => std_logic_vector(to_unsigned(32,8) ,
66082	 => std_logic_vector(to_unsigned(22,8) ,
66083	 => std_logic_vector(to_unsigned(17,8) ,
66084	 => std_logic_vector(to_unsigned(32,8) ,
66085	 => std_logic_vector(to_unsigned(27,8) ,
66086	 => std_logic_vector(to_unsigned(13,8) ,
66087	 => std_logic_vector(to_unsigned(10,8) ,
66088	 => std_logic_vector(to_unsigned(16,8) ,
66089	 => std_logic_vector(to_unsigned(52,8) ,
66090	 => std_logic_vector(to_unsigned(34,8) ,
66091	 => std_logic_vector(to_unsigned(23,8) ,
66092	 => std_logic_vector(to_unsigned(25,8) ,
66093	 => std_logic_vector(to_unsigned(22,8) ,
66094	 => std_logic_vector(to_unsigned(58,8) ,
66095	 => std_logic_vector(to_unsigned(55,8) ,
66096	 => std_logic_vector(to_unsigned(54,8) ,
66097	 => std_logic_vector(to_unsigned(41,8) ,
66098	 => std_logic_vector(to_unsigned(22,8) ,
66099	 => std_logic_vector(to_unsigned(29,8) ,
66100	 => std_logic_vector(to_unsigned(35,8) ,
66101	 => std_logic_vector(to_unsigned(10,8) ,
66102	 => std_logic_vector(to_unsigned(7,8) ,
66103	 => std_logic_vector(to_unsigned(9,8) ,
66104	 => std_logic_vector(to_unsigned(10,8) ,
66105	 => std_logic_vector(to_unsigned(18,8) ,
66106	 => std_logic_vector(to_unsigned(39,8) ,
66107	 => std_logic_vector(to_unsigned(31,8) ,
66108	 => std_logic_vector(to_unsigned(20,8) ,
66109	 => std_logic_vector(to_unsigned(26,8) ,
66110	 => std_logic_vector(to_unsigned(46,8) ,
66111	 => std_logic_vector(to_unsigned(56,8) ,
66112	 => std_logic_vector(to_unsigned(60,8) ,
66113	 => std_logic_vector(to_unsigned(72,8) ,
66114	 => std_logic_vector(to_unsigned(65,8) ,
66115	 => std_logic_vector(to_unsigned(47,8) ,
66116	 => std_logic_vector(to_unsigned(47,8) ,
66117	 => std_logic_vector(to_unsigned(50,8) ,
66118	 => std_logic_vector(to_unsigned(45,8) ,
66119	 => std_logic_vector(to_unsigned(29,8) ,
66120	 => std_logic_vector(to_unsigned(40,8) ,
66121	 => std_logic_vector(to_unsigned(45,8) ,
66122	 => std_logic_vector(to_unsigned(26,8) ,
66123	 => std_logic_vector(to_unsigned(12,8) ,
66124	 => std_logic_vector(to_unsigned(27,8) ,
66125	 => std_logic_vector(to_unsigned(38,8) ,
66126	 => std_logic_vector(to_unsigned(18,8) ,
66127	 => std_logic_vector(to_unsigned(9,8) ,
66128	 => std_logic_vector(to_unsigned(27,8) ,
66129	 => std_logic_vector(to_unsigned(45,8) ,
66130	 => std_logic_vector(to_unsigned(46,8) ,
66131	 => std_logic_vector(to_unsigned(41,8) ,
66132	 => std_logic_vector(to_unsigned(36,8) ,
66133	 => std_logic_vector(to_unsigned(35,8) ,
66134	 => std_logic_vector(to_unsigned(34,8) ,
66135	 => std_logic_vector(to_unsigned(28,8) ,
66136	 => std_logic_vector(to_unsigned(19,8) ,
66137	 => std_logic_vector(to_unsigned(22,8) ,
66138	 => std_logic_vector(to_unsigned(32,8) ,
66139	 => std_logic_vector(to_unsigned(23,8) ,
66140	 => std_logic_vector(to_unsigned(11,8) ,
66141	 => std_logic_vector(to_unsigned(9,8) ,
66142	 => std_logic_vector(to_unsigned(5,8) ,
66143	 => std_logic_vector(to_unsigned(30,8) ,
66144	 => std_logic_vector(to_unsigned(52,8) ,
66145	 => std_logic_vector(to_unsigned(41,8) ,
66146	 => std_logic_vector(to_unsigned(35,8) ,
66147	 => std_logic_vector(to_unsigned(39,8) ,
66148	 => std_logic_vector(to_unsigned(26,8) ,
66149	 => std_logic_vector(to_unsigned(8,8) ,
66150	 => std_logic_vector(to_unsigned(22,8) ,
66151	 => std_logic_vector(to_unsigned(35,8) ,
66152	 => std_logic_vector(to_unsigned(20,8) ,
66153	 => std_logic_vector(to_unsigned(11,8) ,
66154	 => std_logic_vector(to_unsigned(18,8) ,
66155	 => std_logic_vector(to_unsigned(55,8) ,
66156	 => std_logic_vector(to_unsigned(84,8) ,
66157	 => std_logic_vector(to_unsigned(51,8) ,
66158	 => std_logic_vector(to_unsigned(23,8) ,
66159	 => std_logic_vector(to_unsigned(23,8) ,
66160	 => std_logic_vector(to_unsigned(38,8) ,
66161	 => std_logic_vector(to_unsigned(35,8) ,
66162	 => std_logic_vector(to_unsigned(61,8) ,
66163	 => std_logic_vector(to_unsigned(121,8) ,
66164	 => std_logic_vector(to_unsigned(127,8) ,
66165	 => std_logic_vector(to_unsigned(39,8) ,
66166	 => std_logic_vector(to_unsigned(29,8) ,
66167	 => std_logic_vector(to_unsigned(78,8) ,
66168	 => std_logic_vector(to_unsigned(95,8) ,
66169	 => std_logic_vector(to_unsigned(93,8) ,
66170	 => std_logic_vector(to_unsigned(55,8) ,
66171	 => std_logic_vector(to_unsigned(19,8) ,
66172	 => std_logic_vector(to_unsigned(21,8) ,
66173	 => std_logic_vector(to_unsigned(22,8) ,
66174	 => std_logic_vector(to_unsigned(15,8) ,
66175	 => std_logic_vector(to_unsigned(17,8) ,
66176	 => std_logic_vector(to_unsigned(23,8) ,
66177	 => std_logic_vector(to_unsigned(14,8) ,
66178	 => std_logic_vector(to_unsigned(25,8) ,
66179	 => std_logic_vector(to_unsigned(20,8) ,
66180	 => std_logic_vector(to_unsigned(17,8) ,
66181	 => std_logic_vector(to_unsigned(12,8) ,
66182	 => std_logic_vector(to_unsigned(14,8) ,
66183	 => std_logic_vector(to_unsigned(12,8) ,
66184	 => std_logic_vector(to_unsigned(14,8) ,
66185	 => std_logic_vector(to_unsigned(37,8) ,
66186	 => std_logic_vector(to_unsigned(37,8) ,
66187	 => std_logic_vector(to_unsigned(37,8) ,
66188	 => std_logic_vector(to_unsigned(30,8) ,
66189	 => std_logic_vector(to_unsigned(23,8) ,
66190	 => std_logic_vector(to_unsigned(40,8) ,
66191	 => std_logic_vector(to_unsigned(21,8) ,
66192	 => std_logic_vector(to_unsigned(1,8) ,
66193	 => std_logic_vector(to_unsigned(0,8) ,
66194	 => std_logic_vector(to_unsigned(9,8) ,
66195	 => std_logic_vector(to_unsigned(36,8) ,
66196	 => std_logic_vector(to_unsigned(28,8) ,
66197	 => std_logic_vector(to_unsigned(29,8) ,
66198	 => std_logic_vector(to_unsigned(17,8) ,
66199	 => std_logic_vector(to_unsigned(10,8) ,
66200	 => std_logic_vector(to_unsigned(14,8) ,
66201	 => std_logic_vector(to_unsigned(18,8) ,
66202	 => std_logic_vector(to_unsigned(8,8) ,
66203	 => std_logic_vector(to_unsigned(6,8) ,
66204	 => std_logic_vector(to_unsigned(13,8) ,
66205	 => std_logic_vector(to_unsigned(2,8) ,
66206	 => std_logic_vector(to_unsigned(0,8) ,
66207	 => std_logic_vector(to_unsigned(5,8) ,
66208	 => std_logic_vector(to_unsigned(15,8) ,
66209	 => std_logic_vector(to_unsigned(9,8) ,
66210	 => std_logic_vector(to_unsigned(21,8) ,
66211	 => std_logic_vector(to_unsigned(28,8) ,
66212	 => std_logic_vector(to_unsigned(29,8) ,
66213	 => std_logic_vector(to_unsigned(26,8) ,
66214	 => std_logic_vector(to_unsigned(8,8) ,
66215	 => std_logic_vector(to_unsigned(28,8) ,
66216	 => std_logic_vector(to_unsigned(10,8) ,
66217	 => std_logic_vector(to_unsigned(0,8) ,
66218	 => std_logic_vector(to_unsigned(1,8) ,
66219	 => std_logic_vector(to_unsigned(24,8) ,
66220	 => std_logic_vector(to_unsigned(37,8) ,
66221	 => std_logic_vector(to_unsigned(29,8) ,
66222	 => std_logic_vector(to_unsigned(31,8) ,
66223	 => std_logic_vector(to_unsigned(35,8) ,
66224	 => std_logic_vector(to_unsigned(37,8) ,
66225	 => std_logic_vector(to_unsigned(32,8) ,
66226	 => std_logic_vector(to_unsigned(26,8) ,
66227	 => std_logic_vector(to_unsigned(17,8) ,
66228	 => std_logic_vector(to_unsigned(19,8) ,
66229	 => std_logic_vector(to_unsigned(21,8) ,
66230	 => std_logic_vector(to_unsigned(31,8) ,
66231	 => std_logic_vector(to_unsigned(33,8) ,
66232	 => std_logic_vector(to_unsigned(33,8) ,
66233	 => std_logic_vector(to_unsigned(37,8) ,
66234	 => std_logic_vector(to_unsigned(35,8) ,
66235	 => std_logic_vector(to_unsigned(24,8) ,
66236	 => std_logic_vector(to_unsigned(15,8) ,
66237	 => std_logic_vector(to_unsigned(51,8) ,
66238	 => std_logic_vector(to_unsigned(100,8) ,
66239	 => std_logic_vector(to_unsigned(91,8) ,
66240	 => std_logic_vector(to_unsigned(84,8) ,
66241	 => std_logic_vector(to_unsigned(101,8) ,
66242	 => std_logic_vector(to_unsigned(124,8) ,
66243	 => std_logic_vector(to_unsigned(125,8) ,
66244	 => std_logic_vector(to_unsigned(121,8) ,
66245	 => std_logic_vector(to_unsigned(111,8) ,
66246	 => std_logic_vector(to_unsigned(111,8) ,
66247	 => std_logic_vector(to_unsigned(107,8) ,
66248	 => std_logic_vector(to_unsigned(103,8) ,
66249	 => std_logic_vector(to_unsigned(99,8) ,
66250	 => std_logic_vector(to_unsigned(92,8) ,
66251	 => std_logic_vector(to_unsigned(62,8) ,
66252	 => std_logic_vector(to_unsigned(39,8) ,
66253	 => std_logic_vector(to_unsigned(35,8) ,
66254	 => std_logic_vector(to_unsigned(32,8) ,
66255	 => std_logic_vector(to_unsigned(51,8) ,
66256	 => std_logic_vector(to_unsigned(73,8) ,
66257	 => std_logic_vector(to_unsigned(80,8) ,
66258	 => std_logic_vector(to_unsigned(77,8) ,
66259	 => std_logic_vector(to_unsigned(66,8) ,
66260	 => std_logic_vector(to_unsigned(81,8) ,
66261	 => std_logic_vector(to_unsigned(116,8) ,
66262	 => std_logic_vector(to_unsigned(119,8) ,
66263	 => std_logic_vector(to_unsigned(101,8) ,
66264	 => std_logic_vector(to_unsigned(55,8) ,
66265	 => std_logic_vector(to_unsigned(44,8) ,
66266	 => std_logic_vector(to_unsigned(45,8) ,
66267	 => std_logic_vector(to_unsigned(41,8) ,
66268	 => std_logic_vector(to_unsigned(35,8) ,
66269	 => std_logic_vector(to_unsigned(34,8) ,
66270	 => std_logic_vector(to_unsigned(36,8) ,
66271	 => std_logic_vector(to_unsigned(27,8) ,
66272	 => std_logic_vector(to_unsigned(27,8) ,
66273	 => std_logic_vector(to_unsigned(30,8) ,
66274	 => std_logic_vector(to_unsigned(30,8) ,
66275	 => std_logic_vector(to_unsigned(27,8) ,
66276	 => std_logic_vector(to_unsigned(26,8) ,
66277	 => std_logic_vector(to_unsigned(25,8) ,
66278	 => std_logic_vector(to_unsigned(26,8) ,
66279	 => std_logic_vector(to_unsigned(32,8) ,
66280	 => std_logic_vector(to_unsigned(17,8) ,
66281	 => std_logic_vector(to_unsigned(17,8) ,
66282	 => std_logic_vector(to_unsigned(17,8) ,
66283	 => std_logic_vector(to_unsigned(22,8) ,
66284	 => std_logic_vector(to_unsigned(32,8) ,
66285	 => std_logic_vector(to_unsigned(36,8) ,
66286	 => std_logic_vector(to_unsigned(32,8) ,
66287	 => std_logic_vector(to_unsigned(44,8) ,
66288	 => std_logic_vector(to_unsigned(55,8) ,
66289	 => std_logic_vector(to_unsigned(36,8) ,
66290	 => std_logic_vector(to_unsigned(30,8) ,
66291	 => std_logic_vector(to_unsigned(35,8) ,
66292	 => std_logic_vector(to_unsigned(29,8) ,
66293	 => std_logic_vector(to_unsigned(27,8) ,
66294	 => std_logic_vector(to_unsigned(37,8) ,
66295	 => std_logic_vector(to_unsigned(50,8) ,
66296	 => std_logic_vector(to_unsigned(77,8) ,
66297	 => std_logic_vector(to_unsigned(80,8) ,
66298	 => std_logic_vector(to_unsigned(71,8) ,
66299	 => std_logic_vector(to_unsigned(62,8) ,
66300	 => std_logic_vector(to_unsigned(80,8) ,
66301	 => std_logic_vector(to_unsigned(82,8) ,
66302	 => std_logic_vector(to_unsigned(73,8) ,
66303	 => std_logic_vector(to_unsigned(81,8) ,
66304	 => std_logic_vector(to_unsigned(87,8) ,
66305	 => std_logic_vector(to_unsigned(84,8) ,
66306	 => std_logic_vector(to_unsigned(90,8) ,
66307	 => std_logic_vector(to_unsigned(100,8) ,
66308	 => std_logic_vector(to_unsigned(99,8) ,
66309	 => std_logic_vector(to_unsigned(90,8) ,
66310	 => std_logic_vector(to_unsigned(97,8) ,
66311	 => std_logic_vector(to_unsigned(118,8) ,
66312	 => std_logic_vector(to_unsigned(118,8) ,
66313	 => std_logic_vector(to_unsigned(112,8) ,
66314	 => std_logic_vector(to_unsigned(107,8) ,
66315	 => std_logic_vector(to_unsigned(104,8) ,
66316	 => std_logic_vector(to_unsigned(103,8) ,
66317	 => std_logic_vector(to_unsigned(107,8) ,
66318	 => std_logic_vector(to_unsigned(109,8) ,
66319	 => std_logic_vector(to_unsigned(105,8) ,
66320	 => std_logic_vector(to_unsigned(76,8) ,
66321	 => std_logic_vector(to_unsigned(73,8) ,
66322	 => std_logic_vector(to_unsigned(92,8) ,
66323	 => std_logic_vector(to_unsigned(96,8) ,
66324	 => std_logic_vector(to_unsigned(71,8) ,
66325	 => std_logic_vector(to_unsigned(64,8) ,
66326	 => std_logic_vector(to_unsigned(90,8) ,
66327	 => std_logic_vector(to_unsigned(70,8) ,
66328	 => std_logic_vector(to_unsigned(57,8) ,
66329	 => std_logic_vector(to_unsigned(65,8) ,
66330	 => std_logic_vector(to_unsigned(37,8) ,
66331	 => std_logic_vector(to_unsigned(38,8) ,
66332	 => std_logic_vector(to_unsigned(61,8) ,
66333	 => std_logic_vector(to_unsigned(56,8) ,
66334	 => std_logic_vector(to_unsigned(51,8) ,
66335	 => std_logic_vector(to_unsigned(79,8) ,
66336	 => std_logic_vector(to_unsigned(81,8) ,
66337	 => std_logic_vector(to_unsigned(72,8) ,
66338	 => std_logic_vector(to_unsigned(85,8) ,
66339	 => std_logic_vector(to_unsigned(59,8) ,
66340	 => std_logic_vector(to_unsigned(80,8) ,
66341	 => std_logic_vector(to_unsigned(46,8) ,
66342	 => std_logic_vector(to_unsigned(31,8) ,
66343	 => std_logic_vector(to_unsigned(25,8) ,
66344	 => std_logic_vector(to_unsigned(22,8) ,
66345	 => std_logic_vector(to_unsigned(25,8) ,
66346	 => std_logic_vector(to_unsigned(20,8) ,
66347	 => std_logic_vector(to_unsigned(17,8) ,
66348	 => std_logic_vector(to_unsigned(18,8) ,
66349	 => std_logic_vector(to_unsigned(67,8) ,
66350	 => std_logic_vector(to_unsigned(154,8) ,
66351	 => std_logic_vector(to_unsigned(80,8) ,
66352	 => std_logic_vector(to_unsigned(38,8) ,
66353	 => std_logic_vector(to_unsigned(86,8) ,
66354	 => std_logic_vector(to_unsigned(88,8) ,
66355	 => std_logic_vector(to_unsigned(41,8) ,
66356	 => std_logic_vector(to_unsigned(39,8) ,
66357	 => std_logic_vector(to_unsigned(50,8) ,
66358	 => std_logic_vector(to_unsigned(50,8) ,
66359	 => std_logic_vector(to_unsigned(44,8) ,
66360	 => std_logic_vector(to_unsigned(45,8) ,
66361	 => std_logic_vector(to_unsigned(52,8) ,
66362	 => std_logic_vector(to_unsigned(41,8) ,
66363	 => std_logic_vector(to_unsigned(37,8) ,
66364	 => std_logic_vector(to_unsigned(35,8) ,
66365	 => std_logic_vector(to_unsigned(35,8) ,
66366	 => std_logic_vector(to_unsigned(41,8) ,
66367	 => std_logic_vector(to_unsigned(24,8) ,
66368	 => std_logic_vector(to_unsigned(26,8) ,
66369	 => std_logic_vector(to_unsigned(40,8) ,
66370	 => std_logic_vector(to_unsigned(30,8) ,
66371	 => std_logic_vector(to_unsigned(37,8) ,
66372	 => std_logic_vector(to_unsigned(45,8) ,
66373	 => std_logic_vector(to_unsigned(41,8) ,
66374	 => std_logic_vector(to_unsigned(46,8) ,
66375	 => std_logic_vector(to_unsigned(47,8) ,
66376	 => std_logic_vector(to_unsigned(42,8) ,
66377	 => std_logic_vector(to_unsigned(37,8) ,
66378	 => std_logic_vector(to_unsigned(57,8) ,
66379	 => std_logic_vector(to_unsigned(35,8) ,
66380	 => std_logic_vector(to_unsigned(27,8) ,
66381	 => std_logic_vector(to_unsigned(17,8) ,
66382	 => std_logic_vector(to_unsigned(14,8) ,
66383	 => std_logic_vector(to_unsigned(49,8) ,
66384	 => std_logic_vector(to_unsigned(50,8) ,
66385	 => std_logic_vector(to_unsigned(15,8) ,
66386	 => std_logic_vector(to_unsigned(12,8) ,
66387	 => std_logic_vector(to_unsigned(9,8) ,
66388	 => std_logic_vector(to_unsigned(20,8) ,
66389	 => std_logic_vector(to_unsigned(87,8) ,
66390	 => std_logic_vector(to_unsigned(61,8) ,
66391	 => std_logic_vector(to_unsigned(26,8) ,
66392	 => std_logic_vector(to_unsigned(77,8) ,
66393	 => std_logic_vector(to_unsigned(37,8) ,
66394	 => std_logic_vector(to_unsigned(27,8) ,
66395	 => std_logic_vector(to_unsigned(86,8) ,
66396	 => std_logic_vector(to_unsigned(45,8) ,
66397	 => std_logic_vector(to_unsigned(9,8) ,
66398	 => std_logic_vector(to_unsigned(8,8) ,
66399	 => std_logic_vector(to_unsigned(4,8) ,
66400	 => std_logic_vector(to_unsigned(11,8) ,
66401	 => std_logic_vector(to_unsigned(37,8) ,
66402	 => std_logic_vector(to_unsigned(41,8) ,
66403	 => std_logic_vector(to_unsigned(41,8) ,
66404	 => std_logic_vector(to_unsigned(27,8) ,
66405	 => std_logic_vector(to_unsigned(27,8) ,
66406	 => std_logic_vector(to_unsigned(19,8) ,
66407	 => std_logic_vector(to_unsigned(8,8) ,
66408	 => std_logic_vector(to_unsigned(17,8) ,
66409	 => std_logic_vector(to_unsigned(53,8) ,
66410	 => std_logic_vector(to_unsigned(34,8) ,
66411	 => std_logic_vector(to_unsigned(20,8) ,
66412	 => std_logic_vector(to_unsigned(25,8) ,
66413	 => std_logic_vector(to_unsigned(53,8) ,
66414	 => std_logic_vector(to_unsigned(45,8) ,
66415	 => std_logic_vector(to_unsigned(25,8) ,
66416	 => std_logic_vector(to_unsigned(37,8) ,
66417	 => std_logic_vector(to_unsigned(23,8) ,
66418	 => std_logic_vector(to_unsigned(29,8) ,
66419	 => std_logic_vector(to_unsigned(33,8) ,
66420	 => std_logic_vector(to_unsigned(25,8) ,
66421	 => std_logic_vector(to_unsigned(11,8) ,
66422	 => std_logic_vector(to_unsigned(8,8) ,
66423	 => std_logic_vector(to_unsigned(10,8) ,
66424	 => std_logic_vector(to_unsigned(9,8) ,
66425	 => std_logic_vector(to_unsigned(11,8) ,
66426	 => std_logic_vector(to_unsigned(35,8) ,
66427	 => std_logic_vector(to_unsigned(40,8) ,
66428	 => std_logic_vector(to_unsigned(22,8) ,
66429	 => std_logic_vector(to_unsigned(19,8) ,
66430	 => std_logic_vector(to_unsigned(42,8) ,
66431	 => std_logic_vector(to_unsigned(51,8) ,
66432	 => std_logic_vector(to_unsigned(27,8) ,
66433	 => std_logic_vector(to_unsigned(17,8) ,
66434	 => std_logic_vector(to_unsigned(29,8) ,
66435	 => std_logic_vector(to_unsigned(45,8) ,
66436	 => std_logic_vector(to_unsigned(45,8) ,
66437	 => std_logic_vector(to_unsigned(50,8) ,
66438	 => std_logic_vector(to_unsigned(58,8) ,
66439	 => std_logic_vector(to_unsigned(54,8) ,
66440	 => std_logic_vector(to_unsigned(50,8) ,
66441	 => std_logic_vector(to_unsigned(35,8) ,
66442	 => std_logic_vector(to_unsigned(17,8) ,
66443	 => std_logic_vector(to_unsigned(19,8) ,
66444	 => std_logic_vector(to_unsigned(25,8) ,
66445	 => std_logic_vector(to_unsigned(32,8) ,
66446	 => std_logic_vector(to_unsigned(15,8) ,
66447	 => std_logic_vector(to_unsigned(8,8) ,
66448	 => std_logic_vector(to_unsigned(18,8) ,
66449	 => std_logic_vector(to_unsigned(37,8) ,
66450	 => std_logic_vector(to_unsigned(76,8) ,
66451	 => std_logic_vector(to_unsigned(65,8) ,
66452	 => std_logic_vector(to_unsigned(30,8) ,
66453	 => std_logic_vector(to_unsigned(26,8) ,
66454	 => std_logic_vector(to_unsigned(38,8) ,
66455	 => std_logic_vector(to_unsigned(51,8) ,
66456	 => std_logic_vector(to_unsigned(46,8) ,
66457	 => std_logic_vector(to_unsigned(35,8) ,
66458	 => std_logic_vector(to_unsigned(27,8) ,
66459	 => std_logic_vector(to_unsigned(26,8) ,
66460	 => std_logic_vector(to_unsigned(26,8) ,
66461	 => std_logic_vector(to_unsigned(24,8) ,
66462	 => std_logic_vector(to_unsigned(15,8) ,
66463	 => std_logic_vector(to_unsigned(28,8) ,
66464	 => std_logic_vector(to_unsigned(45,8) ,
66465	 => std_logic_vector(to_unsigned(32,8) ,
66466	 => std_logic_vector(to_unsigned(40,8) ,
66467	 => std_logic_vector(to_unsigned(29,8) ,
66468	 => std_logic_vector(to_unsigned(25,8) ,
66469	 => std_logic_vector(to_unsigned(11,8) ,
66470	 => std_logic_vector(to_unsigned(10,8) ,
66471	 => std_logic_vector(to_unsigned(17,8) ,
66472	 => std_logic_vector(to_unsigned(20,8) ,
66473	 => std_logic_vector(to_unsigned(15,8) ,
66474	 => std_logic_vector(to_unsigned(12,8) ,
66475	 => std_logic_vector(to_unsigned(22,8) ,
66476	 => std_logic_vector(to_unsigned(38,8) ,
66477	 => std_logic_vector(to_unsigned(27,8) ,
66478	 => std_logic_vector(to_unsigned(19,8) ,
66479	 => std_logic_vector(to_unsigned(13,8) ,
66480	 => std_logic_vector(to_unsigned(9,8) ,
66481	 => std_logic_vector(to_unsigned(11,8) ,
66482	 => std_logic_vector(to_unsigned(41,8) ,
66483	 => std_logic_vector(to_unsigned(112,8) ,
66484	 => std_logic_vector(to_unsigned(131,8) ,
66485	 => std_logic_vector(to_unsigned(43,8) ,
66486	 => std_logic_vector(to_unsigned(32,8) ,
66487	 => std_logic_vector(to_unsigned(69,8) ,
66488	 => std_logic_vector(to_unsigned(112,8) ,
66489	 => std_logic_vector(to_unsigned(119,8) ,
66490	 => std_logic_vector(to_unsigned(67,8) ,
66491	 => std_logic_vector(to_unsigned(12,8) ,
66492	 => std_logic_vector(to_unsigned(17,8) ,
66493	 => std_logic_vector(to_unsigned(13,8) ,
66494	 => std_logic_vector(to_unsigned(11,8) ,
66495	 => std_logic_vector(to_unsigned(22,8) ,
66496	 => std_logic_vector(to_unsigned(34,8) ,
66497	 => std_logic_vector(to_unsigned(34,8) ,
66498	 => std_logic_vector(to_unsigned(30,8) ,
66499	 => std_logic_vector(to_unsigned(30,8) ,
66500	 => std_logic_vector(to_unsigned(20,8) ,
66501	 => std_logic_vector(to_unsigned(9,8) ,
66502	 => std_logic_vector(to_unsigned(15,8) ,
66503	 => std_logic_vector(to_unsigned(7,8) ,
66504	 => std_logic_vector(to_unsigned(15,8) ,
66505	 => std_logic_vector(to_unsigned(29,8) ,
66506	 => std_logic_vector(to_unsigned(43,8) ,
66507	 => std_logic_vector(to_unsigned(37,8) ,
66508	 => std_logic_vector(to_unsigned(29,8) ,
66509	 => std_logic_vector(to_unsigned(46,8) ,
66510	 => std_logic_vector(to_unsigned(38,8) ,
66511	 => std_logic_vector(to_unsigned(31,8) ,
66512	 => std_logic_vector(to_unsigned(3,8) ,
66513	 => std_logic_vector(to_unsigned(0,8) ,
66514	 => std_logic_vector(to_unsigned(4,8) ,
66515	 => std_logic_vector(to_unsigned(22,8) ,
66516	 => std_logic_vector(to_unsigned(20,8) ,
66517	 => std_logic_vector(to_unsigned(20,8) ,
66518	 => std_logic_vector(to_unsigned(13,8) ,
66519	 => std_logic_vector(to_unsigned(18,8) ,
66520	 => std_logic_vector(to_unsigned(22,8) ,
66521	 => std_logic_vector(to_unsigned(21,8) ,
66522	 => std_logic_vector(to_unsigned(14,8) ,
66523	 => std_logic_vector(to_unsigned(10,8) ,
66524	 => std_logic_vector(to_unsigned(8,8) ,
66525	 => std_logic_vector(to_unsigned(1,8) ,
66526	 => std_logic_vector(to_unsigned(0,8) ,
66527	 => std_logic_vector(to_unsigned(5,8) ,
66528	 => std_logic_vector(to_unsigned(14,8) ,
66529	 => std_logic_vector(to_unsigned(6,8) ,
66530	 => std_logic_vector(to_unsigned(27,8) ,
66531	 => std_logic_vector(to_unsigned(47,8) ,
66532	 => std_logic_vector(to_unsigned(33,8) ,
66533	 => std_logic_vector(to_unsigned(17,8) ,
66534	 => std_logic_vector(to_unsigned(8,8) ,
66535	 => std_logic_vector(to_unsigned(17,8) ,
66536	 => std_logic_vector(to_unsigned(40,8) ,
66537	 => std_logic_vector(to_unsigned(5,8) ,
66538	 => std_logic_vector(to_unsigned(0,8) ,
66539	 => std_logic_vector(to_unsigned(4,8) ,
66540	 => std_logic_vector(to_unsigned(34,8) ,
66541	 => std_logic_vector(to_unsigned(35,8) ,
66542	 => std_logic_vector(to_unsigned(36,8) ,
66543	 => std_logic_vector(to_unsigned(34,8) ,
66544	 => std_logic_vector(to_unsigned(39,8) ,
66545	 => std_logic_vector(to_unsigned(37,8) ,
66546	 => std_logic_vector(to_unsigned(23,8) ,
66547	 => std_logic_vector(to_unsigned(17,8) ,
66548	 => std_logic_vector(to_unsigned(24,8) ,
66549	 => std_logic_vector(to_unsigned(35,8) ,
66550	 => std_logic_vector(to_unsigned(39,8) ,
66551	 => std_logic_vector(to_unsigned(40,8) ,
66552	 => std_logic_vector(to_unsigned(37,8) ,
66553	 => std_logic_vector(to_unsigned(37,8) ,
66554	 => std_logic_vector(to_unsigned(40,8) ,
66555	 => std_logic_vector(to_unsigned(27,8) ,
66556	 => std_logic_vector(to_unsigned(25,8) ,
66557	 => std_logic_vector(to_unsigned(81,8) ,
66558	 => std_logic_vector(to_unsigned(101,8) ,
66559	 => std_logic_vector(to_unsigned(99,8) ,
66560	 => std_logic_vector(to_unsigned(96,8) ,
66561	 => std_logic_vector(to_unsigned(97,8) ,
66562	 => std_logic_vector(to_unsigned(104,8) ,
66563	 => std_logic_vector(to_unsigned(114,8) ,
66564	 => std_logic_vector(to_unsigned(88,8) ,
66565	 => std_logic_vector(to_unsigned(78,8) ,
66566	 => std_logic_vector(to_unsigned(118,8) ,
66567	 => std_logic_vector(to_unsigned(108,8) ,
66568	 => std_logic_vector(to_unsigned(101,8) ,
66569	 => std_logic_vector(to_unsigned(88,8) ,
66570	 => std_logic_vector(to_unsigned(58,8) ,
66571	 => std_logic_vector(to_unsigned(52,8) ,
66572	 => std_logic_vector(to_unsigned(51,8) ,
66573	 => std_logic_vector(to_unsigned(49,8) ,
66574	 => std_logic_vector(to_unsigned(53,8) ,
66575	 => std_logic_vector(to_unsigned(54,8) ,
66576	 => std_logic_vector(to_unsigned(77,8) ,
66577	 => std_logic_vector(to_unsigned(71,8) ,
66578	 => std_logic_vector(to_unsigned(65,8) ,
66579	 => std_logic_vector(to_unsigned(76,8) ,
66580	 => std_logic_vector(to_unsigned(74,8) ,
66581	 => std_logic_vector(to_unsigned(86,8) ,
66582	 => std_logic_vector(to_unsigned(111,8) ,
66583	 => std_logic_vector(to_unsigned(99,8) ,
66584	 => std_logic_vector(to_unsigned(46,8) ,
66585	 => std_logic_vector(to_unsigned(39,8) ,
66586	 => std_logic_vector(to_unsigned(42,8) ,
66587	 => std_logic_vector(to_unsigned(36,8) ,
66588	 => std_logic_vector(to_unsigned(29,8) ,
66589	 => std_logic_vector(to_unsigned(34,8) ,
66590	 => std_logic_vector(to_unsigned(36,8) ,
66591	 => std_logic_vector(to_unsigned(31,8) ,
66592	 => std_logic_vector(to_unsigned(29,8) ,
66593	 => std_logic_vector(to_unsigned(25,8) ,
66594	 => std_logic_vector(to_unsigned(24,8) ,
66595	 => std_logic_vector(to_unsigned(25,8) ,
66596	 => std_logic_vector(to_unsigned(31,8) ,
66597	 => std_logic_vector(to_unsigned(29,8) ,
66598	 => std_logic_vector(to_unsigned(24,8) ,
66599	 => std_logic_vector(to_unsigned(37,8) ,
66600	 => std_logic_vector(to_unsigned(28,8) ,
66601	 => std_logic_vector(to_unsigned(18,8) ,
66602	 => std_logic_vector(to_unsigned(17,8) ,
66603	 => std_logic_vector(to_unsigned(24,8) ,
66604	 => std_logic_vector(to_unsigned(35,8) ,
66605	 => std_logic_vector(to_unsigned(35,8) ,
66606	 => std_logic_vector(to_unsigned(44,8) ,
66607	 => std_logic_vector(to_unsigned(64,8) ,
66608	 => std_logic_vector(to_unsigned(64,8) ,
66609	 => std_logic_vector(to_unsigned(52,8) ,
66610	 => std_logic_vector(to_unsigned(45,8) ,
66611	 => std_logic_vector(to_unsigned(45,8) ,
66612	 => std_logic_vector(to_unsigned(36,8) ,
66613	 => std_logic_vector(to_unsigned(31,8) ,
66614	 => std_logic_vector(to_unsigned(41,8) ,
66615	 => std_logic_vector(to_unsigned(60,8) ,
66616	 => std_logic_vector(to_unsigned(69,8) ,
66617	 => std_logic_vector(to_unsigned(67,8) ,
66618	 => std_logic_vector(to_unsigned(61,8) ,
66619	 => std_logic_vector(to_unsigned(54,8) ,
66620	 => std_logic_vector(to_unsigned(59,8) ,
66621	 => std_logic_vector(to_unsigned(76,8) ,
66622	 => std_logic_vector(to_unsigned(81,8) ,
66623	 => std_logic_vector(to_unsigned(73,8) ,
66624	 => std_logic_vector(to_unsigned(81,8) ,
66625	 => std_logic_vector(to_unsigned(91,8) ,
66626	 => std_logic_vector(to_unsigned(92,8) ,
66627	 => std_logic_vector(to_unsigned(101,8) ,
66628	 => std_logic_vector(to_unsigned(104,8) ,
66629	 => std_logic_vector(to_unsigned(100,8) ,
66630	 => std_logic_vector(to_unsigned(101,8) ,
66631	 => std_logic_vector(to_unsigned(107,8) ,
66632	 => std_logic_vector(to_unsigned(87,8) ,
66633	 => std_logic_vector(to_unsigned(99,8) ,
66634	 => std_logic_vector(to_unsigned(115,8) ,
66635	 => std_logic_vector(to_unsigned(114,8) ,
66636	 => std_logic_vector(to_unsigned(114,8) ,
66637	 => std_logic_vector(to_unsigned(114,8) ,
66638	 => std_logic_vector(to_unsigned(109,8) ,
66639	 => std_logic_vector(to_unsigned(97,8) ,
66640	 => std_logic_vector(to_unsigned(93,8) ,
66641	 => std_logic_vector(to_unsigned(96,8) ,
66642	 => std_logic_vector(to_unsigned(105,8) ,
66643	 => std_logic_vector(to_unsigned(99,8) ,
66644	 => std_logic_vector(to_unsigned(62,8) ,
66645	 => std_logic_vector(to_unsigned(61,8) ,
66646	 => std_logic_vector(to_unsigned(60,8) ,
66647	 => std_logic_vector(to_unsigned(54,8) ,
66648	 => std_logic_vector(to_unsigned(99,8) ,
66649	 => std_logic_vector(to_unsigned(67,8) ,
66650	 => std_logic_vector(to_unsigned(23,8) ,
66651	 => std_logic_vector(to_unsigned(30,8) ,
66652	 => std_logic_vector(to_unsigned(43,8) ,
66653	 => std_logic_vector(to_unsigned(60,8) ,
66654	 => std_logic_vector(to_unsigned(59,8) ,
66655	 => std_logic_vector(to_unsigned(51,8) ,
66656	 => std_logic_vector(to_unsigned(51,8) ,
66657	 => std_logic_vector(to_unsigned(55,8) ,
66658	 => std_logic_vector(to_unsigned(53,8) ,
66659	 => std_logic_vector(to_unsigned(56,8) ,
66660	 => std_logic_vector(to_unsigned(70,8) ,
66661	 => std_logic_vector(to_unsigned(44,8) ,
66662	 => std_logic_vector(to_unsigned(43,8) ,
66663	 => std_logic_vector(to_unsigned(27,8) ,
66664	 => std_logic_vector(to_unsigned(22,8) ,
66665	 => std_logic_vector(to_unsigned(21,8) ,
66666	 => std_logic_vector(to_unsigned(18,8) ,
66667	 => std_logic_vector(to_unsigned(17,8) ,
66668	 => std_logic_vector(to_unsigned(18,8) ,
66669	 => std_logic_vector(to_unsigned(43,8) ,
66670	 => std_logic_vector(to_unsigned(62,8) ,
66671	 => std_logic_vector(to_unsigned(45,8) ,
66672	 => std_logic_vector(to_unsigned(41,8) ,
66673	 => std_logic_vector(to_unsigned(112,8) ,
66674	 => std_logic_vector(to_unsigned(122,8) ,
66675	 => std_logic_vector(to_unsigned(39,8) ,
66676	 => std_logic_vector(to_unsigned(43,8) ,
66677	 => std_logic_vector(to_unsigned(55,8) ,
66678	 => std_logic_vector(to_unsigned(71,8) ,
66679	 => std_logic_vector(to_unsigned(109,8) ,
66680	 => std_logic_vector(to_unsigned(63,8) ,
66681	 => std_logic_vector(to_unsigned(42,8) ,
66682	 => std_logic_vector(to_unsigned(46,8) ,
66683	 => std_logic_vector(to_unsigned(53,8) ,
66684	 => std_logic_vector(to_unsigned(47,8) ,
66685	 => std_logic_vector(to_unsigned(44,8) ,
66686	 => std_logic_vector(to_unsigned(56,8) ,
66687	 => std_logic_vector(to_unsigned(48,8) ,
66688	 => std_logic_vector(to_unsigned(52,8) ,
66689	 => std_logic_vector(to_unsigned(57,8) ,
66690	 => std_logic_vector(to_unsigned(48,8) ,
66691	 => std_logic_vector(to_unsigned(56,8) ,
66692	 => std_logic_vector(to_unsigned(60,8) ,
66693	 => std_logic_vector(to_unsigned(70,8) ,
66694	 => std_logic_vector(to_unsigned(70,8) ,
66695	 => std_logic_vector(to_unsigned(71,8) ,
66696	 => std_logic_vector(to_unsigned(68,8) ,
66697	 => std_logic_vector(to_unsigned(71,8) ,
66698	 => std_logic_vector(to_unsigned(95,8) ,
66699	 => std_logic_vector(to_unsigned(46,8) ,
66700	 => std_logic_vector(to_unsigned(17,8) ,
66701	 => std_logic_vector(to_unsigned(17,8) ,
66702	 => std_logic_vector(to_unsigned(22,8) ,
66703	 => std_logic_vector(to_unsigned(57,8) ,
66704	 => std_logic_vector(to_unsigned(92,8) ,
66705	 => std_logic_vector(to_unsigned(74,8) ,
66706	 => std_logic_vector(to_unsigned(47,8) ,
66707	 => std_logic_vector(to_unsigned(29,8) ,
66708	 => std_logic_vector(to_unsigned(37,8) ,
66709	 => std_logic_vector(to_unsigned(74,8) ,
66710	 => std_logic_vector(to_unsigned(81,8) ,
66711	 => std_logic_vector(to_unsigned(78,8) ,
66712	 => std_logic_vector(to_unsigned(77,8) ,
66713	 => std_logic_vector(to_unsigned(60,8) ,
66714	 => std_logic_vector(to_unsigned(59,8) ,
66715	 => std_logic_vector(to_unsigned(67,8) ,
66716	 => std_logic_vector(to_unsigned(35,8) ,
66717	 => std_logic_vector(to_unsigned(11,8) ,
66718	 => std_logic_vector(to_unsigned(9,8) ,
66719	 => std_logic_vector(to_unsigned(5,8) ,
66720	 => std_logic_vector(to_unsigned(12,8) ,
66721	 => std_logic_vector(to_unsigned(17,8) ,
66722	 => std_logic_vector(to_unsigned(34,8) ,
66723	 => std_logic_vector(to_unsigned(43,8) ,
66724	 => std_logic_vector(to_unsigned(24,8) ,
66725	 => std_logic_vector(to_unsigned(28,8) ,
66726	 => std_logic_vector(to_unsigned(19,8) ,
66727	 => std_logic_vector(to_unsigned(10,8) ,
66728	 => std_logic_vector(to_unsigned(18,8) ,
66729	 => std_logic_vector(to_unsigned(49,8) ,
66730	 => std_logic_vector(to_unsigned(28,8) ,
66731	 => std_logic_vector(to_unsigned(22,8) ,
66732	 => std_logic_vector(to_unsigned(56,8) ,
66733	 => std_logic_vector(to_unsigned(54,8) ,
66734	 => std_logic_vector(to_unsigned(24,8) ,
66735	 => std_logic_vector(to_unsigned(30,8) ,
66736	 => std_logic_vector(to_unsigned(27,8) ,
66737	 => std_logic_vector(to_unsigned(41,8) ,
66738	 => std_logic_vector(to_unsigned(36,8) ,
66739	 => std_logic_vector(to_unsigned(24,8) ,
66740	 => std_logic_vector(to_unsigned(51,8) ,
66741	 => std_logic_vector(to_unsigned(19,8) ,
66742	 => std_logic_vector(to_unsigned(9,8) ,
66743	 => std_logic_vector(to_unsigned(13,8) ,
66744	 => std_logic_vector(to_unsigned(11,8) ,
66745	 => std_logic_vector(to_unsigned(11,8) ,
66746	 => std_logic_vector(to_unsigned(32,8) ,
66747	 => std_logic_vector(to_unsigned(66,8) ,
66748	 => std_logic_vector(to_unsigned(68,8) ,
66749	 => std_logic_vector(to_unsigned(60,8) ,
66750	 => std_logic_vector(to_unsigned(45,8) ,
66751	 => std_logic_vector(to_unsigned(48,8) ,
66752	 => std_logic_vector(to_unsigned(40,8) ,
66753	 => std_logic_vector(to_unsigned(25,8) ,
66754	 => std_logic_vector(to_unsigned(30,8) ,
66755	 => std_logic_vector(to_unsigned(45,8) ,
66756	 => std_logic_vector(to_unsigned(47,8) ,
66757	 => std_logic_vector(to_unsigned(53,8) ,
66758	 => std_logic_vector(to_unsigned(63,8) ,
66759	 => std_logic_vector(to_unsigned(58,8) ,
66760	 => std_logic_vector(to_unsigned(46,8) ,
66761	 => std_logic_vector(to_unsigned(37,8) ,
66762	 => std_logic_vector(to_unsigned(24,8) ,
66763	 => std_logic_vector(to_unsigned(17,8) ,
66764	 => std_logic_vector(to_unsigned(20,8) ,
66765	 => std_logic_vector(to_unsigned(21,8) ,
66766	 => std_logic_vector(to_unsigned(12,8) ,
66767	 => std_logic_vector(to_unsigned(12,8) ,
66768	 => std_logic_vector(to_unsigned(24,8) ,
66769	 => std_logic_vector(to_unsigned(45,8) ,
66770	 => std_logic_vector(to_unsigned(82,8) ,
66771	 => std_logic_vector(to_unsigned(74,8) ,
66772	 => std_logic_vector(to_unsigned(25,8) ,
66773	 => std_logic_vector(to_unsigned(24,8) ,
66774	 => std_logic_vector(to_unsigned(27,8) ,
66775	 => std_logic_vector(to_unsigned(22,8) ,
66776	 => std_logic_vector(to_unsigned(27,8) ,
66777	 => std_logic_vector(to_unsigned(31,8) ,
66778	 => std_logic_vector(to_unsigned(24,8) ,
66779	 => std_logic_vector(to_unsigned(22,8) ,
66780	 => std_logic_vector(to_unsigned(42,8) ,
66781	 => std_logic_vector(to_unsigned(35,8) ,
66782	 => std_logic_vector(to_unsigned(21,8) ,
66783	 => std_logic_vector(to_unsigned(26,8) ,
66784	 => std_logic_vector(to_unsigned(34,8) ,
66785	 => std_logic_vector(to_unsigned(27,8) ,
66786	 => std_logic_vector(to_unsigned(36,8) ,
66787	 => std_logic_vector(to_unsigned(35,8) ,
66788	 => std_logic_vector(to_unsigned(30,8) ,
66789	 => std_logic_vector(to_unsigned(19,8) ,
66790	 => std_logic_vector(to_unsigned(19,8) ,
66791	 => std_logic_vector(to_unsigned(19,8) ,
66792	 => std_logic_vector(to_unsigned(20,8) ,
66793	 => std_logic_vector(to_unsigned(20,8) ,
66794	 => std_logic_vector(to_unsigned(15,8) ,
66795	 => std_logic_vector(to_unsigned(16,8) ,
66796	 => std_logic_vector(to_unsigned(21,8) ,
66797	 => std_logic_vector(to_unsigned(19,8) ,
66798	 => std_logic_vector(to_unsigned(17,8) ,
66799	 => std_logic_vector(to_unsigned(20,8) ,
66800	 => std_logic_vector(to_unsigned(23,8) ,
66801	 => std_logic_vector(to_unsigned(17,8) ,
66802	 => std_logic_vector(to_unsigned(31,8) ,
66803	 => std_logic_vector(to_unsigned(70,8) ,
66804	 => std_logic_vector(to_unsigned(69,8) ,
66805	 => std_logic_vector(to_unsigned(43,8) ,
66806	 => std_logic_vector(to_unsigned(45,8) ,
66807	 => std_logic_vector(to_unsigned(52,8) ,
66808	 => std_logic_vector(to_unsigned(111,8) ,
66809	 => std_logic_vector(to_unsigned(139,8) ,
66810	 => std_logic_vector(to_unsigned(72,8) ,
66811	 => std_logic_vector(to_unsigned(16,8) ,
66812	 => std_logic_vector(to_unsigned(13,8) ,
66813	 => std_logic_vector(to_unsigned(7,8) ,
66814	 => std_logic_vector(to_unsigned(18,8) ,
66815	 => std_logic_vector(to_unsigned(17,8) ,
66816	 => std_logic_vector(to_unsigned(28,8) ,
66817	 => std_logic_vector(to_unsigned(23,8) ,
66818	 => std_logic_vector(to_unsigned(24,8) ,
66819	 => std_logic_vector(to_unsigned(19,8) ,
66820	 => std_logic_vector(to_unsigned(13,8) ,
66821	 => std_logic_vector(to_unsigned(12,8) ,
66822	 => std_logic_vector(to_unsigned(12,8) ,
66823	 => std_logic_vector(to_unsigned(8,8) ,
66824	 => std_logic_vector(to_unsigned(18,8) ,
66825	 => std_logic_vector(to_unsigned(59,8) ,
66826	 => std_logic_vector(to_unsigned(65,8) ,
66827	 => std_logic_vector(to_unsigned(26,8) ,
66828	 => std_logic_vector(to_unsigned(35,8) ,
66829	 => std_logic_vector(to_unsigned(42,8) ,
66830	 => std_logic_vector(to_unsigned(34,8) ,
66831	 => std_logic_vector(to_unsigned(43,8) ,
66832	 => std_logic_vector(to_unsigned(2,8) ,
66833	 => std_logic_vector(to_unsigned(0,8) ,
66834	 => std_logic_vector(to_unsigned(1,8) ,
66835	 => std_logic_vector(to_unsigned(4,8) ,
66836	 => std_logic_vector(to_unsigned(7,8) ,
66837	 => std_logic_vector(to_unsigned(8,8) ,
66838	 => std_logic_vector(to_unsigned(7,8) ,
66839	 => std_logic_vector(to_unsigned(11,8) ,
66840	 => std_logic_vector(to_unsigned(13,8) ,
66841	 => std_logic_vector(to_unsigned(14,8) ,
66842	 => std_logic_vector(to_unsigned(17,8) ,
66843	 => std_logic_vector(to_unsigned(18,8) ,
66844	 => std_logic_vector(to_unsigned(9,8) ,
66845	 => std_logic_vector(to_unsigned(1,8) ,
66846	 => std_logic_vector(to_unsigned(0,8) ,
66847	 => std_logic_vector(to_unsigned(5,8) ,
66848	 => std_logic_vector(to_unsigned(16,8) ,
66849	 => std_logic_vector(to_unsigned(8,8) ,
66850	 => std_logic_vector(to_unsigned(12,8) ,
66851	 => std_logic_vector(to_unsigned(18,8) ,
66852	 => std_logic_vector(to_unsigned(22,8) ,
66853	 => std_logic_vector(to_unsigned(13,8) ,
66854	 => std_logic_vector(to_unsigned(10,8) ,
66855	 => std_logic_vector(to_unsigned(15,8) ,
66856	 => std_logic_vector(to_unsigned(51,8) ,
66857	 => std_logic_vector(to_unsigned(16,8) ,
66858	 => std_logic_vector(to_unsigned(0,8) ,
66859	 => std_logic_vector(to_unsigned(1,8) ,
66860	 => std_logic_vector(to_unsigned(14,8) ,
66861	 => std_logic_vector(to_unsigned(35,8) ,
66862	 => std_logic_vector(to_unsigned(29,8) ,
66863	 => std_logic_vector(to_unsigned(65,8) ,
66864	 => std_logic_vector(to_unsigned(79,8) ,
66865	 => std_logic_vector(to_unsigned(43,8) ,
66866	 => std_logic_vector(to_unsigned(31,8) ,
66867	 => std_logic_vector(to_unsigned(29,8) ,
66868	 => std_logic_vector(to_unsigned(37,8) ,
66869	 => std_logic_vector(to_unsigned(41,8) ,
66870	 => std_logic_vector(to_unsigned(33,8) ,
66871	 => std_logic_vector(to_unsigned(37,8) ,
66872	 => std_logic_vector(to_unsigned(36,8) ,
66873	 => std_logic_vector(to_unsigned(36,8) ,
66874	 => std_logic_vector(to_unsigned(41,8) ,
66875	 => std_logic_vector(to_unsigned(34,8) ,
66876	 => std_logic_vector(to_unsigned(25,8) ,
66877	 => std_logic_vector(to_unsigned(35,8) ,
66878	 => std_logic_vector(to_unsigned(63,8) ,
66879	 => std_logic_vector(to_unsigned(66,8) ,
66880	 => std_logic_vector(to_unsigned(60,8) ,
66881	 => std_logic_vector(to_unsigned(131,8) ,
66882	 => std_logic_vector(to_unsigned(122,8) ,
66883	 => std_logic_vector(to_unsigned(122,8) ,
66884	 => std_logic_vector(to_unsigned(96,8) ,
66885	 => std_logic_vector(to_unsigned(92,8) ,
66886	 => std_logic_vector(to_unsigned(118,8) ,
66887	 => std_logic_vector(to_unsigned(92,8) ,
66888	 => std_logic_vector(to_unsigned(64,8) ,
66889	 => std_logic_vector(to_unsigned(63,8) ,
66890	 => std_logic_vector(to_unsigned(67,8) ,
66891	 => std_logic_vector(to_unsigned(69,8) ,
66892	 => std_logic_vector(to_unsigned(70,8) ,
66893	 => std_logic_vector(to_unsigned(71,8) ,
66894	 => std_logic_vector(to_unsigned(51,8) ,
66895	 => std_logic_vector(to_unsigned(37,8) ,
66896	 => std_logic_vector(to_unsigned(71,8) ,
66897	 => std_logic_vector(to_unsigned(82,8) ,
66898	 => std_logic_vector(to_unsigned(68,8) ,
66899	 => std_logic_vector(to_unsigned(59,8) ,
66900	 => std_logic_vector(to_unsigned(43,8) ,
66901	 => std_logic_vector(to_unsigned(64,8) ,
66902	 => std_logic_vector(to_unsigned(103,8) ,
66903	 => std_logic_vector(to_unsigned(86,8) ,
66904	 => std_logic_vector(to_unsigned(43,8) ,
66905	 => std_logic_vector(to_unsigned(39,8) ,
66906	 => std_logic_vector(to_unsigned(33,8) ,
66907	 => std_logic_vector(to_unsigned(32,8) ,
66908	 => std_logic_vector(to_unsigned(35,8) ,
66909	 => std_logic_vector(to_unsigned(39,8) ,
66910	 => std_logic_vector(to_unsigned(32,8) ,
66911	 => std_logic_vector(to_unsigned(30,8) ,
66912	 => std_logic_vector(to_unsigned(30,8) ,
66913	 => std_logic_vector(to_unsigned(27,8) ,
66914	 => std_logic_vector(to_unsigned(28,8) ,
66915	 => std_logic_vector(to_unsigned(27,8) ,
66916	 => std_logic_vector(to_unsigned(31,8) ,
66917	 => std_logic_vector(to_unsigned(29,8) ,
66918	 => std_logic_vector(to_unsigned(30,8) ,
66919	 => std_logic_vector(to_unsigned(29,8) ,
66920	 => std_logic_vector(to_unsigned(30,8) ,
66921	 => std_logic_vector(to_unsigned(24,8) ,
66922	 => std_logic_vector(to_unsigned(17,8) ,
66923	 => std_logic_vector(to_unsigned(19,8) ,
66924	 => std_logic_vector(to_unsigned(29,8) ,
66925	 => std_logic_vector(to_unsigned(54,8) ,
66926	 => std_logic_vector(to_unsigned(70,8) ,
66927	 => std_logic_vector(to_unsigned(61,8) ,
66928	 => std_logic_vector(to_unsigned(71,8) ,
66929	 => std_logic_vector(to_unsigned(84,8) ,
66930	 => std_logic_vector(to_unsigned(74,8) ,
66931	 => std_logic_vector(to_unsigned(51,8) ,
66932	 => std_logic_vector(to_unsigned(42,8) ,
66933	 => std_logic_vector(to_unsigned(39,8) ,
66934	 => std_logic_vector(to_unsigned(41,8) ,
66935	 => std_logic_vector(to_unsigned(56,8) ,
66936	 => std_logic_vector(to_unsigned(54,8) ,
66937	 => std_logic_vector(to_unsigned(60,8) ,
66938	 => std_logic_vector(to_unsigned(62,8) ,
66939	 => std_logic_vector(to_unsigned(62,8) ,
66940	 => std_logic_vector(to_unsigned(63,8) ,
66941	 => std_logic_vector(to_unsigned(62,8) ,
66942	 => std_logic_vector(to_unsigned(68,8) ,
66943	 => std_logic_vector(to_unsigned(61,8) ,
66944	 => std_logic_vector(to_unsigned(66,8) ,
66945	 => std_logic_vector(to_unsigned(81,8) ,
66946	 => std_logic_vector(to_unsigned(101,8) ,
66947	 => std_logic_vector(to_unsigned(104,8) ,
66948	 => std_logic_vector(to_unsigned(104,8) ,
66949	 => std_logic_vector(to_unsigned(105,8) ,
66950	 => std_logic_vector(to_unsigned(104,8) ,
66951	 => std_logic_vector(to_unsigned(100,8) ,
66952	 => std_logic_vector(to_unsigned(87,8) ,
66953	 => std_logic_vector(to_unsigned(91,8) ,
66954	 => std_logic_vector(to_unsigned(99,8) ,
66955	 => std_logic_vector(to_unsigned(109,8) ,
66956	 => std_logic_vector(to_unsigned(114,8) ,
66957	 => std_logic_vector(to_unsigned(109,8) ,
66958	 => std_logic_vector(to_unsigned(115,8) ,
66959	 => std_logic_vector(to_unsigned(95,8) ,
66960	 => std_logic_vector(to_unsigned(82,8) ,
66961	 => std_logic_vector(to_unsigned(99,8) ,
66962	 => std_logic_vector(to_unsigned(112,8) ,
66963	 => std_logic_vector(to_unsigned(111,8) ,
66964	 => std_logic_vector(to_unsigned(92,8) ,
66965	 => std_logic_vector(to_unsigned(90,8) ,
66966	 => std_logic_vector(to_unsigned(57,8) ,
66967	 => std_logic_vector(to_unsigned(64,8) ,
66968	 => std_logic_vector(to_unsigned(71,8) ,
66969	 => std_logic_vector(to_unsigned(32,8) ,
66970	 => std_logic_vector(to_unsigned(17,8) ,
66971	 => std_logic_vector(to_unsigned(28,8) ,
66972	 => std_logic_vector(to_unsigned(50,8) ,
66973	 => std_logic_vector(to_unsigned(54,8) ,
66974	 => std_logic_vector(to_unsigned(50,8) ,
66975	 => std_logic_vector(to_unsigned(48,8) ,
66976	 => std_logic_vector(to_unsigned(49,8) ,
66977	 => std_logic_vector(to_unsigned(49,8) ,
66978	 => std_logic_vector(to_unsigned(48,8) ,
66979	 => std_logic_vector(to_unsigned(52,8) ,
66980	 => std_logic_vector(to_unsigned(51,8) ,
66981	 => std_logic_vector(to_unsigned(49,8) ,
66982	 => std_logic_vector(to_unsigned(46,8) ,
66983	 => std_logic_vector(to_unsigned(28,8) ,
66984	 => std_logic_vector(to_unsigned(24,8) ,
66985	 => std_logic_vector(to_unsigned(20,8) ,
66986	 => std_logic_vector(to_unsigned(18,8) ,
66987	 => std_logic_vector(to_unsigned(15,8) ,
66988	 => std_logic_vector(to_unsigned(15,8) ,
66989	 => std_logic_vector(to_unsigned(40,8) ,
66990	 => std_logic_vector(to_unsigned(81,8) ,
66991	 => std_logic_vector(to_unsigned(62,8) ,
66992	 => std_logic_vector(to_unsigned(40,8) ,
66993	 => std_logic_vector(to_unsigned(47,8) ,
66994	 => std_logic_vector(to_unsigned(47,8) ,
66995	 => std_logic_vector(to_unsigned(39,8) ,
66996	 => std_logic_vector(to_unsigned(52,8) ,
66997	 => std_logic_vector(to_unsigned(48,8) ,
66998	 => std_logic_vector(to_unsigned(73,8) ,
66999	 => std_logic_vector(to_unsigned(130,8) ,
67000	 => std_logic_vector(to_unsigned(59,8) ,
67001	 => std_logic_vector(to_unsigned(32,8) ,
67002	 => std_logic_vector(to_unsigned(44,8) ,
67003	 => std_logic_vector(to_unsigned(68,8) ,
67004	 => std_logic_vector(to_unsigned(50,8) ,
67005	 => std_logic_vector(to_unsigned(56,8) ,
67006	 => std_logic_vector(to_unsigned(65,8) ,
67007	 => std_logic_vector(to_unsigned(56,8) ,
67008	 => std_logic_vector(to_unsigned(52,8) ,
67009	 => std_logic_vector(to_unsigned(53,8) ,
67010	 => std_logic_vector(to_unsigned(53,8) ,
67011	 => std_logic_vector(to_unsigned(58,8) ,
67012	 => std_logic_vector(to_unsigned(57,8) ,
67013	 => std_logic_vector(to_unsigned(68,8) ,
67014	 => std_logic_vector(to_unsigned(90,8) ,
67015	 => std_logic_vector(to_unsigned(92,8) ,
67016	 => std_logic_vector(to_unsigned(92,8) ,
67017	 => std_logic_vector(to_unsigned(108,8) ,
67018	 => std_logic_vector(to_unsigned(116,8) ,
67019	 => std_logic_vector(to_unsigned(69,8) ,
67020	 => std_logic_vector(to_unsigned(29,8) ,
67021	 => std_logic_vector(to_unsigned(29,8) ,
67022	 => std_logic_vector(to_unsigned(24,8) ,
67023	 => std_logic_vector(to_unsigned(40,8) ,
67024	 => std_logic_vector(to_unsigned(45,8) ,
67025	 => std_logic_vector(to_unsigned(50,8) ,
67026	 => std_logic_vector(to_unsigned(68,8) ,
67027	 => std_logic_vector(to_unsigned(69,8) ,
67028	 => std_logic_vector(to_unsigned(56,8) ,
67029	 => std_logic_vector(to_unsigned(71,8) ,
67030	 => std_logic_vector(to_unsigned(70,8) ,
67031	 => std_logic_vector(to_unsigned(67,8) ,
67032	 => std_logic_vector(to_unsigned(67,8) ,
67033	 => std_logic_vector(to_unsigned(78,8) ,
67034	 => std_logic_vector(to_unsigned(73,8) ,
67035	 => std_logic_vector(to_unsigned(71,8) ,
67036	 => std_logic_vector(to_unsigned(39,8) ,
67037	 => std_logic_vector(to_unsigned(10,8) ,
67038	 => std_logic_vector(to_unsigned(8,8) ,
67039	 => std_logic_vector(to_unsigned(6,8) ,
67040	 => std_logic_vector(to_unsigned(16,8) ,
67041	 => std_logic_vector(to_unsigned(42,8) ,
67042	 => std_logic_vector(to_unsigned(16,8) ,
67043	 => std_logic_vector(to_unsigned(9,8) ,
67044	 => std_logic_vector(to_unsigned(30,8) ,
67045	 => std_logic_vector(to_unsigned(23,8) ,
67046	 => std_logic_vector(to_unsigned(14,8) ,
67047	 => std_logic_vector(to_unsigned(12,8) ,
67048	 => std_logic_vector(to_unsigned(16,8) ,
67049	 => std_logic_vector(to_unsigned(43,8) ,
67050	 => std_logic_vector(to_unsigned(33,8) ,
67051	 => std_logic_vector(to_unsigned(43,8) ,
67052	 => std_logic_vector(to_unsigned(58,8) ,
67053	 => std_logic_vector(to_unsigned(37,8) ,
67054	 => std_logic_vector(to_unsigned(32,8) ,
67055	 => std_logic_vector(to_unsigned(30,8) ,
67056	 => std_logic_vector(to_unsigned(35,8) ,
67057	 => std_logic_vector(to_unsigned(41,8) ,
67058	 => std_logic_vector(to_unsigned(28,8) ,
67059	 => std_logic_vector(to_unsigned(50,8) ,
67060	 => std_logic_vector(to_unsigned(67,8) ,
67061	 => std_logic_vector(to_unsigned(11,8) ,
67062	 => std_logic_vector(to_unsigned(8,8) ,
67063	 => std_logic_vector(to_unsigned(11,8) ,
67064	 => std_logic_vector(to_unsigned(10,8) ,
67065	 => std_logic_vector(to_unsigned(15,8) ,
67066	 => std_logic_vector(to_unsigned(39,8) ,
67067	 => std_logic_vector(to_unsigned(37,8) ,
67068	 => std_logic_vector(to_unsigned(30,8) ,
67069	 => std_logic_vector(to_unsigned(40,8) ,
67070	 => std_logic_vector(to_unsigned(37,8) ,
67071	 => std_logic_vector(to_unsigned(44,8) ,
67072	 => std_logic_vector(to_unsigned(62,8) ,
67073	 => std_logic_vector(to_unsigned(72,8) ,
67074	 => std_logic_vector(to_unsigned(66,8) ,
67075	 => std_logic_vector(to_unsigned(50,8) ,
67076	 => std_logic_vector(to_unsigned(44,8) ,
67077	 => std_logic_vector(to_unsigned(63,8) ,
67078	 => std_logic_vector(to_unsigned(109,8) ,
67079	 => std_logic_vector(to_unsigned(96,8) ,
67080	 => std_logic_vector(to_unsigned(51,8) ,
67081	 => std_logic_vector(to_unsigned(44,8) ,
67082	 => std_logic_vector(to_unsigned(23,8) ,
67083	 => std_logic_vector(to_unsigned(10,8) ,
67084	 => std_logic_vector(to_unsigned(25,8) ,
67085	 => std_logic_vector(to_unsigned(33,8) ,
67086	 => std_logic_vector(to_unsigned(18,8) ,
67087	 => std_logic_vector(to_unsigned(8,8) ,
67088	 => std_logic_vector(to_unsigned(24,8) ,
67089	 => std_logic_vector(to_unsigned(26,8) ,
67090	 => std_logic_vector(to_unsigned(30,8) ,
67091	 => std_logic_vector(to_unsigned(39,8) ,
67092	 => std_logic_vector(to_unsigned(23,8) ,
67093	 => std_logic_vector(to_unsigned(25,8) ,
67094	 => std_logic_vector(to_unsigned(27,8) ,
67095	 => std_logic_vector(to_unsigned(25,8) ,
67096	 => std_logic_vector(to_unsigned(22,8) ,
67097	 => std_logic_vector(to_unsigned(24,8) ,
67098	 => std_logic_vector(to_unsigned(27,8) ,
67099	 => std_logic_vector(to_unsigned(18,8) ,
67100	 => std_logic_vector(to_unsigned(30,8) ,
67101	 => std_logic_vector(to_unsigned(28,8) ,
67102	 => std_logic_vector(to_unsigned(19,8) ,
67103	 => std_logic_vector(to_unsigned(17,8) ,
67104	 => std_logic_vector(to_unsigned(36,8) ,
67105	 => std_logic_vector(to_unsigned(41,8) ,
67106	 => std_logic_vector(to_unsigned(35,8) ,
67107	 => std_logic_vector(to_unsigned(34,8) ,
67108	 => std_logic_vector(to_unsigned(33,8) ,
67109	 => std_logic_vector(to_unsigned(18,8) ,
67110	 => std_logic_vector(to_unsigned(10,8) ,
67111	 => std_logic_vector(to_unsigned(23,8) ,
67112	 => std_logic_vector(to_unsigned(31,8) ,
67113	 => std_logic_vector(to_unsigned(24,8) ,
67114	 => std_logic_vector(to_unsigned(21,8) ,
67115	 => std_logic_vector(to_unsigned(22,8) ,
67116	 => std_logic_vector(to_unsigned(20,8) ,
67117	 => std_logic_vector(to_unsigned(16,8) ,
67118	 => std_logic_vector(to_unsigned(18,8) ,
67119	 => std_logic_vector(to_unsigned(22,8) ,
67120	 => std_logic_vector(to_unsigned(29,8) ,
67121	 => std_logic_vector(to_unsigned(24,8) ,
67122	 => std_logic_vector(to_unsigned(15,8) ,
67123	 => std_logic_vector(to_unsigned(14,8) ,
67124	 => std_logic_vector(to_unsigned(22,8) ,
67125	 => std_logic_vector(to_unsigned(78,8) ,
67126	 => std_logic_vector(to_unsigned(61,8) ,
67127	 => std_logic_vector(to_unsigned(51,8) ,
67128	 => std_logic_vector(to_unsigned(116,8) ,
67129	 => std_logic_vector(to_unsigned(133,8) ,
67130	 => std_logic_vector(to_unsigned(71,8) ,
67131	 => std_logic_vector(to_unsigned(16,8) ,
67132	 => std_logic_vector(to_unsigned(16,8) ,
67133	 => std_logic_vector(to_unsigned(13,8) ,
67134	 => std_logic_vector(to_unsigned(15,8) ,
67135	 => std_logic_vector(to_unsigned(12,8) ,
67136	 => std_logic_vector(to_unsigned(20,8) ,
67137	 => std_logic_vector(to_unsigned(14,8) ,
67138	 => std_logic_vector(to_unsigned(22,8) ,
67139	 => std_logic_vector(to_unsigned(8,8) ,
67140	 => std_logic_vector(to_unsigned(16,8) ,
67141	 => std_logic_vector(to_unsigned(24,8) ,
67142	 => std_logic_vector(to_unsigned(16,8) ,
67143	 => std_logic_vector(to_unsigned(16,8) ,
67144	 => std_logic_vector(to_unsigned(25,8) ,
67145	 => std_logic_vector(to_unsigned(51,8) ,
67146	 => std_logic_vector(to_unsigned(63,8) ,
67147	 => std_logic_vector(to_unsigned(30,8) ,
67148	 => std_logic_vector(to_unsigned(19,8) ,
67149	 => std_logic_vector(to_unsigned(14,8) ,
67150	 => std_logic_vector(to_unsigned(28,8) ,
67151	 => std_logic_vector(to_unsigned(55,8) ,
67152	 => std_logic_vector(to_unsigned(13,8) ,
67153	 => std_logic_vector(to_unsigned(1,8) ,
67154	 => std_logic_vector(to_unsigned(0,8) ,
67155	 => std_logic_vector(to_unsigned(4,8) ,
67156	 => std_logic_vector(to_unsigned(8,8) ,
67157	 => std_logic_vector(to_unsigned(6,8) ,
67158	 => std_logic_vector(to_unsigned(7,8) ,
67159	 => std_logic_vector(to_unsigned(5,8) ,
67160	 => std_logic_vector(to_unsigned(5,8) ,
67161	 => std_logic_vector(to_unsigned(5,8) ,
67162	 => std_logic_vector(to_unsigned(6,8) ,
67163	 => std_logic_vector(to_unsigned(6,8) ,
67164	 => std_logic_vector(to_unsigned(9,8) ,
67165	 => std_logic_vector(to_unsigned(2,8) ,
67166	 => std_logic_vector(to_unsigned(0,8) ,
67167	 => std_logic_vector(to_unsigned(5,8) ,
67168	 => std_logic_vector(to_unsigned(15,8) ,
67169	 => std_logic_vector(to_unsigned(12,8) ,
67170	 => std_logic_vector(to_unsigned(15,8) ,
67171	 => std_logic_vector(to_unsigned(13,8) ,
67172	 => std_logic_vector(to_unsigned(17,8) ,
67173	 => std_logic_vector(to_unsigned(16,8) ,
67174	 => std_logic_vector(to_unsigned(11,8) ,
67175	 => std_logic_vector(to_unsigned(30,8) ,
67176	 => std_logic_vector(to_unsigned(34,8) ,
67177	 => std_logic_vector(to_unsigned(20,8) ,
67178	 => std_logic_vector(to_unsigned(2,8) ,
67179	 => std_logic_vector(to_unsigned(0,8) ,
67180	 => std_logic_vector(to_unsigned(4,8) ,
67181	 => std_logic_vector(to_unsigned(34,8) ,
67182	 => std_logic_vector(to_unsigned(16,8) ,
67183	 => std_logic_vector(to_unsigned(81,8) ,
67184	 => std_logic_vector(to_unsigned(107,8) ,
67185	 => std_logic_vector(to_unsigned(35,8) ,
67186	 => std_logic_vector(to_unsigned(42,8) ,
67187	 => std_logic_vector(to_unsigned(37,8) ,
67188	 => std_logic_vector(to_unsigned(22,8) ,
67189	 => std_logic_vector(to_unsigned(35,8) ,
67190	 => std_logic_vector(to_unsigned(35,8) ,
67191	 => std_logic_vector(to_unsigned(36,8) ,
67192	 => std_logic_vector(to_unsigned(37,8) ,
67193	 => std_logic_vector(to_unsigned(36,8) ,
67194	 => std_logic_vector(to_unsigned(41,8) ,
67195	 => std_logic_vector(to_unsigned(34,8) ,
67196	 => std_logic_vector(to_unsigned(13,8) ,
67197	 => std_logic_vector(to_unsigned(5,8) ,
67198	 => std_logic_vector(to_unsigned(19,8) ,
67199	 => std_logic_vector(to_unsigned(32,8) ,
67200	 => std_logic_vector(to_unsigned(20,8) ,
67201	 => std_logic_vector(to_unsigned(116,8) ,
67202	 => std_logic_vector(to_unsigned(125,8) ,
67203	 => std_logic_vector(to_unsigned(122,8) ,
67204	 => std_logic_vector(to_unsigned(127,8) ,
67205	 => std_logic_vector(to_unsigned(124,8) ,
67206	 => std_logic_vector(to_unsigned(88,8) ,
67207	 => std_logic_vector(to_unsigned(65,8) ,
67208	 => std_logic_vector(to_unsigned(68,8) ,
67209	 => std_logic_vector(to_unsigned(76,8) ,
67210	 => std_logic_vector(to_unsigned(80,8) ,
67211	 => std_logic_vector(to_unsigned(73,8) ,
67212	 => std_logic_vector(to_unsigned(58,8) ,
67213	 => std_logic_vector(to_unsigned(51,8) ,
67214	 => std_logic_vector(to_unsigned(37,8) ,
67215	 => std_logic_vector(to_unsigned(27,8) ,
67216	 => std_logic_vector(to_unsigned(55,8) ,
67217	 => std_logic_vector(to_unsigned(87,8) ,
67218	 => std_logic_vector(to_unsigned(78,8) ,
67219	 => std_logic_vector(to_unsigned(78,8) ,
67220	 => std_logic_vector(to_unsigned(53,8) ,
67221	 => std_logic_vector(to_unsigned(61,8) ,
67222	 => std_logic_vector(to_unsigned(92,8) ,
67223	 => std_logic_vector(to_unsigned(77,8) ,
67224	 => std_logic_vector(to_unsigned(49,8) ,
67225	 => std_logic_vector(to_unsigned(39,8) ,
67226	 => std_logic_vector(to_unsigned(41,8) ,
67227	 => std_logic_vector(to_unsigned(42,8) ,
67228	 => std_logic_vector(to_unsigned(38,8) ,
67229	 => std_logic_vector(to_unsigned(29,8) ,
67230	 => std_logic_vector(to_unsigned(27,8) ,
67231	 => std_logic_vector(to_unsigned(30,8) ,
67232	 => std_logic_vector(to_unsigned(31,8) ,
67233	 => std_logic_vector(to_unsigned(31,8) ,
67234	 => std_logic_vector(to_unsigned(31,8) ,
67235	 => std_logic_vector(to_unsigned(27,8) ,
67236	 => std_logic_vector(to_unsigned(29,8) ,
67237	 => std_logic_vector(to_unsigned(26,8) ,
67238	 => std_logic_vector(to_unsigned(26,8) ,
67239	 => std_logic_vector(to_unsigned(27,8) ,
67240	 => std_logic_vector(to_unsigned(33,8) ,
67241	 => std_logic_vector(to_unsigned(33,8) ,
67242	 => std_logic_vector(to_unsigned(29,8) ,
67243	 => std_logic_vector(to_unsigned(37,8) ,
67244	 => std_logic_vector(to_unsigned(71,8) ,
67245	 => std_logic_vector(to_unsigned(87,8) ,
67246	 => std_logic_vector(to_unsigned(73,8) ,
67247	 => std_logic_vector(to_unsigned(72,8) ,
67248	 => std_logic_vector(to_unsigned(81,8) ,
67249	 => std_logic_vector(to_unsigned(70,8) ,
67250	 => std_logic_vector(to_unsigned(42,8) ,
67251	 => std_logic_vector(to_unsigned(39,8) ,
67252	 => std_logic_vector(to_unsigned(46,8) ,
67253	 => std_logic_vector(to_unsigned(40,8) ,
67254	 => std_logic_vector(to_unsigned(37,8) ,
67255	 => std_logic_vector(to_unsigned(52,8) ,
67256	 => std_logic_vector(to_unsigned(45,8) ,
67257	 => std_logic_vector(to_unsigned(47,8) ,
67258	 => std_logic_vector(to_unsigned(43,8) ,
67259	 => std_logic_vector(to_unsigned(38,8) ,
67260	 => std_logic_vector(to_unsigned(63,8) ,
67261	 => std_logic_vector(to_unsigned(76,8) ,
67262	 => std_logic_vector(to_unsigned(65,8) ,
67263	 => std_logic_vector(to_unsigned(57,8) ,
67264	 => std_logic_vector(to_unsigned(52,8) ,
67265	 => std_logic_vector(to_unsigned(49,8) ,
67266	 => std_logic_vector(to_unsigned(97,8) ,
67267	 => std_logic_vector(to_unsigned(111,8) ,
67268	 => std_logic_vector(to_unsigned(99,8) ,
67269	 => std_logic_vector(to_unsigned(105,8) ,
67270	 => std_logic_vector(to_unsigned(103,8) ,
67271	 => std_logic_vector(to_unsigned(99,8) ,
67272	 => std_logic_vector(to_unsigned(101,8) ,
67273	 => std_logic_vector(to_unsigned(105,8) ,
67274	 => std_logic_vector(to_unsigned(92,8) ,
67275	 => std_logic_vector(to_unsigned(90,8) ,
67276	 => std_logic_vector(to_unsigned(107,8) ,
67277	 => std_logic_vector(to_unsigned(111,8) ,
67278	 => std_logic_vector(to_unsigned(112,8) ,
67279	 => std_logic_vector(to_unsigned(114,8) ,
67280	 => std_logic_vector(to_unsigned(104,8) ,
67281	 => std_logic_vector(to_unsigned(105,8) ,
67282	 => std_logic_vector(to_unsigned(97,8) ,
67283	 => std_logic_vector(to_unsigned(101,8) ,
67284	 => std_logic_vector(to_unsigned(109,8) ,
67285	 => std_logic_vector(to_unsigned(86,8) ,
67286	 => std_logic_vector(to_unsigned(72,8) ,
67287	 => std_logic_vector(to_unsigned(74,8) ,
67288	 => std_logic_vector(to_unsigned(40,8) ,
67289	 => std_logic_vector(to_unsigned(28,8) ,
67290	 => std_logic_vector(to_unsigned(25,8) ,
67291	 => std_logic_vector(to_unsigned(30,8) ,
67292	 => std_logic_vector(to_unsigned(52,8) ,
67293	 => std_logic_vector(to_unsigned(48,8) ,
67294	 => std_logic_vector(to_unsigned(51,8) ,
67295	 => std_logic_vector(to_unsigned(49,8) ,
67296	 => std_logic_vector(to_unsigned(51,8) ,
67297	 => std_logic_vector(to_unsigned(48,8) ,
67298	 => std_logic_vector(to_unsigned(32,8) ,
67299	 => std_logic_vector(to_unsigned(46,8) ,
67300	 => std_logic_vector(to_unsigned(41,8) ,
67301	 => std_logic_vector(to_unsigned(37,8) ,
67302	 => std_logic_vector(to_unsigned(37,8) ,
67303	 => std_logic_vector(to_unsigned(26,8) ,
67304	 => std_logic_vector(to_unsigned(24,8) ,
67305	 => std_logic_vector(to_unsigned(22,8) ,
67306	 => std_logic_vector(to_unsigned(18,8) ,
67307	 => std_logic_vector(to_unsigned(12,8) ,
67308	 => std_logic_vector(to_unsigned(12,8) ,
67309	 => std_logic_vector(to_unsigned(53,8) ,
67310	 => std_logic_vector(to_unsigned(149,8) ,
67311	 => std_logic_vector(to_unsigned(82,8) ,
67312	 => std_logic_vector(to_unsigned(35,8) ,
67313	 => std_logic_vector(to_unsigned(95,8) ,
67314	 => std_logic_vector(to_unsigned(119,8) ,
67315	 => std_logic_vector(to_unsigned(55,8) ,
67316	 => std_logic_vector(to_unsigned(38,8) ,
67317	 => std_logic_vector(to_unsigned(52,8) ,
67318	 => std_logic_vector(to_unsigned(43,8) ,
67319	 => std_logic_vector(to_unsigned(37,8) ,
67320	 => std_logic_vector(to_unsigned(39,8) ,
67321	 => std_logic_vector(to_unsigned(43,8) ,
67322	 => std_logic_vector(to_unsigned(59,8) ,
67323	 => std_logic_vector(to_unsigned(60,8) ,
67324	 => std_logic_vector(to_unsigned(51,8) ,
67325	 => std_logic_vector(to_unsigned(61,8) ,
67326	 => std_logic_vector(to_unsigned(52,8) ,
67327	 => std_logic_vector(to_unsigned(51,8) ,
67328	 => std_logic_vector(to_unsigned(53,8) ,
67329	 => std_logic_vector(to_unsigned(56,8) ,
67330	 => std_logic_vector(to_unsigned(65,8) ,
67331	 => std_logic_vector(to_unsigned(59,8) ,
67332	 => std_logic_vector(to_unsigned(33,8) ,
67333	 => std_logic_vector(to_unsigned(43,8) ,
67334	 => std_logic_vector(to_unsigned(81,8) ,
67335	 => std_logic_vector(to_unsigned(90,8) ,
67336	 => std_logic_vector(to_unsigned(104,8) ,
67337	 => std_logic_vector(to_unsigned(119,8) ,
67338	 => std_logic_vector(to_unsigned(116,8) ,
67339	 => std_logic_vector(to_unsigned(62,8) ,
67340	 => std_logic_vector(to_unsigned(43,8) ,
67341	 => std_logic_vector(to_unsigned(38,8) ,
67342	 => std_logic_vector(to_unsigned(30,8) ,
67343	 => std_logic_vector(to_unsigned(36,8) ,
67344	 => std_logic_vector(to_unsigned(41,8) ,
67345	 => std_logic_vector(to_unsigned(56,8) ,
67346	 => std_logic_vector(to_unsigned(55,8) ,
67347	 => std_logic_vector(to_unsigned(47,8) ,
67348	 => std_logic_vector(to_unsigned(41,8) ,
67349	 => std_logic_vector(to_unsigned(66,8) ,
67350	 => std_logic_vector(to_unsigned(54,8) ,
67351	 => std_logic_vector(to_unsigned(32,8) ,
67352	 => std_logic_vector(to_unsigned(60,8) ,
67353	 => std_logic_vector(to_unsigned(79,8) ,
67354	 => std_logic_vector(to_unsigned(57,8) ,
67355	 => std_logic_vector(to_unsigned(70,8) ,
67356	 => std_logic_vector(to_unsigned(50,8) ,
67357	 => std_logic_vector(to_unsigned(10,8) ,
67358	 => std_logic_vector(to_unsigned(7,8) ,
67359	 => std_logic_vector(to_unsigned(4,8) ,
67360	 => std_logic_vector(to_unsigned(12,8) ,
67361	 => std_logic_vector(to_unsigned(43,8) ,
67362	 => std_logic_vector(to_unsigned(12,8) ,
67363	 => std_logic_vector(to_unsigned(10,8) ,
67364	 => std_logic_vector(to_unsigned(31,8) ,
67365	 => std_logic_vector(to_unsigned(27,8) ,
67366	 => std_logic_vector(to_unsigned(19,8) ,
67367	 => std_logic_vector(to_unsigned(15,8) ,
67368	 => std_logic_vector(to_unsigned(24,8) ,
67369	 => std_logic_vector(to_unsigned(39,8) ,
67370	 => std_logic_vector(to_unsigned(44,8) ,
67371	 => std_logic_vector(to_unsigned(39,8) ,
67372	 => std_logic_vector(to_unsigned(24,8) ,
67373	 => std_logic_vector(to_unsigned(31,8) ,
67374	 => std_logic_vector(to_unsigned(16,8) ,
67375	 => std_logic_vector(to_unsigned(23,8) ,
67376	 => std_logic_vector(to_unsigned(38,8) ,
67377	 => std_logic_vector(to_unsigned(20,8) ,
67378	 => std_logic_vector(to_unsigned(51,8) ,
67379	 => std_logic_vector(to_unsigned(72,8) ,
67380	 => std_logic_vector(to_unsigned(37,8) ,
67381	 => std_logic_vector(to_unsigned(10,8) ,
67382	 => std_logic_vector(to_unsigned(9,8) ,
67383	 => std_logic_vector(to_unsigned(11,8) ,
67384	 => std_logic_vector(to_unsigned(7,8) ,
67385	 => std_logic_vector(to_unsigned(9,8) ,
67386	 => std_logic_vector(to_unsigned(36,8) ,
67387	 => std_logic_vector(to_unsigned(31,8) ,
67388	 => std_logic_vector(to_unsigned(13,8) ,
67389	 => std_logic_vector(to_unsigned(17,8) ,
67390	 => std_logic_vector(to_unsigned(39,8) ,
67391	 => std_logic_vector(to_unsigned(45,8) ,
67392	 => std_logic_vector(to_unsigned(28,8) ,
67393	 => std_logic_vector(to_unsigned(22,8) ,
67394	 => std_logic_vector(to_unsigned(35,8) ,
67395	 => std_logic_vector(to_unsigned(43,8) ,
67396	 => std_logic_vector(to_unsigned(39,8) ,
67397	 => std_logic_vector(to_unsigned(46,8) ,
67398	 => std_logic_vector(to_unsigned(65,8) ,
67399	 => std_logic_vector(to_unsigned(70,8) ,
67400	 => std_logic_vector(to_unsigned(45,8) ,
67401	 => std_logic_vector(to_unsigned(28,8) ,
67402	 => std_logic_vector(to_unsigned(16,8) ,
67403	 => std_logic_vector(to_unsigned(15,8) ,
67404	 => std_logic_vector(to_unsigned(18,8) ,
67405	 => std_logic_vector(to_unsigned(24,8) ,
67406	 => std_logic_vector(to_unsigned(17,8) ,
67407	 => std_logic_vector(to_unsigned(11,8) ,
67408	 => std_logic_vector(to_unsigned(30,8) ,
67409	 => std_logic_vector(to_unsigned(20,8) ,
67410	 => std_logic_vector(to_unsigned(13,8) ,
67411	 => std_logic_vector(to_unsigned(16,8) ,
67412	 => std_logic_vector(to_unsigned(22,8) ,
67413	 => std_logic_vector(to_unsigned(28,8) ,
67414	 => std_logic_vector(to_unsigned(28,8) ,
67415	 => std_logic_vector(to_unsigned(43,8) ,
67416	 => std_logic_vector(to_unsigned(49,8) ,
67417	 => std_logic_vector(to_unsigned(32,8) ,
67418	 => std_logic_vector(to_unsigned(28,8) ,
67419	 => std_logic_vector(to_unsigned(23,8) ,
67420	 => std_logic_vector(to_unsigned(20,8) ,
67421	 => std_logic_vector(to_unsigned(19,8) ,
67422	 => std_logic_vector(to_unsigned(13,8) ,
67423	 => std_logic_vector(to_unsigned(23,8) ,
67424	 => std_logic_vector(to_unsigned(41,8) ,
67425	 => std_logic_vector(to_unsigned(37,8) ,
67426	 => std_logic_vector(to_unsigned(38,8) ,
67427	 => std_logic_vector(to_unsigned(28,8) ,
67428	 => std_logic_vector(to_unsigned(23,8) ,
67429	 => std_logic_vector(to_unsigned(6,8) ,
67430	 => std_logic_vector(to_unsigned(8,8) ,
67431	 => std_logic_vector(to_unsigned(51,8) ,
67432	 => std_logic_vector(to_unsigned(53,8) ,
67433	 => std_logic_vector(to_unsigned(41,8) ,
67434	 => std_logic_vector(to_unsigned(32,8) ,
67435	 => std_logic_vector(to_unsigned(30,8) ,
67436	 => std_logic_vector(to_unsigned(30,8) ,
67437	 => std_logic_vector(to_unsigned(25,8) ,
67438	 => std_logic_vector(to_unsigned(20,8) ,
67439	 => std_logic_vector(to_unsigned(24,8) ,
67440	 => std_logic_vector(to_unsigned(29,8) ,
67441	 => std_logic_vector(to_unsigned(21,8) ,
67442	 => std_logic_vector(to_unsigned(17,8) ,
67443	 => std_logic_vector(to_unsigned(22,8) ,
67444	 => std_logic_vector(to_unsigned(61,8) ,
67445	 => std_logic_vector(to_unsigned(109,8) ,
67446	 => std_logic_vector(to_unsigned(56,8) ,
67447	 => std_logic_vector(to_unsigned(55,8) ,
67448	 => std_logic_vector(to_unsigned(124,8) ,
67449	 => std_logic_vector(to_unsigned(125,8) ,
67450	 => std_logic_vector(to_unsigned(61,8) ,
67451	 => std_logic_vector(to_unsigned(10,8) ,
67452	 => std_logic_vector(to_unsigned(13,8) ,
67453	 => std_logic_vector(to_unsigned(12,8) ,
67454	 => std_logic_vector(to_unsigned(7,8) ,
67455	 => std_logic_vector(to_unsigned(10,8) ,
67456	 => std_logic_vector(to_unsigned(13,8) ,
67457	 => std_logic_vector(to_unsigned(12,8) ,
67458	 => std_logic_vector(to_unsigned(18,8) ,
67459	 => std_logic_vector(to_unsigned(19,8) ,
67460	 => std_logic_vector(to_unsigned(22,8) ,
67461	 => std_logic_vector(to_unsigned(32,8) ,
67462	 => std_logic_vector(to_unsigned(48,8) ,
67463	 => std_logic_vector(to_unsigned(67,8) ,
67464	 => std_logic_vector(to_unsigned(34,8) ,
67465	 => std_logic_vector(to_unsigned(17,8) ,
67466	 => std_logic_vector(to_unsigned(52,8) ,
67467	 => std_logic_vector(to_unsigned(26,8) ,
67468	 => std_logic_vector(to_unsigned(20,8) ,
67469	 => std_logic_vector(to_unsigned(17,8) ,
67470	 => std_logic_vector(to_unsigned(27,8) ,
67471	 => std_logic_vector(to_unsigned(72,8) ,
67472	 => std_logic_vector(to_unsigned(31,8) ,
67473	 => std_logic_vector(to_unsigned(2,8) ,
67474	 => std_logic_vector(to_unsigned(0,8) ,
67475	 => std_logic_vector(to_unsigned(2,8) ,
67476	 => std_logic_vector(to_unsigned(12,8) ,
67477	 => std_logic_vector(to_unsigned(9,8) ,
67478	 => std_logic_vector(to_unsigned(8,8) ,
67479	 => std_logic_vector(to_unsigned(8,8) ,
67480	 => std_logic_vector(to_unsigned(6,8) ,
67481	 => std_logic_vector(to_unsigned(5,8) ,
67482	 => std_logic_vector(to_unsigned(6,8) ,
67483	 => std_logic_vector(to_unsigned(4,8) ,
67484	 => std_logic_vector(to_unsigned(6,8) ,
67485	 => std_logic_vector(to_unsigned(2,8) ,
67486	 => std_logic_vector(to_unsigned(0,8) ,
67487	 => std_logic_vector(to_unsigned(6,8) ,
67488	 => std_logic_vector(to_unsigned(18,8) ,
67489	 => std_logic_vector(to_unsigned(17,8) ,
67490	 => std_logic_vector(to_unsigned(23,8) ,
67491	 => std_logic_vector(to_unsigned(32,8) ,
67492	 => std_logic_vector(to_unsigned(36,8) ,
67493	 => std_logic_vector(to_unsigned(35,8) ,
67494	 => std_logic_vector(to_unsigned(34,8) ,
67495	 => std_logic_vector(to_unsigned(38,8) ,
67496	 => std_logic_vector(to_unsigned(37,8) ,
67497	 => std_logic_vector(to_unsigned(37,8) ,
67498	 => std_logic_vector(to_unsigned(9,8) ,
67499	 => std_logic_vector(to_unsigned(0,8) ,
67500	 => std_logic_vector(to_unsigned(1,8) ,
67501	 => std_logic_vector(to_unsigned(32,8) ,
67502	 => std_logic_vector(to_unsigned(78,8) ,
67503	 => std_logic_vector(to_unsigned(82,8) ,
67504	 => std_logic_vector(to_unsigned(73,8) ,
67505	 => std_logic_vector(to_unsigned(45,8) ,
67506	 => std_logic_vector(to_unsigned(52,8) ,
67507	 => std_logic_vector(to_unsigned(35,8) ,
67508	 => std_logic_vector(to_unsigned(21,8) ,
67509	 => std_logic_vector(to_unsigned(35,8) ,
67510	 => std_logic_vector(to_unsigned(40,8) ,
67511	 => std_logic_vector(to_unsigned(39,8) ,
67512	 => std_logic_vector(to_unsigned(42,8) ,
67513	 => std_logic_vector(to_unsigned(41,8) ,
67514	 => std_logic_vector(to_unsigned(32,8) ,
67515	 => std_logic_vector(to_unsigned(17,8) ,
67516	 => std_logic_vector(to_unsigned(14,8) ,
67517	 => std_logic_vector(to_unsigned(16,8) ,
67518	 => std_logic_vector(to_unsigned(35,8) ,
67519	 => std_logic_vector(to_unsigned(74,8) ,
67520	 => std_logic_vector(to_unsigned(51,8) ,
67521	 => std_logic_vector(to_unsigned(96,8) ,
67522	 => std_logic_vector(to_unsigned(104,8) ,
67523	 => std_logic_vector(to_unsigned(96,8) ,
67524	 => std_logic_vector(to_unsigned(107,8) ,
67525	 => std_logic_vector(to_unsigned(85,8) ,
67526	 => std_logic_vector(to_unsigned(86,8) ,
67527	 => std_logic_vector(to_unsigned(82,8) ,
67528	 => std_logic_vector(to_unsigned(87,8) ,
67529	 => std_logic_vector(to_unsigned(79,8) ,
67530	 => std_logic_vector(to_unsigned(78,8) ,
67531	 => std_logic_vector(to_unsigned(77,8) ,
67532	 => std_logic_vector(to_unsigned(49,8) ,
67533	 => std_logic_vector(to_unsigned(36,8) ,
67534	 => std_logic_vector(to_unsigned(32,8) ,
67535	 => std_logic_vector(to_unsigned(27,8) ,
67536	 => std_logic_vector(to_unsigned(53,8) ,
67537	 => std_logic_vector(to_unsigned(80,8) ,
67538	 => std_logic_vector(to_unsigned(61,8) ,
67539	 => std_logic_vector(to_unsigned(57,8) ,
67540	 => std_logic_vector(to_unsigned(53,8) ,
67541	 => std_logic_vector(to_unsigned(58,8) ,
67542	 => std_logic_vector(to_unsigned(77,8) ,
67543	 => std_logic_vector(to_unsigned(58,8) ,
67544	 => std_logic_vector(to_unsigned(42,8) ,
67545	 => std_logic_vector(to_unsigned(43,8) ,
67546	 => std_logic_vector(to_unsigned(48,8) ,
67547	 => std_logic_vector(to_unsigned(40,8) ,
67548	 => std_logic_vector(to_unsigned(32,8) ,
67549	 => std_logic_vector(to_unsigned(28,8) ,
67550	 => std_logic_vector(to_unsigned(31,8) ,
67551	 => std_logic_vector(to_unsigned(34,8) ,
67552	 => std_logic_vector(to_unsigned(30,8) ,
67553	 => std_logic_vector(to_unsigned(32,8) ,
67554	 => std_logic_vector(to_unsigned(30,8) ,
67555	 => std_logic_vector(to_unsigned(26,8) ,
67556	 => std_logic_vector(to_unsigned(26,8) ,
67557	 => std_logic_vector(to_unsigned(29,8) ,
67558	 => std_logic_vector(to_unsigned(27,8) ,
67559	 => std_logic_vector(to_unsigned(34,8) ,
67560	 => std_logic_vector(to_unsigned(32,8) ,
67561	 => std_logic_vector(to_unsigned(30,8) ,
67562	 => std_logic_vector(to_unsigned(50,8) ,
67563	 => std_logic_vector(to_unsigned(72,8) ,
67564	 => std_logic_vector(to_unsigned(91,8) ,
67565	 => std_logic_vector(to_unsigned(80,8) ,
67566	 => std_logic_vector(to_unsigned(72,8) ,
67567	 => std_logic_vector(to_unsigned(82,8) ,
67568	 => std_logic_vector(to_unsigned(62,8) ,
67569	 => std_logic_vector(to_unsigned(42,8) ,
67570	 => std_logic_vector(to_unsigned(30,8) ,
67571	 => std_logic_vector(to_unsigned(32,8) ,
67572	 => std_logic_vector(to_unsigned(44,8) ,
67573	 => std_logic_vector(to_unsigned(33,8) ,
67574	 => std_logic_vector(to_unsigned(27,8) ,
67575	 => std_logic_vector(to_unsigned(53,8) ,
67576	 => std_logic_vector(to_unsigned(63,8) ,
67577	 => std_logic_vector(to_unsigned(54,8) ,
67578	 => std_logic_vector(to_unsigned(41,8) ,
67579	 => std_logic_vector(to_unsigned(39,8) ,
67580	 => std_logic_vector(to_unsigned(41,8) ,
67581	 => std_logic_vector(to_unsigned(66,8) ,
67582	 => std_logic_vector(to_unsigned(70,8) ,
67583	 => std_logic_vector(to_unsigned(47,8) ,
67584	 => std_logic_vector(to_unsigned(33,8) ,
67585	 => std_logic_vector(to_unsigned(41,8) ,
67586	 => std_logic_vector(to_unsigned(90,8) ,
67587	 => std_logic_vector(to_unsigned(99,8) ,
67588	 => std_logic_vector(to_unsigned(81,8) ,
67589	 => std_logic_vector(to_unsigned(92,8) ,
67590	 => std_logic_vector(to_unsigned(104,8) ,
67591	 => std_logic_vector(to_unsigned(104,8) ,
67592	 => std_logic_vector(to_unsigned(108,8) ,
67593	 => std_logic_vector(to_unsigned(112,8) ,
67594	 => std_logic_vector(to_unsigned(95,8) ,
67595	 => std_logic_vector(to_unsigned(88,8) ,
67596	 => std_logic_vector(to_unsigned(104,8) ,
67597	 => std_logic_vector(to_unsigned(104,8) ,
67598	 => std_logic_vector(to_unsigned(97,8) ,
67599	 => std_logic_vector(to_unsigned(105,8) ,
67600	 => std_logic_vector(to_unsigned(103,8) ,
67601	 => std_logic_vector(to_unsigned(105,8) ,
67602	 => std_logic_vector(to_unsigned(71,8) ,
67603	 => std_logic_vector(to_unsigned(67,8) ,
67604	 => std_logic_vector(to_unsigned(92,8) ,
67605	 => std_logic_vector(to_unsigned(90,8) ,
67606	 => std_logic_vector(to_unsigned(92,8) ,
67607	 => std_logic_vector(to_unsigned(82,8) ,
67608	 => std_logic_vector(to_unsigned(49,8) ,
67609	 => std_logic_vector(to_unsigned(48,8) ,
67610	 => std_logic_vector(to_unsigned(33,8) ,
67611	 => std_logic_vector(to_unsigned(25,8) ,
67612	 => std_logic_vector(to_unsigned(41,8) ,
67613	 => std_logic_vector(to_unsigned(41,8) ,
67614	 => std_logic_vector(to_unsigned(38,8) ,
67615	 => std_logic_vector(to_unsigned(51,8) ,
67616	 => std_logic_vector(to_unsigned(46,8) ,
67617	 => std_logic_vector(to_unsigned(47,8) ,
67618	 => std_logic_vector(to_unsigned(48,8) ,
67619	 => std_logic_vector(to_unsigned(45,8) ,
67620	 => std_logic_vector(to_unsigned(35,8) ,
67621	 => std_logic_vector(to_unsigned(38,8) ,
67622	 => std_logic_vector(to_unsigned(49,8) ,
67623	 => std_logic_vector(to_unsigned(27,8) ,
67624	 => std_logic_vector(to_unsigned(23,8) ,
67625	 => std_logic_vector(to_unsigned(20,8) ,
67626	 => std_logic_vector(to_unsigned(15,8) ,
67627	 => std_logic_vector(to_unsigned(13,8) ,
67628	 => std_logic_vector(to_unsigned(13,8) ,
67629	 => std_logic_vector(to_unsigned(32,8) ,
67630	 => std_logic_vector(to_unsigned(46,8) ,
67631	 => std_logic_vector(to_unsigned(41,8) ,
67632	 => std_logic_vector(to_unsigned(44,8) ,
67633	 => std_logic_vector(to_unsigned(92,8) ,
67634	 => std_logic_vector(to_unsigned(107,8) ,
67635	 => std_logic_vector(to_unsigned(52,8) ,
67636	 => std_logic_vector(to_unsigned(86,8) ,
67637	 => std_logic_vector(to_unsigned(136,8) ,
67638	 => std_logic_vector(to_unsigned(68,8) ,
67639	 => std_logic_vector(to_unsigned(10,8) ,
67640	 => std_logic_vector(to_unsigned(24,8) ,
67641	 => std_logic_vector(to_unsigned(54,8) ,
67642	 => std_logic_vector(to_unsigned(54,8) ,
67643	 => std_logic_vector(to_unsigned(54,8) ,
67644	 => std_logic_vector(to_unsigned(55,8) ,
67645	 => std_logic_vector(to_unsigned(51,8) ,
67646	 => std_logic_vector(to_unsigned(46,8) ,
67647	 => std_logic_vector(to_unsigned(45,8) ,
67648	 => std_logic_vector(to_unsigned(48,8) ,
67649	 => std_logic_vector(to_unsigned(64,8) ,
67650	 => std_logic_vector(to_unsigned(56,8) ,
67651	 => std_logic_vector(to_unsigned(28,8) ,
67652	 => std_logic_vector(to_unsigned(38,8) ,
67653	 => std_logic_vector(to_unsigned(79,8) ,
67654	 => std_logic_vector(to_unsigned(95,8) ,
67655	 => std_logic_vector(to_unsigned(105,8) ,
67656	 => std_logic_vector(to_unsigned(107,8) ,
67657	 => std_logic_vector(to_unsigned(114,8) ,
67658	 => std_logic_vector(to_unsigned(114,8) ,
67659	 => std_logic_vector(to_unsigned(45,8) ,
67660	 => std_logic_vector(to_unsigned(20,8) ,
67661	 => std_logic_vector(to_unsigned(38,8) ,
67662	 => std_logic_vector(to_unsigned(55,8) ,
67663	 => std_logic_vector(to_unsigned(48,8) ,
67664	 => std_logic_vector(to_unsigned(67,8) ,
67665	 => std_logic_vector(to_unsigned(73,8) ,
67666	 => std_logic_vector(to_unsigned(63,8) ,
67667	 => std_logic_vector(to_unsigned(45,8) ,
67668	 => std_logic_vector(to_unsigned(25,8) ,
67669	 => std_logic_vector(to_unsigned(45,8) ,
67670	 => std_logic_vector(to_unsigned(53,8) ,
67671	 => std_logic_vector(to_unsigned(57,8) ,
67672	 => std_logic_vector(to_unsigned(72,8) ,
67673	 => std_logic_vector(to_unsigned(50,8) ,
67674	 => std_logic_vector(to_unsigned(42,8) ,
67675	 => std_logic_vector(to_unsigned(63,8) ,
67676	 => std_logic_vector(to_unsigned(39,8) ,
67677	 => std_logic_vector(to_unsigned(8,8) ,
67678	 => std_logic_vector(to_unsigned(7,8) ,
67679	 => std_logic_vector(to_unsigned(5,8) ,
67680	 => std_logic_vector(to_unsigned(9,8) ,
67681	 => std_logic_vector(to_unsigned(17,8) ,
67682	 => std_logic_vector(to_unsigned(11,8) ,
67683	 => std_logic_vector(to_unsigned(12,8) ,
67684	 => std_logic_vector(to_unsigned(25,8) ,
67685	 => std_logic_vector(to_unsigned(23,8) ,
67686	 => std_logic_vector(to_unsigned(13,8) ,
67687	 => std_logic_vector(to_unsigned(22,8) ,
67688	 => std_logic_vector(to_unsigned(34,8) ,
67689	 => std_logic_vector(to_unsigned(38,8) ,
67690	 => std_logic_vector(to_unsigned(25,8) ,
67691	 => std_logic_vector(to_unsigned(21,8) ,
67692	 => std_logic_vector(to_unsigned(27,8) ,
67693	 => std_logic_vector(to_unsigned(19,8) ,
67694	 => std_logic_vector(to_unsigned(26,8) ,
67695	 => std_logic_vector(to_unsigned(30,8) ,
67696	 => std_logic_vector(to_unsigned(20,8) ,
67697	 => std_logic_vector(to_unsigned(51,8) ,
67698	 => std_logic_vector(to_unsigned(74,8) ,
67699	 => std_logic_vector(to_unsigned(35,8) ,
67700	 => std_logic_vector(to_unsigned(29,8) ,
67701	 => std_logic_vector(to_unsigned(21,8) ,
67702	 => std_logic_vector(to_unsigned(14,8) ,
67703	 => std_logic_vector(to_unsigned(13,8) ,
67704	 => std_logic_vector(to_unsigned(12,8) ,
67705	 => std_logic_vector(to_unsigned(12,8) ,
67706	 => std_logic_vector(to_unsigned(30,8) ,
67707	 => std_logic_vector(to_unsigned(51,8) ,
67708	 => std_logic_vector(to_unsigned(54,8) ,
67709	 => std_logic_vector(to_unsigned(42,8) ,
67710	 => std_logic_vector(to_unsigned(40,8) ,
67711	 => std_logic_vector(to_unsigned(48,8) ,
67712	 => std_logic_vector(to_unsigned(29,8) ,
67713	 => std_logic_vector(to_unsigned(13,8) ,
67714	 => std_logic_vector(to_unsigned(17,8) ,
67715	 => std_logic_vector(to_unsigned(43,8) ,
67716	 => std_logic_vector(to_unsigned(40,8) ,
67717	 => std_logic_vector(to_unsigned(49,8) ,
67718	 => std_logic_vector(to_unsigned(61,8) ,
67719	 => std_logic_vector(to_unsigned(50,8) ,
67720	 => std_logic_vector(to_unsigned(47,8) ,
67721	 => std_logic_vector(to_unsigned(31,8) ,
67722	 => std_logic_vector(to_unsigned(22,8) ,
67723	 => std_logic_vector(to_unsigned(18,8) ,
67724	 => std_logic_vector(to_unsigned(14,8) ,
67725	 => std_logic_vector(to_unsigned(17,8) ,
67726	 => std_logic_vector(to_unsigned(13,8) ,
67727	 => std_logic_vector(to_unsigned(12,8) ,
67728	 => std_logic_vector(to_unsigned(27,8) ,
67729	 => std_logic_vector(to_unsigned(41,8) ,
67730	 => std_logic_vector(to_unsigned(45,8) ,
67731	 => std_logic_vector(to_unsigned(34,8) ,
67732	 => std_logic_vector(to_unsigned(25,8) ,
67733	 => std_logic_vector(to_unsigned(34,8) ,
67734	 => std_logic_vector(to_unsigned(25,8) ,
67735	 => std_logic_vector(to_unsigned(12,8) ,
67736	 => std_logic_vector(to_unsigned(15,8) ,
67737	 => std_logic_vector(to_unsigned(25,8) ,
67738	 => std_logic_vector(to_unsigned(33,8) ,
67739	 => std_logic_vector(to_unsigned(25,8) ,
67740	 => std_logic_vector(to_unsigned(22,8) ,
67741	 => std_logic_vector(to_unsigned(27,8) ,
67742	 => std_logic_vector(to_unsigned(20,8) ,
67743	 => std_logic_vector(to_unsigned(29,8) ,
67744	 => std_logic_vector(to_unsigned(38,8) ,
67745	 => std_logic_vector(to_unsigned(31,8) ,
67746	 => std_logic_vector(to_unsigned(39,8) ,
67747	 => std_logic_vector(to_unsigned(30,8) ,
67748	 => std_logic_vector(to_unsigned(19,8) ,
67749	 => std_logic_vector(to_unsigned(5,8) ,
67750	 => std_logic_vector(to_unsigned(15,8) ,
67751	 => std_logic_vector(to_unsigned(45,8) ,
67752	 => std_logic_vector(to_unsigned(17,8) ,
67753	 => std_logic_vector(to_unsigned(28,8) ,
67754	 => std_logic_vector(to_unsigned(47,8) ,
67755	 => std_logic_vector(to_unsigned(54,8) ,
67756	 => std_logic_vector(to_unsigned(59,8) ,
67757	 => std_logic_vector(to_unsigned(69,8) ,
67758	 => std_logic_vector(to_unsigned(55,8) ,
67759	 => std_logic_vector(to_unsigned(50,8) ,
67760	 => std_logic_vector(to_unsigned(55,8) ,
67761	 => std_logic_vector(to_unsigned(57,8) ,
67762	 => std_logic_vector(to_unsigned(51,8) ,
67763	 => std_logic_vector(to_unsigned(51,8) ,
67764	 => std_logic_vector(to_unsigned(86,8) ,
67765	 => std_logic_vector(to_unsigned(111,8) ,
67766	 => std_logic_vector(to_unsigned(53,8) ,
67767	 => std_logic_vector(to_unsigned(56,8) ,
67768	 => std_logic_vector(to_unsigned(119,8) ,
67769	 => std_logic_vector(to_unsigned(127,8) ,
67770	 => std_logic_vector(to_unsigned(60,8) ,
67771	 => std_logic_vector(to_unsigned(13,8) ,
67772	 => std_logic_vector(to_unsigned(16,8) ,
67773	 => std_logic_vector(to_unsigned(10,8) ,
67774	 => std_logic_vector(to_unsigned(7,8) ,
67775	 => std_logic_vector(to_unsigned(12,8) ,
67776	 => std_logic_vector(to_unsigned(13,8) ,
67777	 => std_logic_vector(to_unsigned(24,8) ,
67778	 => std_logic_vector(to_unsigned(49,8) ,
67779	 => std_logic_vector(to_unsigned(19,8) ,
67780	 => std_logic_vector(to_unsigned(11,8) ,
67781	 => std_logic_vector(to_unsigned(9,8) ,
67782	 => std_logic_vector(to_unsigned(11,8) ,
67783	 => std_logic_vector(to_unsigned(14,8) ,
67784	 => std_logic_vector(to_unsigned(14,8) ,
67785	 => std_logic_vector(to_unsigned(30,8) ,
67786	 => std_logic_vector(to_unsigned(39,8) ,
67787	 => std_logic_vector(to_unsigned(16,8) ,
67788	 => std_logic_vector(to_unsigned(20,8) ,
67789	 => std_logic_vector(to_unsigned(14,8) ,
67790	 => std_logic_vector(to_unsigned(29,8) ,
67791	 => std_logic_vector(to_unsigned(37,8) ,
67792	 => std_logic_vector(to_unsigned(11,8) ,
67793	 => std_logic_vector(to_unsigned(4,8) ,
67794	 => std_logic_vector(to_unsigned(0,8) ,
67795	 => std_logic_vector(to_unsigned(1,8) ,
67796	 => std_logic_vector(to_unsigned(8,8) ,
67797	 => std_logic_vector(to_unsigned(8,8) ,
67798	 => std_logic_vector(to_unsigned(7,8) ,
67799	 => std_logic_vector(to_unsigned(10,8) ,
67800	 => std_logic_vector(to_unsigned(5,8) ,
67801	 => std_logic_vector(to_unsigned(4,8) ,
67802	 => std_logic_vector(to_unsigned(5,8) ,
67803	 => std_logic_vector(to_unsigned(6,8) ,
67804	 => std_logic_vector(to_unsigned(8,8) ,
67805	 => std_logic_vector(to_unsigned(2,8) ,
67806	 => std_logic_vector(to_unsigned(0,8) ,
67807	 => std_logic_vector(to_unsigned(4,8) ,
67808	 => std_logic_vector(to_unsigned(10,8) ,
67809	 => std_logic_vector(to_unsigned(10,8) ,
67810	 => std_logic_vector(to_unsigned(35,8) ,
67811	 => std_logic_vector(to_unsigned(57,8) ,
67812	 => std_logic_vector(to_unsigned(45,8) ,
67813	 => std_logic_vector(to_unsigned(37,8) ,
67814	 => std_logic_vector(to_unsigned(31,8) ,
67815	 => std_logic_vector(to_unsigned(30,8) ,
67816	 => std_logic_vector(to_unsigned(39,8) ,
67817	 => std_logic_vector(to_unsigned(39,8) ,
67818	 => std_logic_vector(to_unsigned(27,8) ,
67819	 => std_logic_vector(to_unsigned(2,8) ,
67820	 => std_logic_vector(to_unsigned(0,8) ,
67821	 => std_logic_vector(to_unsigned(14,8) ,
67822	 => std_logic_vector(to_unsigned(119,8) ,
67823	 => std_logic_vector(to_unsigned(100,8) ,
67824	 => std_logic_vector(to_unsigned(96,8) ,
67825	 => std_logic_vector(to_unsigned(104,8) ,
67826	 => std_logic_vector(to_unsigned(55,8) ,
67827	 => std_logic_vector(to_unsigned(30,8) ,
67828	 => std_logic_vector(to_unsigned(34,8) ,
67829	 => std_logic_vector(to_unsigned(46,8) ,
67830	 => std_logic_vector(to_unsigned(52,8) ,
67831	 => std_logic_vector(to_unsigned(51,8) ,
67832	 => std_logic_vector(to_unsigned(50,8) ,
67833	 => std_logic_vector(to_unsigned(49,8) ,
67834	 => std_logic_vector(to_unsigned(32,8) ,
67835	 => std_logic_vector(to_unsigned(20,8) ,
67836	 => std_logic_vector(to_unsigned(68,8) ,
67837	 => std_logic_vector(to_unsigned(92,8) ,
67838	 => std_logic_vector(to_unsigned(93,8) ,
67839	 => std_logic_vector(to_unsigned(99,8) ,
67840	 => std_logic_vector(to_unsigned(92,8) ,
67841	 => std_logic_vector(to_unsigned(115,8) ,
67842	 => std_logic_vector(to_unsigned(116,8) ,
67843	 => std_logic_vector(to_unsigned(109,8) ,
67844	 => std_logic_vector(to_unsigned(103,8) ,
67845	 => std_logic_vector(to_unsigned(84,8) ,
67846	 => std_logic_vector(to_unsigned(109,8) ,
67847	 => std_logic_vector(to_unsigned(104,8) ,
67848	 => std_logic_vector(to_unsigned(93,8) ,
67849	 => std_logic_vector(to_unsigned(82,8) ,
67850	 => std_logic_vector(to_unsigned(87,8) ,
67851	 => std_logic_vector(to_unsigned(69,8) ,
67852	 => std_logic_vector(to_unsigned(45,8) ,
67853	 => std_logic_vector(to_unsigned(38,8) ,
67854	 => std_logic_vector(to_unsigned(37,8) ,
67855	 => std_logic_vector(to_unsigned(27,8) ,
67856	 => std_logic_vector(to_unsigned(46,8) ,
67857	 => std_logic_vector(to_unsigned(81,8) ,
67858	 => std_logic_vector(to_unsigned(58,8) ,
67859	 => std_logic_vector(to_unsigned(51,8) ,
67860	 => std_logic_vector(to_unsigned(40,8) ,
67861	 => std_logic_vector(to_unsigned(38,8) ,
67862	 => std_logic_vector(to_unsigned(53,8) ,
67863	 => std_logic_vector(to_unsigned(46,8) ,
67864	 => std_logic_vector(to_unsigned(36,8) ,
67865	 => std_logic_vector(to_unsigned(41,8) ,
67866	 => std_logic_vector(to_unsigned(41,8) ,
67867	 => std_logic_vector(to_unsigned(34,8) ,
67868	 => std_logic_vector(to_unsigned(34,8) ,
67869	 => std_logic_vector(to_unsigned(32,8) ,
67870	 => std_logic_vector(to_unsigned(34,8) ,
67871	 => std_logic_vector(to_unsigned(37,8) ,
67872	 => std_logic_vector(to_unsigned(37,8) ,
67873	 => std_logic_vector(to_unsigned(31,8) ,
67874	 => std_logic_vector(to_unsigned(30,8) ,
67875	 => std_logic_vector(to_unsigned(34,8) ,
67876	 => std_logic_vector(to_unsigned(32,8) ,
67877	 => std_logic_vector(to_unsigned(29,8) ,
67878	 => std_logic_vector(to_unsigned(30,8) ,
67879	 => std_logic_vector(to_unsigned(29,8) ,
67880	 => std_logic_vector(to_unsigned(35,8) ,
67881	 => std_logic_vector(to_unsigned(58,8) ,
67882	 => std_logic_vector(to_unsigned(59,8) ,
67883	 => std_logic_vector(to_unsigned(46,8) ,
67884	 => std_logic_vector(to_unsigned(74,8) ,
67885	 => std_logic_vector(to_unsigned(64,8) ,
67886	 => std_logic_vector(to_unsigned(54,8) ,
67887	 => std_logic_vector(to_unsigned(56,8) ,
67888	 => std_logic_vector(to_unsigned(39,8) ,
67889	 => std_logic_vector(to_unsigned(27,8) ,
67890	 => std_logic_vector(to_unsigned(37,8) ,
67891	 => std_logic_vector(to_unsigned(45,8) ,
67892	 => std_logic_vector(to_unsigned(49,8) ,
67893	 => std_logic_vector(to_unsigned(43,8) ,
67894	 => std_logic_vector(to_unsigned(32,8) ,
67895	 => std_logic_vector(to_unsigned(56,8) ,
67896	 => std_logic_vector(to_unsigned(81,8) ,
67897	 => std_logic_vector(to_unsigned(76,8) ,
67898	 => std_logic_vector(to_unsigned(47,8) ,
67899	 => std_logic_vector(to_unsigned(41,8) ,
67900	 => std_logic_vector(to_unsigned(38,8) ,
67901	 => std_logic_vector(to_unsigned(43,8) ,
67902	 => std_logic_vector(to_unsigned(46,8) ,
67903	 => std_logic_vector(to_unsigned(35,8) ,
67904	 => std_logic_vector(to_unsigned(29,8) ,
67905	 => std_logic_vector(to_unsigned(38,8) ,
67906	 => std_logic_vector(to_unsigned(71,8) ,
67907	 => std_logic_vector(to_unsigned(80,8) ,
67908	 => std_logic_vector(to_unsigned(85,8) ,
67909	 => std_logic_vector(to_unsigned(96,8) ,
67910	 => std_logic_vector(to_unsigned(107,8) ,
67911	 => std_logic_vector(to_unsigned(109,8) ,
67912	 => std_logic_vector(to_unsigned(95,8) ,
67913	 => std_logic_vector(to_unsigned(90,8) ,
67914	 => std_logic_vector(to_unsigned(88,8) ,
67915	 => std_logic_vector(to_unsigned(87,8) ,
67916	 => std_logic_vector(to_unsigned(93,8) ,
67917	 => std_logic_vector(to_unsigned(82,8) ,
67918	 => std_logic_vector(to_unsigned(81,8) ,
67919	 => std_logic_vector(to_unsigned(92,8) ,
67920	 => std_logic_vector(to_unsigned(91,8) ,
67921	 => std_logic_vector(to_unsigned(86,8) ,
67922	 => std_logic_vector(to_unsigned(76,8) ,
67923	 => std_logic_vector(to_unsigned(77,8) ,
67924	 => std_logic_vector(to_unsigned(92,8) ,
67925	 => std_logic_vector(to_unsigned(105,8) ,
67926	 => std_logic_vector(to_unsigned(88,8) ,
67927	 => std_logic_vector(to_unsigned(80,8) ,
67928	 => std_logic_vector(to_unsigned(80,8) ,
67929	 => std_logic_vector(to_unsigned(62,8) ,
67930	 => std_logic_vector(to_unsigned(22,8) ,
67931	 => std_logic_vector(to_unsigned(19,8) ,
67932	 => std_logic_vector(to_unsigned(45,8) ,
67933	 => std_logic_vector(to_unsigned(42,8) ,
67934	 => std_logic_vector(to_unsigned(39,8) ,
67935	 => std_logic_vector(to_unsigned(49,8) ,
67936	 => std_logic_vector(to_unsigned(33,8) ,
67937	 => std_logic_vector(to_unsigned(42,8) ,
67938	 => std_logic_vector(to_unsigned(54,8) ,
67939	 => std_logic_vector(to_unsigned(44,8) ,
67940	 => std_logic_vector(to_unsigned(51,8) ,
67941	 => std_logic_vector(to_unsigned(51,8) ,
67942	 => std_logic_vector(to_unsigned(39,8) ,
67943	 => std_logic_vector(to_unsigned(27,8) ,
67944	 => std_logic_vector(to_unsigned(21,8) ,
67945	 => std_logic_vector(to_unsigned(21,8) ,
67946	 => std_logic_vector(to_unsigned(17,8) ,
67947	 => std_logic_vector(to_unsigned(12,8) ,
67948	 => std_logic_vector(to_unsigned(9,8) ,
67949	 => std_logic_vector(to_unsigned(26,8) ,
67950	 => std_logic_vector(to_unsigned(67,8) ,
67951	 => std_logic_vector(to_unsigned(60,8) ,
67952	 => std_logic_vector(to_unsigned(41,8) ,
67953	 => std_logic_vector(to_unsigned(45,8) ,
67954	 => std_logic_vector(to_unsigned(41,8) ,
67955	 => std_logic_vector(to_unsigned(45,8) ,
67956	 => std_logic_vector(to_unsigned(116,8) ,
67957	 => std_logic_vector(to_unsigned(147,8) ,
67958	 => std_logic_vector(to_unsigned(79,8) ,
67959	 => std_logic_vector(to_unsigned(21,8) ,
67960	 => std_logic_vector(to_unsigned(34,8) ,
67961	 => std_logic_vector(to_unsigned(56,8) ,
67962	 => std_logic_vector(to_unsigned(51,8) ,
67963	 => std_logic_vector(to_unsigned(45,8) ,
67964	 => std_logic_vector(to_unsigned(45,8) ,
67965	 => std_logic_vector(to_unsigned(51,8) ,
67966	 => std_logic_vector(to_unsigned(51,8) ,
67967	 => std_logic_vector(to_unsigned(49,8) ,
67968	 => std_logic_vector(to_unsigned(51,8) ,
67969	 => std_logic_vector(to_unsigned(50,8) ,
67970	 => std_logic_vector(to_unsigned(27,8) ,
67971	 => std_logic_vector(to_unsigned(36,8) ,
67972	 => std_logic_vector(to_unsigned(80,8) ,
67973	 => std_logic_vector(to_unsigned(100,8) ,
67974	 => std_logic_vector(to_unsigned(116,8) ,
67975	 => std_logic_vector(to_unsigned(116,8) ,
67976	 => std_logic_vector(to_unsigned(107,8) ,
67977	 => std_logic_vector(to_unsigned(107,8) ,
67978	 => std_logic_vector(to_unsigned(107,8) ,
67979	 => std_logic_vector(to_unsigned(57,8) ,
67980	 => std_logic_vector(to_unsigned(23,8) ,
67981	 => std_logic_vector(to_unsigned(36,8) ,
67982	 => std_logic_vector(to_unsigned(46,8) ,
67983	 => std_logic_vector(to_unsigned(51,8) ,
67984	 => std_logic_vector(to_unsigned(48,8) ,
67985	 => std_logic_vector(to_unsigned(50,8) ,
67986	 => std_logic_vector(to_unsigned(67,8) ,
67987	 => std_logic_vector(to_unsigned(48,8) ,
67988	 => std_logic_vector(to_unsigned(17,8) ,
67989	 => std_logic_vector(to_unsigned(40,8) ,
67990	 => std_logic_vector(to_unsigned(64,8) ,
67991	 => std_logic_vector(to_unsigned(82,8) ,
67992	 => std_logic_vector(to_unsigned(65,8) ,
67993	 => std_logic_vector(to_unsigned(60,8) ,
67994	 => std_logic_vector(to_unsigned(56,8) ,
67995	 => std_logic_vector(to_unsigned(61,8) ,
67996	 => std_logic_vector(to_unsigned(37,8) ,
67997	 => std_logic_vector(to_unsigned(8,8) ,
67998	 => std_logic_vector(to_unsigned(7,8) ,
67999	 => std_logic_vector(to_unsigned(6,8) ,
68000	 => std_logic_vector(to_unsigned(13,8) ,
68001	 => std_logic_vector(to_unsigned(29,8) ,
68002	 => std_logic_vector(to_unsigned(18,8) ,
68003	 => std_logic_vector(to_unsigned(16,8) ,
68004	 => std_logic_vector(to_unsigned(29,8) ,
68005	 => std_logic_vector(to_unsigned(19,8) ,
68006	 => std_logic_vector(to_unsigned(9,8) ,
68007	 => std_logic_vector(to_unsigned(11,8) ,
68008	 => std_logic_vector(to_unsigned(15,8) ,
68009	 => std_logic_vector(to_unsigned(35,8) ,
68010	 => std_logic_vector(to_unsigned(27,8) ,
68011	 => std_logic_vector(to_unsigned(27,8) ,
68012	 => std_logic_vector(to_unsigned(24,8) ,
68013	 => std_logic_vector(to_unsigned(24,8) ,
68014	 => std_logic_vector(to_unsigned(36,8) ,
68015	 => std_logic_vector(to_unsigned(25,8) ,
68016	 => std_logic_vector(to_unsigned(38,8) ,
68017	 => std_logic_vector(to_unsigned(65,8) ,
68018	 => std_logic_vector(to_unsigned(35,8) ,
68019	 => std_logic_vector(to_unsigned(29,8) ,
68020	 => std_logic_vector(to_unsigned(31,8) ,
68021	 => std_logic_vector(to_unsigned(12,8) ,
68022	 => std_logic_vector(to_unsigned(13,8) ,
68023	 => std_logic_vector(to_unsigned(17,8) ,
68024	 => std_logic_vector(to_unsigned(15,8) ,
68025	 => std_logic_vector(to_unsigned(20,8) ,
68026	 => std_logic_vector(to_unsigned(35,8) ,
68027	 => std_logic_vector(to_unsigned(37,8) ,
68028	 => std_logic_vector(to_unsigned(42,8) ,
68029	 => std_logic_vector(to_unsigned(43,8) ,
68030	 => std_logic_vector(to_unsigned(35,8) ,
68031	 => std_logic_vector(to_unsigned(37,8) ,
68032	 => std_logic_vector(to_unsigned(47,8) ,
68033	 => std_logic_vector(to_unsigned(53,8) ,
68034	 => std_logic_vector(to_unsigned(43,8) ,
68035	 => std_logic_vector(to_unsigned(38,8) ,
68036	 => std_logic_vector(to_unsigned(36,8) ,
68037	 => std_logic_vector(to_unsigned(59,8) ,
68038	 => std_logic_vector(to_unsigned(93,8) ,
68039	 => std_logic_vector(to_unsigned(77,8) ,
68040	 => std_logic_vector(to_unsigned(41,8) ,
68041	 => std_logic_vector(to_unsigned(36,8) ,
68042	 => std_logic_vector(to_unsigned(22,8) ,
68043	 => std_logic_vector(to_unsigned(8,8) ,
68044	 => std_logic_vector(to_unsigned(18,8) ,
68045	 => std_logic_vector(to_unsigned(22,8) ,
68046	 => std_logic_vector(to_unsigned(13,8) ,
68047	 => std_logic_vector(to_unsigned(9,8) ,
68048	 => std_logic_vector(to_unsigned(23,8) ,
68049	 => std_logic_vector(to_unsigned(41,8) ,
68050	 => std_logic_vector(to_unsigned(65,8) ,
68051	 => std_logic_vector(to_unsigned(52,8) ,
68052	 => std_logic_vector(to_unsigned(30,8) ,
68053	 => std_logic_vector(to_unsigned(33,8) ,
68054	 => std_logic_vector(to_unsigned(35,8) ,
68055	 => std_logic_vector(to_unsigned(19,8) ,
68056	 => std_logic_vector(to_unsigned(15,8) ,
68057	 => std_logic_vector(to_unsigned(23,8) ,
68058	 => std_logic_vector(to_unsigned(31,8) ,
68059	 => std_logic_vector(to_unsigned(28,8) ,
68060	 => std_logic_vector(to_unsigned(16,8) ,
68061	 => std_logic_vector(to_unsigned(9,8) ,
68062	 => std_logic_vector(to_unsigned(16,8) ,
68063	 => std_logic_vector(to_unsigned(31,8) ,
68064	 => std_logic_vector(to_unsigned(44,8) ,
68065	 => std_logic_vector(to_unsigned(37,8) ,
68066	 => std_logic_vector(to_unsigned(35,8) ,
68067	 => std_logic_vector(to_unsigned(38,8) ,
68068	 => std_logic_vector(to_unsigned(27,8) ,
68069	 => std_logic_vector(to_unsigned(5,8) ,
68070	 => std_logic_vector(to_unsigned(13,8) ,
68071	 => std_logic_vector(to_unsigned(35,8) ,
68072	 => std_logic_vector(to_unsigned(5,8) ,
68073	 => std_logic_vector(to_unsigned(17,8) ,
68074	 => std_logic_vector(to_unsigned(50,8) ,
68075	 => std_logic_vector(to_unsigned(68,8) ,
68076	 => std_logic_vector(to_unsigned(35,8) ,
68077	 => std_logic_vector(to_unsigned(29,8) ,
68078	 => std_logic_vector(to_unsigned(67,8) ,
68079	 => std_logic_vector(to_unsigned(67,8) ,
68080	 => std_logic_vector(to_unsigned(51,8) ,
68081	 => std_logic_vector(to_unsigned(31,8) ,
68082	 => std_logic_vector(to_unsigned(41,8) ,
68083	 => std_logic_vector(to_unsigned(66,8) ,
68084	 => std_logic_vector(to_unsigned(90,8) ,
68085	 => std_logic_vector(to_unsigned(114,8) ,
68086	 => std_logic_vector(to_unsigned(52,8) ,
68087	 => std_logic_vector(to_unsigned(53,8) ,
68088	 => std_logic_vector(to_unsigned(116,8) ,
68089	 => std_logic_vector(to_unsigned(122,8) ,
68090	 => std_logic_vector(to_unsigned(78,8) ,
68091	 => std_logic_vector(to_unsigned(32,8) ,
68092	 => std_logic_vector(to_unsigned(30,8) ,
68093	 => std_logic_vector(to_unsigned(25,8) ,
68094	 => std_logic_vector(to_unsigned(15,8) ,
68095	 => std_logic_vector(to_unsigned(14,8) ,
68096	 => std_logic_vector(to_unsigned(13,8) ,
68097	 => std_logic_vector(to_unsigned(30,8) ,
68098	 => std_logic_vector(to_unsigned(41,8) ,
68099	 => std_logic_vector(to_unsigned(12,8) ,
68100	 => std_logic_vector(to_unsigned(12,8) ,
68101	 => std_logic_vector(to_unsigned(10,8) ,
68102	 => std_logic_vector(to_unsigned(8,8) ,
68103	 => std_logic_vector(to_unsigned(6,8) ,
68104	 => std_logic_vector(to_unsigned(9,8) ,
68105	 => std_logic_vector(to_unsigned(21,8) ,
68106	 => std_logic_vector(to_unsigned(30,8) ,
68107	 => std_logic_vector(to_unsigned(26,8) ,
68108	 => std_logic_vector(to_unsigned(15,8) ,
68109	 => std_logic_vector(to_unsigned(11,8) ,
68110	 => std_logic_vector(to_unsigned(32,8) ,
68111	 => std_logic_vector(to_unsigned(48,8) ,
68112	 => std_logic_vector(to_unsigned(22,8) ,
68113	 => std_logic_vector(to_unsigned(8,8) ,
68114	 => std_logic_vector(to_unsigned(0,8) ,
68115	 => std_logic_vector(to_unsigned(1,8) ,
68116	 => std_logic_vector(to_unsigned(6,8) ,
68117	 => std_logic_vector(to_unsigned(6,8) ,
68118	 => std_logic_vector(to_unsigned(7,8) ,
68119	 => std_logic_vector(to_unsigned(11,8) ,
68120	 => std_logic_vector(to_unsigned(8,8) ,
68121	 => std_logic_vector(to_unsigned(8,8) ,
68122	 => std_logic_vector(to_unsigned(6,8) ,
68123	 => std_logic_vector(to_unsigned(8,8) ,
68124	 => std_logic_vector(to_unsigned(8,8) ,
68125	 => std_logic_vector(to_unsigned(1,8) ,
68126	 => std_logic_vector(to_unsigned(0,8) ,
68127	 => std_logic_vector(to_unsigned(2,8) ,
68128	 => std_logic_vector(to_unsigned(6,8) ,
68129	 => std_logic_vector(to_unsigned(9,8) ,
68130	 => std_logic_vector(to_unsigned(25,8) ,
68131	 => std_logic_vector(to_unsigned(43,8) ,
68132	 => std_logic_vector(to_unsigned(67,8) ,
68133	 => std_logic_vector(to_unsigned(58,8) ,
68134	 => std_logic_vector(to_unsigned(54,8) ,
68135	 => std_logic_vector(to_unsigned(45,8) ,
68136	 => std_logic_vector(to_unsigned(35,8) ,
68137	 => std_logic_vector(to_unsigned(36,8) ,
68138	 => std_logic_vector(to_unsigned(33,8) ,
68139	 => std_logic_vector(to_unsigned(8,8) ,
68140	 => std_logic_vector(to_unsigned(0,8) ,
68141	 => std_logic_vector(to_unsigned(1,8) ,
68142	 => std_logic_vector(to_unsigned(25,8) ,
68143	 => std_logic_vector(to_unsigned(69,8) ,
68144	 => std_logic_vector(to_unsigned(78,8) ,
68145	 => std_logic_vector(to_unsigned(105,8) ,
68146	 => std_logic_vector(to_unsigned(45,8) ,
68147	 => std_logic_vector(to_unsigned(22,8) ,
68148	 => std_logic_vector(to_unsigned(24,8) ,
68149	 => std_logic_vector(to_unsigned(17,8) ,
68150	 => std_logic_vector(to_unsigned(22,8) ,
68151	 => std_logic_vector(to_unsigned(23,8) ,
68152	 => std_logic_vector(to_unsigned(25,8) ,
68153	 => std_logic_vector(to_unsigned(33,8) ,
68154	 => std_logic_vector(to_unsigned(35,8) ,
68155	 => std_logic_vector(to_unsigned(49,8) ,
68156	 => std_logic_vector(to_unsigned(116,8) ,
68157	 => std_logic_vector(to_unsigned(114,8) ,
68158	 => std_logic_vector(to_unsigned(109,8) ,
68159	 => std_logic_vector(to_unsigned(105,8) ,
68160	 => std_logic_vector(to_unsigned(103,8) ,
68161	 => std_logic_vector(to_unsigned(112,8) ,
68162	 => std_logic_vector(to_unsigned(118,8) ,
68163	 => std_logic_vector(to_unsigned(115,8) ,
68164	 => std_logic_vector(to_unsigned(108,8) ,
68165	 => std_logic_vector(to_unsigned(104,8) ,
68166	 => std_logic_vector(to_unsigned(107,8) ,
68167	 => std_logic_vector(to_unsigned(105,8) ,
68168	 => std_logic_vector(to_unsigned(107,8) ,
68169	 => std_logic_vector(to_unsigned(101,8) ,
68170	 => std_logic_vector(to_unsigned(107,8) ,
68171	 => std_logic_vector(to_unsigned(77,8) ,
68172	 => std_logic_vector(to_unsigned(46,8) ,
68173	 => std_logic_vector(to_unsigned(42,8) ,
68174	 => std_logic_vector(to_unsigned(31,8) ,
68175	 => std_logic_vector(to_unsigned(29,8) ,
68176	 => std_logic_vector(to_unsigned(42,8) ,
68177	 => std_logic_vector(to_unsigned(67,8) ,
68178	 => std_logic_vector(to_unsigned(67,8) ,
68179	 => std_logic_vector(to_unsigned(64,8) ,
68180	 => std_logic_vector(to_unsigned(54,8) ,
68181	 => std_logic_vector(to_unsigned(41,8) ,
68182	 => std_logic_vector(to_unsigned(42,8) ,
68183	 => std_logic_vector(to_unsigned(48,8) ,
68184	 => std_logic_vector(to_unsigned(42,8) ,
68185	 => std_logic_vector(to_unsigned(40,8) ,
68186	 => std_logic_vector(to_unsigned(37,8) ,
68187	 => std_logic_vector(to_unsigned(35,8) ,
68188	 => std_logic_vector(to_unsigned(37,8) ,
68189	 => std_logic_vector(to_unsigned(31,8) ,
68190	 => std_logic_vector(to_unsigned(34,8) ,
68191	 => std_logic_vector(to_unsigned(29,8) ,
68192	 => std_logic_vector(to_unsigned(29,8) ,
68193	 => std_logic_vector(to_unsigned(25,8) ,
68194	 => std_logic_vector(to_unsigned(30,8) ,
68195	 => std_logic_vector(to_unsigned(33,8) ,
68196	 => std_logic_vector(to_unsigned(29,8) ,
68197	 => std_logic_vector(to_unsigned(26,8) ,
68198	 => std_logic_vector(to_unsigned(25,8) ,
68199	 => std_logic_vector(to_unsigned(42,8) ,
68200	 => std_logic_vector(to_unsigned(64,8) ,
68201	 => std_logic_vector(to_unsigned(74,8) ,
68202	 => std_logic_vector(to_unsigned(58,8) ,
68203	 => std_logic_vector(to_unsigned(65,8) ,
68204	 => std_logic_vector(to_unsigned(72,8) ,
68205	 => std_logic_vector(to_unsigned(52,8) ,
68206	 => std_logic_vector(to_unsigned(38,8) ,
68207	 => std_logic_vector(to_unsigned(34,8) ,
68208	 => std_logic_vector(to_unsigned(38,8) ,
68209	 => std_logic_vector(to_unsigned(30,8) ,
68210	 => std_logic_vector(to_unsigned(30,8) ,
68211	 => std_logic_vector(to_unsigned(44,8) ,
68212	 => std_logic_vector(to_unsigned(53,8) ,
68213	 => std_logic_vector(to_unsigned(62,8) ,
68214	 => std_logic_vector(to_unsigned(67,8) ,
68215	 => std_logic_vector(to_unsigned(77,8) ,
68216	 => std_logic_vector(to_unsigned(79,8) ,
68217	 => std_logic_vector(to_unsigned(95,8) ,
68218	 => std_logic_vector(to_unsigned(57,8) ,
68219	 => std_logic_vector(to_unsigned(30,8) ,
68220	 => std_logic_vector(to_unsigned(37,8) ,
68221	 => std_logic_vector(to_unsigned(35,8) ,
68222	 => std_logic_vector(to_unsigned(35,8) ,
68223	 => std_logic_vector(to_unsigned(31,8) ,
68224	 => std_logic_vector(to_unsigned(33,8) ,
68225	 => std_logic_vector(to_unsigned(36,8) ,
68226	 => std_logic_vector(to_unsigned(61,8) ,
68227	 => std_logic_vector(to_unsigned(85,8) ,
68228	 => std_logic_vector(to_unsigned(96,8) ,
68229	 => std_logic_vector(to_unsigned(101,8) ,
68230	 => std_logic_vector(to_unsigned(101,8) ,
68231	 => std_logic_vector(to_unsigned(100,8) ,
68232	 => std_logic_vector(to_unsigned(91,8) ,
68233	 => std_logic_vector(to_unsigned(87,8) ,
68234	 => std_logic_vector(to_unsigned(81,8) ,
68235	 => std_logic_vector(to_unsigned(80,8) ,
68236	 => std_logic_vector(to_unsigned(84,8) ,
68237	 => std_logic_vector(to_unsigned(84,8) ,
68238	 => std_logic_vector(to_unsigned(91,8) ,
68239	 => std_logic_vector(to_unsigned(80,8) ,
68240	 => std_logic_vector(to_unsigned(87,8) ,
68241	 => std_logic_vector(to_unsigned(80,8) ,
68242	 => std_logic_vector(to_unsigned(76,8) ,
68243	 => std_logic_vector(to_unsigned(90,8) ,
68244	 => std_logic_vector(to_unsigned(95,8) ,
68245	 => std_logic_vector(to_unsigned(84,8) ,
68246	 => std_logic_vector(to_unsigned(71,8) ,
68247	 => std_logic_vector(to_unsigned(74,8) ,
68248	 => std_logic_vector(to_unsigned(72,8) ,
68249	 => std_logic_vector(to_unsigned(37,8) ,
68250	 => std_logic_vector(to_unsigned(18,8) ,
68251	 => std_logic_vector(to_unsigned(22,8) ,
68252	 => std_logic_vector(to_unsigned(38,8) ,
68253	 => std_logic_vector(to_unsigned(43,8) ,
68254	 => std_logic_vector(to_unsigned(45,8) ,
68255	 => std_logic_vector(to_unsigned(46,8) ,
68256	 => std_logic_vector(to_unsigned(46,8) ,
68257	 => std_logic_vector(to_unsigned(45,8) ,
68258	 => std_logic_vector(to_unsigned(60,8) ,
68259	 => std_logic_vector(to_unsigned(52,8) ,
68260	 => std_logic_vector(to_unsigned(73,8) ,
68261	 => std_logic_vector(to_unsigned(56,8) ,
68262	 => std_logic_vector(to_unsigned(32,8) ,
68263	 => std_logic_vector(to_unsigned(27,8) ,
68264	 => std_logic_vector(to_unsigned(18,8) ,
68265	 => std_logic_vector(to_unsigned(22,8) ,
68266	 => std_logic_vector(to_unsigned(19,8) ,
68267	 => std_logic_vector(to_unsigned(10,8) ,
68268	 => std_logic_vector(to_unsigned(10,8) ,
68269	 => std_logic_vector(to_unsigned(32,8) ,
68270	 => std_logic_vector(to_unsigned(91,8) ,
68271	 => std_logic_vector(to_unsigned(61,8) ,
68272	 => std_logic_vector(to_unsigned(32,8) ,
68273	 => std_logic_vector(to_unsigned(107,8) ,
68274	 => std_logic_vector(to_unsigned(139,8) ,
68275	 => std_logic_vector(to_unsigned(57,8) ,
68276	 => std_logic_vector(to_unsigned(90,8) ,
68277	 => std_logic_vector(to_unsigned(118,8) ,
68278	 => std_logic_vector(to_unsigned(76,8) ,
68279	 => std_logic_vector(to_unsigned(61,8) ,
68280	 => std_logic_vector(to_unsigned(70,8) ,
68281	 => std_logic_vector(to_unsigned(85,8) ,
68282	 => std_logic_vector(to_unsigned(49,8) ,
68283	 => std_logic_vector(to_unsigned(20,8) ,
68284	 => std_logic_vector(to_unsigned(25,8) ,
68285	 => std_logic_vector(to_unsigned(27,8) ,
68286	 => std_logic_vector(to_unsigned(32,8) ,
68287	 => std_logic_vector(to_unsigned(35,8) ,
68288	 => std_logic_vector(to_unsigned(37,8) ,
68289	 => std_logic_vector(to_unsigned(29,8) ,
68290	 => std_logic_vector(to_unsigned(43,8) ,
68291	 => std_logic_vector(to_unsigned(87,8) ,
68292	 => std_logic_vector(to_unsigned(108,8) ,
68293	 => std_logic_vector(to_unsigned(107,8) ,
68294	 => std_logic_vector(to_unsigned(116,8) ,
68295	 => std_logic_vector(to_unsigned(118,8) ,
68296	 => std_logic_vector(to_unsigned(104,8) ,
68297	 => std_logic_vector(to_unsigned(114,8) ,
68298	 => std_logic_vector(to_unsigned(116,8) ,
68299	 => std_logic_vector(to_unsigned(72,8) ,
68300	 => std_logic_vector(to_unsigned(62,8) ,
68301	 => std_logic_vector(to_unsigned(42,8) ,
68302	 => std_logic_vector(to_unsigned(16,8) ,
68303	 => std_logic_vector(to_unsigned(45,8) ,
68304	 => std_logic_vector(to_unsigned(23,8) ,
68305	 => std_logic_vector(to_unsigned(23,8) ,
68306	 => std_logic_vector(to_unsigned(72,8) ,
68307	 => std_logic_vector(to_unsigned(52,8) ,
68308	 => std_logic_vector(to_unsigned(13,8) ,
68309	 => std_logic_vector(to_unsigned(32,8) ,
68310	 => std_logic_vector(to_unsigned(47,8) ,
68311	 => std_logic_vector(to_unsigned(47,8) ,
68312	 => std_logic_vector(to_unsigned(50,8) ,
68313	 => std_logic_vector(to_unsigned(42,8) ,
68314	 => std_logic_vector(to_unsigned(37,8) ,
68315	 => std_logic_vector(to_unsigned(57,8) ,
68316	 => std_logic_vector(to_unsigned(39,8) ,
68317	 => std_logic_vector(to_unsigned(8,8) ,
68318	 => std_logic_vector(to_unsigned(6,8) ,
68319	 => std_logic_vector(to_unsigned(6,8) ,
68320	 => std_logic_vector(to_unsigned(8,8) ,
68321	 => std_logic_vector(to_unsigned(23,8) ,
68322	 => std_logic_vector(to_unsigned(13,8) ,
68323	 => std_logic_vector(to_unsigned(9,8) ,
68324	 => std_logic_vector(to_unsigned(27,8) ,
68325	 => std_logic_vector(to_unsigned(23,8) ,
68326	 => std_logic_vector(to_unsigned(12,8) ,
68327	 => std_logic_vector(to_unsigned(5,8) ,
68328	 => std_logic_vector(to_unsigned(10,8) ,
68329	 => std_logic_vector(to_unsigned(34,8) ,
68330	 => std_logic_vector(to_unsigned(24,8) ,
68331	 => std_logic_vector(to_unsigned(16,8) ,
68332	 => std_logic_vector(to_unsigned(23,8) ,
68333	 => std_logic_vector(to_unsigned(33,8) ,
68334	 => std_logic_vector(to_unsigned(15,8) ,
68335	 => std_logic_vector(to_unsigned(31,8) ,
68336	 => std_logic_vector(to_unsigned(67,8) ,
68337	 => std_logic_vector(to_unsigned(34,8) ,
68338	 => std_logic_vector(to_unsigned(23,8) ,
68339	 => std_logic_vector(to_unsigned(27,8) ,
68340	 => std_logic_vector(to_unsigned(22,8) ,
68341	 => std_logic_vector(to_unsigned(12,8) ,
68342	 => std_logic_vector(to_unsigned(17,8) ,
68343	 => std_logic_vector(to_unsigned(30,8) ,
68344	 => std_logic_vector(to_unsigned(25,8) ,
68345	 => std_logic_vector(to_unsigned(15,8) ,
68346	 => std_logic_vector(to_unsigned(33,8) ,
68347	 => std_logic_vector(to_unsigned(26,8) ,
68348	 => std_logic_vector(to_unsigned(12,8) ,
68349	 => std_logic_vector(to_unsigned(18,8) ,
68350	 => std_logic_vector(to_unsigned(34,8) ,
68351	 => std_logic_vector(to_unsigned(37,8) ,
68352	 => std_logic_vector(to_unsigned(31,8) ,
68353	 => std_logic_vector(to_unsigned(32,8) ,
68354	 => std_logic_vector(to_unsigned(41,8) ,
68355	 => std_logic_vector(to_unsigned(38,8) ,
68356	 => std_logic_vector(to_unsigned(37,8) ,
68357	 => std_logic_vector(to_unsigned(45,8) ,
68358	 => std_logic_vector(to_unsigned(67,8) ,
68359	 => std_logic_vector(to_unsigned(67,8) ,
68360	 => std_logic_vector(to_unsigned(37,8) ,
68361	 => std_logic_vector(to_unsigned(27,8) ,
68362	 => std_logic_vector(to_unsigned(16,8) ,
68363	 => std_logic_vector(to_unsigned(11,8) ,
68364	 => std_logic_vector(to_unsigned(20,8) ,
68365	 => std_logic_vector(to_unsigned(19,8) ,
68366	 => std_logic_vector(to_unsigned(12,8) ,
68367	 => std_logic_vector(to_unsigned(9,8) ,
68368	 => std_logic_vector(to_unsigned(24,8) ,
68369	 => std_logic_vector(to_unsigned(41,8) ,
68370	 => std_logic_vector(to_unsigned(61,8) ,
68371	 => std_logic_vector(to_unsigned(44,8) ,
68372	 => std_logic_vector(to_unsigned(25,8) ,
68373	 => std_logic_vector(to_unsigned(32,8) ,
68374	 => std_logic_vector(to_unsigned(40,8) ,
68375	 => std_logic_vector(to_unsigned(43,8) ,
68376	 => std_logic_vector(to_unsigned(39,8) ,
68377	 => std_logic_vector(to_unsigned(26,8) ,
68378	 => std_logic_vector(to_unsigned(27,8) ,
68379	 => std_logic_vector(to_unsigned(35,8) ,
68380	 => std_logic_vector(to_unsigned(46,8) ,
68381	 => std_logic_vector(to_unsigned(40,8) ,
68382	 => std_logic_vector(to_unsigned(25,8) ,
68383	 => std_logic_vector(to_unsigned(27,8) ,
68384	 => std_logic_vector(to_unsigned(48,8) ,
68385	 => std_logic_vector(to_unsigned(37,8) ,
68386	 => std_logic_vector(to_unsigned(32,8) ,
68387	 => std_logic_vector(to_unsigned(32,8) ,
68388	 => std_logic_vector(to_unsigned(20,8) ,
68389	 => std_logic_vector(to_unsigned(4,8) ,
68390	 => std_logic_vector(to_unsigned(10,8) ,
68391	 => std_logic_vector(to_unsigned(45,8) ,
68392	 => std_logic_vector(to_unsigned(25,8) ,
68393	 => std_logic_vector(to_unsigned(30,8) ,
68394	 => std_logic_vector(to_unsigned(44,8) ,
68395	 => std_logic_vector(to_unsigned(58,8) ,
68396	 => std_logic_vector(to_unsigned(29,8) ,
68397	 => std_logic_vector(to_unsigned(19,8) ,
68398	 => std_logic_vector(to_unsigned(68,8) ,
68399	 => std_logic_vector(to_unsigned(74,8) ,
68400	 => std_logic_vector(to_unsigned(46,8) ,
68401	 => std_logic_vector(to_unsigned(13,8) ,
68402	 => std_logic_vector(to_unsigned(32,8) ,
68403	 => std_logic_vector(to_unsigned(69,8) ,
68404	 => std_logic_vector(to_unsigned(95,8) ,
68405	 => std_logic_vector(to_unsigned(112,8) ,
68406	 => std_logic_vector(to_unsigned(49,8) ,
68407	 => std_logic_vector(to_unsigned(57,8) ,
68408	 => std_logic_vector(to_unsigned(127,8) ,
68409	 => std_logic_vector(to_unsigned(111,8) ,
68410	 => std_logic_vector(to_unsigned(78,8) ,
68411	 => std_logic_vector(to_unsigned(48,8) ,
68412	 => std_logic_vector(to_unsigned(24,8) ,
68413	 => std_logic_vector(to_unsigned(37,8) ,
68414	 => std_logic_vector(to_unsigned(48,8) ,
68415	 => std_logic_vector(to_unsigned(42,8) ,
68416	 => std_logic_vector(to_unsigned(45,8) ,
68417	 => std_logic_vector(to_unsigned(37,8) ,
68418	 => std_logic_vector(to_unsigned(31,8) ,
68419	 => std_logic_vector(to_unsigned(28,8) ,
68420	 => std_logic_vector(to_unsigned(29,8) ,
68421	 => std_logic_vector(to_unsigned(21,8) ,
68422	 => std_logic_vector(to_unsigned(29,8) ,
68423	 => std_logic_vector(to_unsigned(40,8) ,
68424	 => std_logic_vector(to_unsigned(34,8) ,
68425	 => std_logic_vector(to_unsigned(32,8) ,
68426	 => std_logic_vector(to_unsigned(39,8) ,
68427	 => std_logic_vector(to_unsigned(43,8) ,
68428	 => std_logic_vector(to_unsigned(35,8) ,
68429	 => std_logic_vector(to_unsigned(13,8) ,
68430	 => std_logic_vector(to_unsigned(29,8) ,
68431	 => std_logic_vector(to_unsigned(50,8) ,
68432	 => std_logic_vector(to_unsigned(18,8) ,
68433	 => std_logic_vector(to_unsigned(12,8) ,
68434	 => std_logic_vector(to_unsigned(1,8) ,
68435	 => std_logic_vector(to_unsigned(0,8) ,
68436	 => std_logic_vector(to_unsigned(5,8) ,
68437	 => std_logic_vector(to_unsigned(8,8) ,
68438	 => std_logic_vector(to_unsigned(6,8) ,
68439	 => std_logic_vector(to_unsigned(7,8) ,
68440	 => std_logic_vector(to_unsigned(8,8) ,
68441	 => std_logic_vector(to_unsigned(8,8) ,
68442	 => std_logic_vector(to_unsigned(8,8) ,
68443	 => std_logic_vector(to_unsigned(8,8) ,
68444	 => std_logic_vector(to_unsigned(6,8) ,
68445	 => std_logic_vector(to_unsigned(1,8) ,
68446	 => std_logic_vector(to_unsigned(0,8) ,
68447	 => std_logic_vector(to_unsigned(1,8) ,
68448	 => std_logic_vector(to_unsigned(12,8) ,
68449	 => std_logic_vector(to_unsigned(16,8) ,
68450	 => std_logic_vector(to_unsigned(9,8) ,
68451	 => std_logic_vector(to_unsigned(25,8) ,
68452	 => std_logic_vector(to_unsigned(100,8) ,
68453	 => std_logic_vector(to_unsigned(92,8) ,
68454	 => std_logic_vector(to_unsigned(95,8) ,
68455	 => std_logic_vector(to_unsigned(51,8) ,
68456	 => std_logic_vector(to_unsigned(37,8) ,
68457	 => std_logic_vector(to_unsigned(32,8) ,
68458	 => std_logic_vector(to_unsigned(54,8) ,
68459	 => std_logic_vector(to_unsigned(29,8) ,
68460	 => std_logic_vector(to_unsigned(1,8) ,
68461	 => std_logic_vector(to_unsigned(0,8) ,
68462	 => std_logic_vector(to_unsigned(8,8) ,
68463	 => std_logic_vector(to_unsigned(37,8) ,
68464	 => std_logic_vector(to_unsigned(42,8) ,
68465	 => std_logic_vector(to_unsigned(97,8) ,
68466	 => std_logic_vector(to_unsigned(24,8) ,
68467	 => std_logic_vector(to_unsigned(32,8) ,
68468	 => std_logic_vector(to_unsigned(42,8) ,
68469	 => std_logic_vector(to_unsigned(8,8) ,
68470	 => std_logic_vector(to_unsigned(9,8) ,
68471	 => std_logic_vector(to_unsigned(8,8) ,
68472	 => std_logic_vector(to_unsigned(7,8) ,
68473	 => std_logic_vector(to_unsigned(9,8) ,
68474	 => std_logic_vector(to_unsigned(10,8) ,
68475	 => std_logic_vector(to_unsigned(17,8) ,
68476	 => std_logic_vector(to_unsigned(32,8) ,
68477	 => std_logic_vector(to_unsigned(39,8) ,
68478	 => std_logic_vector(to_unsigned(48,8) ,
68479	 => std_logic_vector(to_unsigned(55,8) ,
68480	 => std_logic_vector(to_unsigned(69,8) ,
68481	 => std_logic_vector(to_unsigned(97,8) ,
68482	 => std_logic_vector(to_unsigned(100,8) ,
68483	 => std_logic_vector(to_unsigned(100,8) ,
68484	 => std_logic_vector(to_unsigned(103,8) ,
68485	 => std_logic_vector(to_unsigned(88,8) ,
68486	 => std_logic_vector(to_unsigned(107,8) ,
68487	 => std_logic_vector(to_unsigned(114,8) ,
68488	 => std_logic_vector(to_unsigned(100,8) ,
68489	 => std_logic_vector(to_unsigned(97,8) ,
68490	 => std_logic_vector(to_unsigned(105,8) ,
68491	 => std_logic_vector(to_unsigned(81,8) ,
68492	 => std_logic_vector(to_unsigned(43,8) ,
68493	 => std_logic_vector(to_unsigned(43,8) ,
68494	 => std_logic_vector(to_unsigned(43,8) ,
68495	 => std_logic_vector(to_unsigned(46,8) ,
68496	 => std_logic_vector(to_unsigned(53,8) ,
68497	 => std_logic_vector(to_unsigned(70,8) ,
68498	 => std_logic_vector(to_unsigned(63,8) ,
68499	 => std_logic_vector(to_unsigned(52,8) ,
68500	 => std_logic_vector(to_unsigned(51,8) ,
68501	 => std_logic_vector(to_unsigned(47,8) ,
68502	 => std_logic_vector(to_unsigned(44,8) ,
68503	 => std_logic_vector(to_unsigned(35,8) ,
68504	 => std_logic_vector(to_unsigned(25,8) ,
68505	 => std_logic_vector(to_unsigned(25,8) ,
68506	 => std_logic_vector(to_unsigned(43,8) ,
68507	 => std_logic_vector(to_unsigned(55,8) ,
68508	 => std_logic_vector(to_unsigned(43,8) ,
68509	 => std_logic_vector(to_unsigned(35,8) ,
68510	 => std_logic_vector(to_unsigned(37,8) ,
68511	 => std_logic_vector(to_unsigned(33,8) ,
68512	 => std_logic_vector(to_unsigned(33,8) ,
68513	 => std_logic_vector(to_unsigned(29,8) ,
68514	 => std_logic_vector(to_unsigned(26,8) ,
68515	 => std_logic_vector(to_unsigned(27,8) ,
68516	 => std_logic_vector(to_unsigned(32,8) ,
68517	 => std_logic_vector(to_unsigned(38,8) ,
68518	 => std_logic_vector(to_unsigned(63,8) ,
68519	 => std_logic_vector(to_unsigned(73,8) ,
68520	 => std_logic_vector(to_unsigned(37,8) ,
68521	 => std_logic_vector(to_unsigned(35,8) ,
68522	 => std_logic_vector(to_unsigned(56,8) ,
68523	 => std_logic_vector(to_unsigned(74,8) ,
68524	 => std_logic_vector(to_unsigned(51,8) ,
68525	 => std_logic_vector(to_unsigned(37,8) ,
68526	 => std_logic_vector(to_unsigned(32,8) ,
68527	 => std_logic_vector(to_unsigned(39,8) ,
68528	 => std_logic_vector(to_unsigned(52,8) ,
68529	 => std_logic_vector(to_unsigned(37,8) ,
68530	 => std_logic_vector(to_unsigned(32,8) ,
68531	 => std_logic_vector(to_unsigned(34,8) ,
68532	 => std_logic_vector(to_unsigned(40,8) ,
68533	 => std_logic_vector(to_unsigned(69,8) ,
68534	 => std_logic_vector(to_unsigned(85,8) ,
68535	 => std_logic_vector(to_unsigned(99,8) ,
68536	 => std_logic_vector(to_unsigned(88,8) ,
68537	 => std_logic_vector(to_unsigned(72,8) ,
68538	 => std_logic_vector(to_unsigned(57,8) ,
68539	 => std_logic_vector(to_unsigned(35,8) ,
68540	 => std_logic_vector(to_unsigned(40,8) ,
68541	 => std_logic_vector(to_unsigned(37,8) ,
68542	 => std_logic_vector(to_unsigned(39,8) ,
68543	 => std_logic_vector(to_unsigned(34,8) ,
68544	 => std_logic_vector(to_unsigned(35,8) ,
68545	 => std_logic_vector(to_unsigned(35,8) ,
68546	 => std_logic_vector(to_unsigned(68,8) ,
68547	 => std_logic_vector(to_unsigned(100,8) ,
68548	 => std_logic_vector(to_unsigned(91,8) ,
68549	 => std_logic_vector(to_unsigned(100,8) ,
68550	 => std_logic_vector(to_unsigned(97,8) ,
68551	 => std_logic_vector(to_unsigned(97,8) ,
68552	 => std_logic_vector(to_unsigned(99,8) ,
68553	 => std_logic_vector(to_unsigned(95,8) ,
68554	 => std_logic_vector(to_unsigned(79,8) ,
68555	 => std_logic_vector(to_unsigned(78,8) ,
68556	 => std_logic_vector(to_unsigned(90,8) ,
68557	 => std_logic_vector(to_unsigned(88,8) ,
68558	 => std_logic_vector(to_unsigned(87,8) ,
68559	 => std_logic_vector(to_unsigned(78,8) ,
68560	 => std_logic_vector(to_unsigned(93,8) ,
68561	 => std_logic_vector(to_unsigned(96,8) ,
68562	 => std_logic_vector(to_unsigned(79,8) ,
68563	 => std_logic_vector(to_unsigned(97,8) ,
68564	 => std_logic_vector(to_unsigned(88,8) ,
68565	 => std_logic_vector(to_unsigned(79,8) ,
68566	 => std_logic_vector(to_unsigned(76,8) ,
68567	 => std_logic_vector(to_unsigned(73,8) ,
68568	 => std_logic_vector(to_unsigned(43,8) ,
68569	 => std_logic_vector(to_unsigned(20,8) ,
68570	 => std_logic_vector(to_unsigned(23,8) ,
68571	 => std_logic_vector(to_unsigned(24,8) ,
68572	 => std_logic_vector(to_unsigned(36,8) ,
68573	 => std_logic_vector(to_unsigned(35,8) ,
68574	 => std_logic_vector(to_unsigned(35,8) ,
68575	 => std_logic_vector(to_unsigned(41,8) ,
68576	 => std_logic_vector(to_unsigned(48,8) ,
68577	 => std_logic_vector(to_unsigned(46,8) ,
68578	 => std_logic_vector(to_unsigned(49,8) ,
68579	 => std_logic_vector(to_unsigned(43,8) ,
68580	 => std_logic_vector(to_unsigned(46,8) ,
68581	 => std_logic_vector(to_unsigned(48,8) ,
68582	 => std_logic_vector(to_unsigned(50,8) ,
68583	 => std_logic_vector(to_unsigned(27,8) ,
68584	 => std_logic_vector(to_unsigned(19,8) ,
68585	 => std_logic_vector(to_unsigned(22,8) ,
68586	 => std_logic_vector(to_unsigned(19,8) ,
68587	 => std_logic_vector(to_unsigned(14,8) ,
68588	 => std_logic_vector(to_unsigned(14,8) ,
68589	 => std_logic_vector(to_unsigned(31,8) ,
68590	 => std_logic_vector(to_unsigned(51,8) ,
68591	 => std_logic_vector(to_unsigned(41,8) ,
68592	 => std_logic_vector(to_unsigned(37,8) ,
68593	 => std_logic_vector(to_unsigned(78,8) ,
68594	 => std_logic_vector(to_unsigned(82,8) ,
68595	 => std_logic_vector(to_unsigned(42,8) ,
68596	 => std_logic_vector(to_unsigned(95,8) ,
68597	 => std_logic_vector(to_unsigned(119,8) ,
68598	 => std_logic_vector(to_unsigned(82,8) ,
68599	 => std_logic_vector(to_unsigned(66,8) ,
68600	 => std_logic_vector(to_unsigned(85,8) ,
68601	 => std_logic_vector(to_unsigned(92,8) ,
68602	 => std_logic_vector(to_unsigned(73,8) ,
68603	 => std_logic_vector(to_unsigned(51,8) ,
68604	 => std_logic_vector(to_unsigned(45,8) ,
68605	 => std_logic_vector(to_unsigned(37,8) ,
68606	 => std_logic_vector(to_unsigned(30,8) ,
68607	 => std_logic_vector(to_unsigned(27,8) ,
68608	 => std_logic_vector(to_unsigned(28,8) ,
68609	 => std_logic_vector(to_unsigned(52,8) ,
68610	 => std_logic_vector(to_unsigned(90,8) ,
68611	 => std_logic_vector(to_unsigned(104,8) ,
68612	 => std_logic_vector(to_unsigned(122,8) ,
68613	 => std_logic_vector(to_unsigned(115,8) ,
68614	 => std_logic_vector(to_unsigned(114,8) ,
68615	 => std_logic_vector(to_unsigned(116,8) ,
68616	 => std_logic_vector(to_unsigned(97,8) ,
68617	 => std_logic_vector(to_unsigned(58,8) ,
68618	 => std_logic_vector(to_unsigned(53,8) ,
68619	 => std_logic_vector(to_unsigned(56,8) ,
68620	 => std_logic_vector(to_unsigned(60,8) ,
68621	 => std_logic_vector(to_unsigned(47,8) ,
68622	 => std_logic_vector(to_unsigned(23,8) ,
68623	 => std_logic_vector(to_unsigned(38,8) ,
68624	 => std_logic_vector(to_unsigned(28,8) ,
68625	 => std_logic_vector(to_unsigned(15,8) ,
68626	 => std_logic_vector(to_unsigned(63,8) ,
68627	 => std_logic_vector(to_unsigned(38,8) ,
68628	 => std_logic_vector(to_unsigned(6,8) ,
68629	 => std_logic_vector(to_unsigned(33,8) ,
68630	 => std_logic_vector(to_unsigned(37,8) ,
68631	 => std_logic_vector(to_unsigned(21,8) ,
68632	 => std_logic_vector(to_unsigned(46,8) ,
68633	 => std_logic_vector(to_unsigned(44,8) ,
68634	 => std_logic_vector(to_unsigned(41,8) ,
68635	 => std_logic_vector(to_unsigned(52,8) ,
68636	 => std_logic_vector(to_unsigned(35,8) ,
68637	 => std_logic_vector(to_unsigned(7,8) ,
68638	 => std_logic_vector(to_unsigned(4,8) ,
68639	 => std_logic_vector(to_unsigned(8,8) ,
68640	 => std_logic_vector(to_unsigned(6,8) ,
68641	 => std_logic_vector(to_unsigned(17,8) ,
68642	 => std_logic_vector(to_unsigned(13,8) ,
68643	 => std_logic_vector(to_unsigned(9,8) ,
68644	 => std_logic_vector(to_unsigned(20,8) ,
68645	 => std_logic_vector(to_unsigned(17,8) ,
68646	 => std_logic_vector(to_unsigned(10,8) ,
68647	 => std_logic_vector(to_unsigned(5,8) ,
68648	 => std_logic_vector(to_unsigned(10,8) ,
68649	 => std_logic_vector(to_unsigned(30,8) ,
68650	 => std_logic_vector(to_unsigned(20,8) ,
68651	 => std_logic_vector(to_unsigned(23,8) ,
68652	 => std_logic_vector(to_unsigned(31,8) ,
68653	 => std_logic_vector(to_unsigned(19,8) ,
68654	 => std_logic_vector(to_unsigned(31,8) ,
68655	 => std_logic_vector(to_unsigned(60,8) ,
68656	 => std_logic_vector(to_unsigned(30,8) ,
68657	 => std_logic_vector(to_unsigned(38,8) ,
68658	 => std_logic_vector(to_unsigned(27,8) ,
68659	 => std_logic_vector(to_unsigned(24,8) ,
68660	 => std_logic_vector(to_unsigned(29,8) ,
68661	 => std_logic_vector(to_unsigned(12,8) ,
68662	 => std_logic_vector(to_unsigned(12,8) ,
68663	 => std_logic_vector(to_unsigned(19,8) ,
68664	 => std_logic_vector(to_unsigned(20,8) ,
68665	 => std_logic_vector(to_unsigned(23,8) ,
68666	 => std_logic_vector(to_unsigned(41,8) ,
68667	 => std_logic_vector(to_unsigned(45,8) ,
68668	 => std_logic_vector(to_unsigned(43,8) ,
68669	 => std_logic_vector(to_unsigned(35,8) ,
68670	 => std_logic_vector(to_unsigned(35,8) ,
68671	 => std_logic_vector(to_unsigned(39,8) ,
68672	 => std_logic_vector(to_unsigned(21,8) ,
68673	 => std_logic_vector(to_unsigned(12,8) ,
68674	 => std_logic_vector(to_unsigned(22,8) ,
68675	 => std_logic_vector(to_unsigned(40,8) ,
68676	 => std_logic_vector(to_unsigned(38,8) ,
68677	 => std_logic_vector(to_unsigned(43,8) ,
68678	 => std_logic_vector(to_unsigned(56,8) ,
68679	 => std_logic_vector(to_unsigned(45,8) ,
68680	 => std_logic_vector(to_unsigned(41,8) ,
68681	 => std_logic_vector(to_unsigned(20,8) ,
68682	 => std_logic_vector(to_unsigned(16,8) ,
68683	 => std_logic_vector(to_unsigned(16,8) ,
68684	 => std_logic_vector(to_unsigned(13,8) ,
68685	 => std_logic_vector(to_unsigned(16,8) ,
68686	 => std_logic_vector(to_unsigned(11,8) ,
68687	 => std_logic_vector(to_unsigned(10,8) ,
68688	 => std_logic_vector(to_unsigned(19,8) ,
68689	 => std_logic_vector(to_unsigned(55,8) ,
68690	 => std_logic_vector(to_unsigned(107,8) ,
68691	 => std_logic_vector(to_unsigned(79,8) ,
68692	 => std_logic_vector(to_unsigned(29,8) ,
68693	 => std_logic_vector(to_unsigned(24,8) ,
68694	 => std_logic_vector(to_unsigned(37,8) ,
68695	 => std_logic_vector(to_unsigned(50,8) ,
68696	 => std_logic_vector(to_unsigned(44,8) ,
68697	 => std_logic_vector(to_unsigned(29,8) ,
68698	 => std_logic_vector(to_unsigned(24,8) ,
68699	 => std_logic_vector(to_unsigned(29,8) ,
68700	 => std_logic_vector(to_unsigned(45,8) ,
68701	 => std_logic_vector(to_unsigned(50,8) ,
68702	 => std_logic_vector(to_unsigned(28,8) ,
68703	 => std_logic_vector(to_unsigned(27,8) ,
68704	 => std_logic_vector(to_unsigned(37,8) ,
68705	 => std_logic_vector(to_unsigned(31,8) ,
68706	 => std_logic_vector(to_unsigned(35,8) ,
68707	 => std_logic_vector(to_unsigned(29,8) ,
68708	 => std_logic_vector(to_unsigned(16,8) ,
68709	 => std_logic_vector(to_unsigned(4,8) ,
68710	 => std_logic_vector(to_unsigned(11,8) ,
68711	 => std_logic_vector(to_unsigned(48,8) ,
68712	 => std_logic_vector(to_unsigned(41,8) ,
68713	 => std_logic_vector(to_unsigned(33,8) ,
68714	 => std_logic_vector(to_unsigned(35,8) ,
68715	 => std_logic_vector(to_unsigned(50,8) ,
68716	 => std_logic_vector(to_unsigned(51,8) ,
68717	 => std_logic_vector(to_unsigned(63,8) ,
68718	 => std_logic_vector(to_unsigned(72,8) ,
68719	 => std_logic_vector(to_unsigned(65,8) ,
68720	 => std_logic_vector(to_unsigned(51,8) ,
68721	 => std_logic_vector(to_unsigned(45,8) ,
68722	 => std_logic_vector(to_unsigned(47,8) ,
68723	 => std_logic_vector(to_unsigned(71,8) ,
68724	 => std_logic_vector(to_unsigned(107,8) ,
68725	 => std_logic_vector(to_unsigned(111,8) ,
68726	 => std_logic_vector(to_unsigned(48,8) ,
68727	 => std_logic_vector(to_unsigned(57,8) ,
68728	 => std_logic_vector(to_unsigned(124,8) ,
68729	 => std_logic_vector(to_unsigned(115,8) ,
68730	 => std_logic_vector(to_unsigned(59,8) ,
68731	 => std_logic_vector(to_unsigned(27,8) ,
68732	 => std_logic_vector(to_unsigned(26,8) ,
68733	 => std_logic_vector(to_unsigned(44,8) ,
68734	 => std_logic_vector(to_unsigned(48,8) ,
68735	 => std_logic_vector(to_unsigned(51,8) ,
68736	 => std_logic_vector(to_unsigned(56,8) ,
68737	 => std_logic_vector(to_unsigned(31,8) ,
68738	 => std_logic_vector(to_unsigned(36,8) ,
68739	 => std_logic_vector(to_unsigned(49,8) ,
68740	 => std_logic_vector(to_unsigned(45,8) ,
68741	 => std_logic_vector(to_unsigned(34,8) ,
68742	 => std_logic_vector(to_unsigned(43,8) ,
68743	 => std_logic_vector(to_unsigned(65,8) ,
68744	 => std_logic_vector(to_unsigned(58,8) ,
68745	 => std_logic_vector(to_unsigned(54,8) ,
68746	 => std_logic_vector(to_unsigned(42,8) ,
68747	 => std_logic_vector(to_unsigned(56,8) ,
68748	 => std_logic_vector(to_unsigned(44,8) ,
68749	 => std_logic_vector(to_unsigned(8,8) ,
68750	 => std_logic_vector(to_unsigned(17,8) ,
68751	 => std_logic_vector(to_unsigned(20,8) ,
68752	 => std_logic_vector(to_unsigned(7,8) ,
68753	 => std_logic_vector(to_unsigned(15,8) ,
68754	 => std_logic_vector(to_unsigned(1,8) ,
68755	 => std_logic_vector(to_unsigned(0,8) ,
68756	 => std_logic_vector(to_unsigned(4,8) ,
68757	 => std_logic_vector(to_unsigned(7,8) ,
68758	 => std_logic_vector(to_unsigned(9,8) ,
68759	 => std_logic_vector(to_unsigned(13,8) ,
68760	 => std_logic_vector(to_unsigned(6,8) ,
68761	 => std_logic_vector(to_unsigned(7,8) ,
68762	 => std_logic_vector(to_unsigned(5,8) ,
68763	 => std_logic_vector(to_unsigned(5,8) ,
68764	 => std_logic_vector(to_unsigned(8,8) ,
68765	 => std_logic_vector(to_unsigned(2,8) ,
68766	 => std_logic_vector(to_unsigned(0,8) ,
68767	 => std_logic_vector(to_unsigned(1,8) ,
68768	 => std_logic_vector(to_unsigned(19,8) ,
68769	 => std_logic_vector(to_unsigned(37,8) ,
68770	 => std_logic_vector(to_unsigned(37,8) ,
68771	 => std_logic_vector(to_unsigned(67,8) ,
68772	 => std_logic_vector(to_unsigned(104,8) ,
68773	 => std_logic_vector(to_unsigned(87,8) ,
68774	 => std_logic_vector(to_unsigned(79,8) ,
68775	 => std_logic_vector(to_unsigned(37,8) ,
68776	 => std_logic_vector(to_unsigned(41,8) ,
68777	 => std_logic_vector(to_unsigned(17,8) ,
68778	 => std_logic_vector(to_unsigned(58,8) ,
68779	 => std_logic_vector(to_unsigned(26,8) ,
68780	 => std_logic_vector(to_unsigned(2,8) ,
68781	 => std_logic_vector(to_unsigned(0,8) ,
68782	 => std_logic_vector(to_unsigned(4,8) ,
68783	 => std_logic_vector(to_unsigned(17,8) ,
68784	 => std_logic_vector(to_unsigned(41,8) ,
68785	 => std_logic_vector(to_unsigned(101,8) ,
68786	 => std_logic_vector(to_unsigned(27,8) ,
68787	 => std_logic_vector(to_unsigned(40,8) ,
68788	 => std_logic_vector(to_unsigned(35,8) ,
68789	 => std_logic_vector(to_unsigned(9,8) ,
68790	 => std_logic_vector(to_unsigned(13,8) ,
68791	 => std_logic_vector(to_unsigned(13,8) ,
68792	 => std_logic_vector(to_unsigned(10,8) ,
68793	 => std_logic_vector(to_unsigned(12,8) ,
68794	 => std_logic_vector(to_unsigned(7,8) ,
68795	 => std_logic_vector(to_unsigned(9,8) ,
68796	 => std_logic_vector(to_unsigned(18,8) ,
68797	 => std_logic_vector(to_unsigned(8,8) ,
68798	 => std_logic_vector(to_unsigned(8,8) ,
68799	 => std_logic_vector(to_unsigned(11,8) ,
68800	 => std_logic_vector(to_unsigned(13,8) ,
68801	 => std_logic_vector(to_unsigned(101,8) ,
68802	 => std_logic_vector(to_unsigned(105,8) ,
68803	 => std_logic_vector(to_unsigned(103,8) ,
68804	 => std_logic_vector(to_unsigned(104,8) ,
68805	 => std_logic_vector(to_unsigned(97,8) ,
68806	 => std_logic_vector(to_unsigned(122,8) ,
68807	 => std_logic_vector(to_unsigned(121,8) ,
68808	 => std_logic_vector(to_unsigned(88,8) ,
68809	 => std_logic_vector(to_unsigned(95,8) ,
68810	 => std_logic_vector(to_unsigned(112,8) ,
68811	 => std_logic_vector(to_unsigned(74,8) ,
68812	 => std_logic_vector(to_unsigned(42,8) ,
68813	 => std_logic_vector(to_unsigned(54,8) ,
68814	 => std_logic_vector(to_unsigned(63,8) ,
68815	 => std_logic_vector(to_unsigned(66,8) ,
68816	 => std_logic_vector(to_unsigned(66,8) ,
68817	 => std_logic_vector(to_unsigned(79,8) ,
68818	 => std_logic_vector(to_unsigned(64,8) ,
68819	 => std_logic_vector(to_unsigned(59,8) ,
68820	 => std_logic_vector(to_unsigned(66,8) ,
68821	 => std_logic_vector(to_unsigned(46,8) ,
68822	 => std_logic_vector(to_unsigned(45,8) ,
68823	 => std_logic_vector(to_unsigned(31,8) ,
68824	 => std_logic_vector(to_unsigned(18,8) ,
68825	 => std_logic_vector(to_unsigned(25,8) ,
68826	 => std_logic_vector(to_unsigned(48,8) ,
68827	 => std_logic_vector(to_unsigned(37,8) ,
68828	 => std_logic_vector(to_unsigned(31,8) ,
68829	 => std_logic_vector(to_unsigned(34,8) ,
68830	 => std_logic_vector(to_unsigned(37,8) ,
68831	 => std_logic_vector(to_unsigned(39,8) ,
68832	 => std_logic_vector(to_unsigned(41,8) ,
68833	 => std_logic_vector(to_unsigned(29,8) ,
68834	 => std_logic_vector(to_unsigned(27,8) ,
68835	 => std_logic_vector(to_unsigned(45,8) ,
68836	 => std_logic_vector(to_unsigned(68,8) ,
68837	 => std_logic_vector(to_unsigned(80,8) ,
68838	 => std_logic_vector(to_unsigned(84,8) ,
68839	 => std_logic_vector(to_unsigned(78,8) ,
68840	 => std_logic_vector(to_unsigned(69,8) ,
68841	 => std_logic_vector(to_unsigned(55,8) ,
68842	 => std_logic_vector(to_unsigned(40,8) ,
68843	 => std_logic_vector(to_unsigned(37,8) ,
68844	 => std_logic_vector(to_unsigned(35,8) ,
68845	 => std_logic_vector(to_unsigned(39,8) ,
68846	 => std_logic_vector(to_unsigned(51,8) ,
68847	 => std_logic_vector(to_unsigned(53,8) ,
68848	 => std_logic_vector(to_unsigned(54,8) ,
68849	 => std_logic_vector(to_unsigned(41,8) ,
68850	 => std_logic_vector(to_unsigned(32,8) ,
68851	 => std_logic_vector(to_unsigned(28,8) ,
68852	 => std_logic_vector(to_unsigned(26,8) ,
68853	 => std_logic_vector(to_unsigned(39,8) ,
68854	 => std_logic_vector(to_unsigned(61,8) ,
68855	 => std_logic_vector(to_unsigned(80,8) ,
68856	 => std_logic_vector(to_unsigned(87,8) ,
68857	 => std_logic_vector(to_unsigned(81,8) ,
68858	 => std_logic_vector(to_unsigned(60,8) ,
68859	 => std_logic_vector(to_unsigned(42,8) ,
68860	 => std_logic_vector(to_unsigned(41,8) ,
68861	 => std_logic_vector(to_unsigned(45,8) ,
68862	 => std_logic_vector(to_unsigned(37,8) ,
68863	 => std_logic_vector(to_unsigned(29,8) ,
68864	 => std_logic_vector(to_unsigned(37,8) ,
68865	 => std_logic_vector(to_unsigned(38,8) ,
68866	 => std_logic_vector(to_unsigned(66,8) ,
68867	 => std_logic_vector(to_unsigned(100,8) ,
68868	 => std_logic_vector(to_unsigned(93,8) ,
68869	 => std_logic_vector(to_unsigned(93,8) ,
68870	 => std_logic_vector(to_unsigned(99,8) ,
68871	 => std_logic_vector(to_unsigned(99,8) ,
68872	 => std_logic_vector(to_unsigned(95,8) ,
68873	 => std_logic_vector(to_unsigned(77,8) ,
68874	 => std_logic_vector(to_unsigned(69,8) ,
68875	 => std_logic_vector(to_unsigned(77,8) ,
68876	 => std_logic_vector(to_unsigned(57,8) ,
68877	 => std_logic_vector(to_unsigned(62,8) ,
68878	 => std_logic_vector(to_unsigned(88,8) ,
68879	 => std_logic_vector(to_unsigned(73,8) ,
68880	 => std_logic_vector(to_unsigned(81,8) ,
68881	 => std_logic_vector(to_unsigned(72,8) ,
68882	 => std_logic_vector(to_unsigned(52,8) ,
68883	 => std_logic_vector(to_unsigned(100,8) ,
68884	 => std_logic_vector(to_unsigned(82,8) ,
68885	 => std_logic_vector(to_unsigned(74,8) ,
68886	 => std_logic_vector(to_unsigned(76,8) ,
68887	 => std_logic_vector(to_unsigned(74,8) ,
68888	 => std_logic_vector(to_unsigned(45,8) ,
68889	 => std_logic_vector(to_unsigned(33,8) ,
68890	 => std_logic_vector(to_unsigned(33,8) ,
68891	 => std_logic_vector(to_unsigned(19,8) ,
68892	 => std_logic_vector(to_unsigned(35,8) ,
68893	 => std_logic_vector(to_unsigned(39,8) ,
68894	 => std_logic_vector(to_unsigned(31,8) ,
68895	 => std_logic_vector(to_unsigned(35,8) ,
68896	 => std_logic_vector(to_unsigned(44,8) ,
68897	 => std_logic_vector(to_unsigned(39,8) ,
68898	 => std_logic_vector(to_unsigned(51,8) ,
68899	 => std_logic_vector(to_unsigned(45,8) ,
68900	 => std_logic_vector(to_unsigned(36,8) ,
68901	 => std_logic_vector(to_unsigned(45,8) ,
68902	 => std_logic_vector(to_unsigned(38,8) ,
68903	 => std_logic_vector(to_unsigned(28,8) ,
68904	 => std_logic_vector(to_unsigned(22,8) ,
68905	 => std_logic_vector(to_unsigned(19,8) ,
68906	 => std_logic_vector(to_unsigned(16,8) ,
68907	 => std_logic_vector(to_unsigned(15,8) ,
68908	 => std_logic_vector(to_unsigned(14,8) ,
68909	 => std_logic_vector(to_unsigned(27,8) ,
68910	 => std_logic_vector(to_unsigned(60,8) ,
68911	 => std_logic_vector(to_unsigned(65,8) ,
68912	 => std_logic_vector(to_unsigned(41,8) ,
68913	 => std_logic_vector(to_unsigned(43,8) ,
68914	 => std_logic_vector(to_unsigned(50,8) ,
68915	 => std_logic_vector(to_unsigned(45,8) ,
68916	 => std_logic_vector(to_unsigned(96,8) ,
68917	 => std_logic_vector(to_unsigned(130,8) ,
68918	 => std_logic_vector(to_unsigned(74,8) ,
68919	 => std_logic_vector(to_unsigned(67,8) ,
68920	 => std_logic_vector(to_unsigned(92,8) ,
68921	 => std_logic_vector(to_unsigned(84,8) ,
68922	 => std_logic_vector(to_unsigned(90,8) ,
68923	 => std_logic_vector(to_unsigned(90,8) ,
68924	 => std_logic_vector(to_unsigned(78,8) ,
68925	 => std_logic_vector(to_unsigned(73,8) ,
68926	 => std_logic_vector(to_unsigned(63,8) ,
68927	 => std_logic_vector(to_unsigned(54,8) ,
68928	 => std_logic_vector(to_unsigned(56,8) ,
68929	 => std_logic_vector(to_unsigned(86,8) ,
68930	 => std_logic_vector(to_unsigned(111,8) ,
68931	 => std_logic_vector(to_unsigned(114,8) ,
68932	 => std_logic_vector(to_unsigned(118,8) ,
68933	 => std_logic_vector(to_unsigned(114,8) ,
68934	 => std_logic_vector(to_unsigned(105,8) ,
68935	 => std_logic_vector(to_unsigned(122,8) ,
68936	 => std_logic_vector(to_unsigned(86,8) ,
68937	 => std_logic_vector(to_unsigned(23,8) ,
68938	 => std_logic_vector(to_unsigned(32,8) ,
68939	 => std_logic_vector(to_unsigned(74,8) ,
68940	 => std_logic_vector(to_unsigned(81,8) ,
68941	 => std_logic_vector(to_unsigned(79,8) ,
68942	 => std_logic_vector(to_unsigned(73,8) ,
68943	 => std_logic_vector(to_unsigned(61,8) ,
68944	 => std_logic_vector(to_unsigned(51,8) ,
68945	 => std_logic_vector(to_unsigned(44,8) ,
68946	 => std_logic_vector(to_unsigned(51,8) ,
68947	 => std_logic_vector(to_unsigned(29,8) ,
68948	 => std_logic_vector(to_unsigned(16,8) ,
68949	 => std_logic_vector(to_unsigned(29,8) ,
68950	 => std_logic_vector(to_unsigned(27,8) ,
68951	 => std_logic_vector(to_unsigned(13,8) ,
68952	 => std_logic_vector(to_unsigned(36,8) ,
68953	 => std_logic_vector(to_unsigned(29,8) ,
68954	 => std_logic_vector(to_unsigned(23,8) ,
68955	 => std_logic_vector(to_unsigned(51,8) ,
68956	 => std_logic_vector(to_unsigned(40,8) ,
68957	 => std_logic_vector(to_unsigned(18,8) ,
68958	 => std_logic_vector(to_unsigned(22,8) ,
68959	 => std_logic_vector(to_unsigned(24,8) ,
68960	 => std_logic_vector(to_unsigned(27,8) ,
68961	 => std_logic_vector(to_unsigned(40,8) ,
68962	 => std_logic_vector(to_unsigned(16,8) ,
68963	 => std_logic_vector(to_unsigned(20,8) ,
68964	 => std_logic_vector(to_unsigned(33,8) ,
68965	 => std_logic_vector(to_unsigned(22,8) ,
68966	 => std_logic_vector(to_unsigned(6,8) ,
68967	 => std_logic_vector(to_unsigned(6,8) ,
68968	 => std_logic_vector(to_unsigned(13,8) ,
68969	 => std_logic_vector(to_unsigned(27,8) ,
68970	 => std_logic_vector(to_unsigned(24,8) ,
68971	 => std_logic_vector(to_unsigned(26,8) ,
68972	 => std_logic_vector(to_unsigned(20,8) ,
68973	 => std_logic_vector(to_unsigned(24,8) ,
68974	 => std_logic_vector(to_unsigned(56,8) ,
68975	 => std_logic_vector(to_unsigned(32,8) ,
68976	 => std_logic_vector(to_unsigned(29,8) ,
68977	 => std_logic_vector(to_unsigned(23,8) ,
68978	 => std_logic_vector(to_unsigned(22,8) ,
68979	 => std_logic_vector(to_unsigned(35,8) ,
68980	 => std_logic_vector(to_unsigned(24,8) ,
68981	 => std_logic_vector(to_unsigned(9,8) ,
68982	 => std_logic_vector(to_unsigned(11,8) ,
68983	 => std_logic_vector(to_unsigned(13,8) ,
68984	 => std_logic_vector(to_unsigned(10,8) ,
68985	 => std_logic_vector(to_unsigned(16,8) ,
68986	 => std_logic_vector(to_unsigned(37,8) ,
68987	 => std_logic_vector(to_unsigned(49,8) ,
68988	 => std_logic_vector(to_unsigned(54,8) ,
68989	 => std_logic_vector(to_unsigned(46,8) ,
68990	 => std_logic_vector(to_unsigned(36,8) ,
68991	 => std_logic_vector(to_unsigned(35,8) ,
68992	 => std_logic_vector(to_unsigned(37,8) ,
68993	 => std_logic_vector(to_unsigned(44,8) ,
68994	 => std_logic_vector(to_unsigned(35,8) ,
68995	 => std_logic_vector(to_unsigned(37,8) ,
68996	 => std_logic_vector(to_unsigned(38,8) ,
68997	 => std_logic_vector(to_unsigned(56,8) ,
68998	 => std_logic_vector(to_unsigned(70,8) ,
68999	 => std_logic_vector(to_unsigned(54,8) ,
69000	 => std_logic_vector(to_unsigned(39,8) ,
69001	 => std_logic_vector(to_unsigned(30,8) ,
69002	 => std_logic_vector(to_unsigned(17,8) ,
69003	 => std_logic_vector(to_unsigned(7,8) ,
69004	 => std_logic_vector(to_unsigned(14,8) ,
69005	 => std_logic_vector(to_unsigned(20,8) ,
69006	 => std_logic_vector(to_unsigned(12,8) ,
69007	 => std_logic_vector(to_unsigned(9,8) ,
69008	 => std_logic_vector(to_unsigned(20,8) ,
69009	 => std_logic_vector(to_unsigned(47,8) ,
69010	 => std_logic_vector(to_unsigned(80,8) ,
69011	 => std_logic_vector(to_unsigned(68,8) ,
69012	 => std_logic_vector(to_unsigned(32,8) ,
69013	 => std_logic_vector(to_unsigned(30,8) ,
69014	 => std_logic_vector(to_unsigned(32,8) ,
69015	 => std_logic_vector(to_unsigned(29,8) ,
69016	 => std_logic_vector(to_unsigned(24,8) ,
69017	 => std_logic_vector(to_unsigned(25,8) ,
69018	 => std_logic_vector(to_unsigned(23,8) ,
69019	 => std_logic_vector(to_unsigned(28,8) ,
69020	 => std_logic_vector(to_unsigned(55,8) ,
69021	 => std_logic_vector(to_unsigned(42,8) ,
69022	 => std_logic_vector(to_unsigned(30,8) ,
69023	 => std_logic_vector(to_unsigned(31,8) ,
69024	 => std_logic_vector(to_unsigned(40,8) ,
69025	 => std_logic_vector(to_unsigned(30,8) ,
69026	 => std_logic_vector(to_unsigned(31,8) ,
69027	 => std_logic_vector(to_unsigned(40,8) ,
69028	 => std_logic_vector(to_unsigned(26,8) ,
69029	 => std_logic_vector(to_unsigned(4,8) ,
69030	 => std_logic_vector(to_unsigned(13,8) ,
69031	 => std_logic_vector(to_unsigned(45,8) ,
69032	 => std_logic_vector(to_unsigned(29,8) ,
69033	 => std_logic_vector(to_unsigned(28,8) ,
69034	 => std_logic_vector(to_unsigned(39,8) ,
69035	 => std_logic_vector(to_unsigned(59,8) ,
69036	 => std_logic_vector(to_unsigned(30,8) ,
69037	 => std_logic_vector(to_unsigned(30,8) ,
69038	 => std_logic_vector(to_unsigned(60,8) ,
69039	 => std_logic_vector(to_unsigned(64,8) ,
69040	 => std_logic_vector(to_unsigned(49,8) ,
69041	 => std_logic_vector(to_unsigned(60,8) ,
69042	 => std_logic_vector(to_unsigned(45,8) ,
69043	 => std_logic_vector(to_unsigned(71,8) ,
69044	 => std_logic_vector(to_unsigned(108,8) ,
69045	 => std_logic_vector(to_unsigned(105,8) ,
69046	 => std_logic_vector(to_unsigned(51,8) ,
69047	 => std_logic_vector(to_unsigned(59,8) ,
69048	 => std_logic_vector(to_unsigned(118,8) ,
69049	 => std_logic_vector(to_unsigned(127,8) ,
69050	 => std_logic_vector(to_unsigned(51,8) ,
69051	 => std_logic_vector(to_unsigned(15,8) ,
69052	 => std_logic_vector(to_unsigned(39,8) ,
69053	 => std_logic_vector(to_unsigned(51,8) ,
69054	 => std_logic_vector(to_unsigned(35,8) ,
69055	 => std_logic_vector(to_unsigned(31,8) ,
69056	 => std_logic_vector(to_unsigned(32,8) ,
69057	 => std_logic_vector(to_unsigned(37,8) ,
69058	 => std_logic_vector(to_unsigned(41,8) ,
69059	 => std_logic_vector(to_unsigned(45,8) ,
69060	 => std_logic_vector(to_unsigned(45,8) ,
69061	 => std_logic_vector(to_unsigned(12,8) ,
69062	 => std_logic_vector(to_unsigned(9,8) ,
69063	 => std_logic_vector(to_unsigned(23,8) ,
69064	 => std_logic_vector(to_unsigned(33,8) ,
69065	 => std_logic_vector(to_unsigned(43,8) ,
69066	 => std_logic_vector(to_unsigned(44,8) ,
69067	 => std_logic_vector(to_unsigned(37,8) ,
69068	 => std_logic_vector(to_unsigned(33,8) ,
69069	 => std_logic_vector(to_unsigned(25,8) ,
69070	 => std_logic_vector(to_unsigned(24,8) ,
69071	 => std_logic_vector(to_unsigned(14,8) ,
69072	 => std_logic_vector(to_unsigned(8,8) ,
69073	 => std_logic_vector(to_unsigned(9,8) ,
69074	 => std_logic_vector(to_unsigned(2,8) ,
69075	 => std_logic_vector(to_unsigned(0,8) ,
69076	 => std_logic_vector(to_unsigned(2,8) ,
69077	 => std_logic_vector(to_unsigned(4,8) ,
69078	 => std_logic_vector(to_unsigned(9,8) ,
69079	 => std_logic_vector(to_unsigned(20,8) ,
69080	 => std_logic_vector(to_unsigned(9,8) ,
69081	 => std_logic_vector(to_unsigned(14,8) ,
69082	 => std_logic_vector(to_unsigned(10,8) ,
69083	 => std_logic_vector(to_unsigned(8,8) ,
69084	 => std_logic_vector(to_unsigned(5,8) ,
69085	 => std_logic_vector(to_unsigned(4,8) ,
69086	 => std_logic_vector(to_unsigned(1,8) ,
69087	 => std_logic_vector(to_unsigned(1,8) ,
69088	 => std_logic_vector(to_unsigned(10,8) ,
69089	 => std_logic_vector(to_unsigned(27,8) ,
69090	 => std_logic_vector(to_unsigned(30,8) ,
69091	 => std_logic_vector(to_unsigned(40,8) ,
69092	 => std_logic_vector(to_unsigned(43,8) ,
69093	 => std_logic_vector(to_unsigned(51,8) ,
69094	 => std_logic_vector(to_unsigned(53,8) ,
69095	 => std_logic_vector(to_unsigned(37,8) ,
69096	 => std_logic_vector(to_unsigned(58,8) ,
69097	 => std_logic_vector(to_unsigned(55,8) ,
69098	 => std_logic_vector(to_unsigned(72,8) ,
69099	 => std_logic_vector(to_unsigned(43,8) ,
69100	 => std_logic_vector(to_unsigned(26,8) ,
69101	 => std_logic_vector(to_unsigned(2,8) ,
69102	 => std_logic_vector(to_unsigned(0,8) ,
69103	 => std_logic_vector(to_unsigned(9,8) ,
69104	 => std_logic_vector(to_unsigned(62,8) ,
69105	 => std_logic_vector(to_unsigned(91,8) ,
69106	 => std_logic_vector(to_unsigned(35,8) ,
69107	 => std_logic_vector(to_unsigned(62,8) ,
69108	 => std_logic_vector(to_unsigned(28,8) ,
69109	 => std_logic_vector(to_unsigned(7,8) ,
69110	 => std_logic_vector(to_unsigned(10,8) ,
69111	 => std_logic_vector(to_unsigned(12,8) ,
69112	 => std_logic_vector(to_unsigned(12,8) ,
69113	 => std_logic_vector(to_unsigned(13,8) ,
69114	 => std_logic_vector(to_unsigned(10,8) ,
69115	 => std_logic_vector(to_unsigned(11,8) ,
69116	 => std_logic_vector(to_unsigned(17,8) ,
69117	 => std_logic_vector(to_unsigned(8,8) ,
69118	 => std_logic_vector(to_unsigned(9,8) ,
69119	 => std_logic_vector(to_unsigned(11,8) ,
69120	 => std_logic_vector(to_unsigned(8,8) ,
69121	 => std_logic_vector(to_unsigned(114,8) ,
69122	 => std_logic_vector(to_unsigned(125,8) ,
69123	 => std_logic_vector(to_unsigned(121,8) ,
69124	 => std_logic_vector(to_unsigned(109,8) ,
69125	 => std_logic_vector(to_unsigned(107,8) ,
69126	 => std_logic_vector(to_unsigned(118,8) ,
69127	 => std_logic_vector(to_unsigned(111,8) ,
69128	 => std_logic_vector(to_unsigned(86,8) ,
69129	 => std_logic_vector(to_unsigned(95,8) ,
69130	 => std_logic_vector(to_unsigned(116,8) ,
69131	 => std_logic_vector(to_unsigned(85,8) ,
69132	 => std_logic_vector(to_unsigned(48,8) ,
69133	 => std_logic_vector(to_unsigned(51,8) ,
69134	 => std_logic_vector(to_unsigned(46,8) ,
69135	 => std_logic_vector(to_unsigned(49,8) ,
69136	 => std_logic_vector(to_unsigned(53,8) ,
69137	 => std_logic_vector(to_unsigned(74,8) ,
69138	 => std_logic_vector(to_unsigned(70,8) ,
69139	 => std_logic_vector(to_unsigned(64,8) ,
69140	 => std_logic_vector(to_unsigned(74,8) ,
69141	 => std_logic_vector(to_unsigned(55,8) ,
69142	 => std_logic_vector(to_unsigned(41,8) ,
69143	 => std_logic_vector(to_unsigned(45,8) ,
69144	 => std_logic_vector(to_unsigned(41,8) ,
69145	 => std_logic_vector(to_unsigned(32,8) ,
69146	 => std_logic_vector(to_unsigned(34,8) ,
69147	 => std_logic_vector(to_unsigned(35,8) ,
69148	 => std_logic_vector(to_unsigned(41,8) ,
69149	 => std_logic_vector(to_unsigned(41,8) ,
69150	 => std_logic_vector(to_unsigned(44,8) ,
69151	 => std_logic_vector(to_unsigned(35,8) ,
69152	 => std_logic_vector(to_unsigned(35,8) ,
69153	 => std_logic_vector(to_unsigned(45,8) ,
69154	 => std_logic_vector(to_unsigned(62,8) ,
69155	 => std_logic_vector(to_unsigned(79,8) ,
69156	 => std_logic_vector(to_unsigned(79,8) ,
69157	 => std_logic_vector(to_unsigned(77,8) ,
69158	 => std_logic_vector(to_unsigned(80,8) ,
69159	 => std_logic_vector(to_unsigned(79,8) ,
69160	 => std_logic_vector(to_unsigned(68,8) ,
69161	 => std_logic_vector(to_unsigned(47,8) ,
69162	 => std_logic_vector(to_unsigned(35,8) ,
69163	 => std_logic_vector(to_unsigned(41,8) ,
69164	 => std_logic_vector(to_unsigned(52,8) ,
69165	 => std_logic_vector(to_unsigned(56,8) ,
69166	 => std_logic_vector(to_unsigned(54,8) ,
69167	 => std_logic_vector(to_unsigned(61,8) ,
69168	 => std_logic_vector(to_unsigned(51,8) ,
69169	 => std_logic_vector(to_unsigned(30,8) ,
69170	 => std_logic_vector(to_unsigned(24,8) ,
69171	 => std_logic_vector(to_unsigned(25,8) ,
69172	 => std_logic_vector(to_unsigned(23,8) ,
69173	 => std_logic_vector(to_unsigned(27,8) ,
69174	 => std_logic_vector(to_unsigned(37,8) ,
69175	 => std_logic_vector(to_unsigned(50,8) ,
69176	 => std_logic_vector(to_unsigned(56,8) ,
69177	 => std_logic_vector(to_unsigned(69,8) ,
69178	 => std_logic_vector(to_unsigned(53,8) ,
69179	 => std_logic_vector(to_unsigned(37,8) ,
69180	 => std_logic_vector(to_unsigned(41,8) ,
69181	 => std_logic_vector(to_unsigned(45,8) ,
69182	 => std_logic_vector(to_unsigned(37,8) ,
69183	 => std_logic_vector(to_unsigned(30,8) ,
69184	 => std_logic_vector(to_unsigned(46,8) ,
69185	 => std_logic_vector(to_unsigned(79,8) ,
69186	 => std_logic_vector(to_unsigned(85,8) ,
69187	 => std_logic_vector(to_unsigned(88,8) ,
69188	 => std_logic_vector(to_unsigned(104,8) ,
69189	 => std_logic_vector(to_unsigned(96,8) ,
69190	 => std_logic_vector(to_unsigned(101,8) ,
69191	 => std_logic_vector(to_unsigned(112,8) ,
69192	 => std_logic_vector(to_unsigned(124,8) ,
69193	 => std_logic_vector(to_unsigned(104,8) ,
69194	 => std_logic_vector(to_unsigned(90,8) ,
69195	 => std_logic_vector(to_unsigned(87,8) ,
69196	 => std_logic_vector(to_unsigned(45,8) ,
69197	 => std_logic_vector(to_unsigned(57,8) ,
69198	 => std_logic_vector(to_unsigned(104,8) ,
69199	 => std_logic_vector(to_unsigned(95,8) ,
69200	 => std_logic_vector(to_unsigned(97,8) ,
69201	 => std_logic_vector(to_unsigned(84,8) ,
69202	 => std_logic_vector(to_unsigned(59,8) ,
69203	 => std_logic_vector(to_unsigned(84,8) ,
69204	 => std_logic_vector(to_unsigned(84,8) ,
69205	 => std_logic_vector(to_unsigned(78,8) ,
69206	 => std_logic_vector(to_unsigned(72,8) ,
69207	 => std_logic_vector(to_unsigned(72,8) ,
69208	 => std_logic_vector(to_unsigned(70,8) ,
69209	 => std_logic_vector(to_unsigned(58,8) ,
69210	 => std_logic_vector(to_unsigned(36,8) ,
69211	 => std_logic_vector(to_unsigned(20,8) ,
69212	 => std_logic_vector(to_unsigned(29,8) ,
69213	 => std_logic_vector(to_unsigned(34,8) ,
69214	 => std_logic_vector(to_unsigned(32,8) ,
69215	 => std_logic_vector(to_unsigned(38,8) ,
69216	 => std_logic_vector(to_unsigned(45,8) ,
69217	 => std_logic_vector(to_unsigned(35,8) ,
69218	 => std_logic_vector(to_unsigned(50,8) ,
69219	 => std_logic_vector(to_unsigned(50,8) ,
69220	 => std_logic_vector(to_unsigned(45,8) ,
69221	 => std_logic_vector(to_unsigned(45,8) ,
69222	 => std_logic_vector(to_unsigned(35,8) ,
69223	 => std_logic_vector(to_unsigned(32,8) ,
69224	 => std_logic_vector(to_unsigned(24,8) ,
69225	 => std_logic_vector(to_unsigned(19,8) ,
69226	 => std_logic_vector(to_unsigned(14,8) ,
69227	 => std_logic_vector(to_unsigned(19,8) ,
69228	 => std_logic_vector(to_unsigned(19,8) ,
69229	 => std_logic_vector(to_unsigned(32,8) ,
69230	 => std_logic_vector(to_unsigned(43,8) ,
69231	 => std_logic_vector(to_unsigned(41,8) ,
69232	 => std_logic_vector(to_unsigned(43,8) ,
69233	 => std_logic_vector(to_unsigned(56,8) ,
69234	 => std_logic_vector(to_unsigned(74,8) ,
69235	 => std_logic_vector(to_unsigned(46,8) ,
69236	 => std_logic_vector(to_unsigned(80,8) ,
69237	 => std_logic_vector(to_unsigned(128,8) ,
69238	 => std_logic_vector(to_unsigned(108,8) ,
69239	 => std_logic_vector(to_unsigned(112,8) ,
69240	 => std_logic_vector(to_unsigned(118,8) ,
69241	 => std_logic_vector(to_unsigned(107,8) ,
69242	 => std_logic_vector(to_unsigned(104,8) ,
69243	 => std_logic_vector(to_unsigned(91,8) ,
69244	 => std_logic_vector(to_unsigned(81,8) ,
69245	 => std_logic_vector(to_unsigned(80,8) ,
69246	 => std_logic_vector(to_unsigned(76,8) ,
69247	 => std_logic_vector(to_unsigned(73,8) ,
69248	 => std_logic_vector(to_unsigned(78,8) ,
69249	 => std_logic_vector(to_unsigned(101,8) ,
69250	 => std_logic_vector(to_unsigned(109,8) ,
69251	 => std_logic_vector(to_unsigned(107,8) ,
69252	 => std_logic_vector(to_unsigned(112,8) ,
69253	 => std_logic_vector(to_unsigned(111,8) ,
69254	 => std_logic_vector(to_unsigned(115,8) ,
69255	 => std_logic_vector(to_unsigned(112,8) ,
69256	 => std_logic_vector(to_unsigned(87,8) ,
69257	 => std_logic_vector(to_unsigned(53,8) ,
69258	 => std_logic_vector(to_unsigned(51,8) ,
69259	 => std_logic_vector(to_unsigned(70,8) ,
69260	 => std_logic_vector(to_unsigned(72,8) ,
69261	 => std_logic_vector(to_unsigned(51,8) ,
69262	 => std_logic_vector(to_unsigned(77,8) ,
69263	 => std_logic_vector(to_unsigned(91,8) ,
69264	 => std_logic_vector(to_unsigned(61,8) ,
69265	 => std_logic_vector(to_unsigned(54,8) ,
69266	 => std_logic_vector(to_unsigned(25,8) ,
69267	 => std_logic_vector(to_unsigned(10,8) ,
69268	 => std_logic_vector(to_unsigned(20,8) ,
69269	 => std_logic_vector(to_unsigned(20,8) ,
69270	 => std_logic_vector(to_unsigned(22,8) ,
69271	 => std_logic_vector(to_unsigned(17,8) ,
69272	 => std_logic_vector(to_unsigned(27,8) ,
69273	 => std_logic_vector(to_unsigned(21,8) ,
69274	 => std_logic_vector(to_unsigned(16,8) ,
69275	 => std_logic_vector(to_unsigned(57,8) ,
69276	 => std_logic_vector(to_unsigned(47,8) ,
69277	 => std_logic_vector(to_unsigned(30,8) ,
69278	 => std_logic_vector(to_unsigned(21,8) ,
69279	 => std_logic_vector(to_unsigned(14,8) ,
69280	 => std_logic_vector(to_unsigned(16,8) ,
69281	 => std_logic_vector(to_unsigned(13,8) ,
69282	 => std_logic_vector(to_unsigned(8,8) ,
69283	 => std_logic_vector(to_unsigned(6,8) ,
69284	 => std_logic_vector(to_unsigned(13,8) ,
69285	 => std_logic_vector(to_unsigned(37,8) ,
69286	 => std_logic_vector(to_unsigned(12,8) ,
69287	 => std_logic_vector(to_unsigned(5,8) ,
69288	 => std_logic_vector(to_unsigned(7,8) ,
69289	 => std_logic_vector(to_unsigned(24,8) ,
69290	 => std_logic_vector(to_unsigned(27,8) ,
69291	 => std_logic_vector(to_unsigned(13,8) ,
69292	 => std_logic_vector(to_unsigned(22,8) ,
69293	 => std_logic_vector(to_unsigned(58,8) ,
69294	 => std_logic_vector(to_unsigned(22,8) ,
69295	 => std_logic_vector(to_unsigned(20,8) ,
69296	 => std_logic_vector(to_unsigned(30,8) ,
69297	 => std_logic_vector(to_unsigned(21,8) ,
69298	 => std_logic_vector(to_unsigned(28,8) ,
69299	 => std_logic_vector(to_unsigned(25,8) ,
69300	 => std_logic_vector(to_unsigned(32,8) ,
69301	 => std_logic_vector(to_unsigned(18,8) ,
69302	 => std_logic_vector(to_unsigned(11,8) ,
69303	 => std_logic_vector(to_unsigned(19,8) ,
69304	 => std_logic_vector(to_unsigned(14,8) ,
69305	 => std_logic_vector(to_unsigned(14,8) ,
69306	 => std_logic_vector(to_unsigned(30,8) ,
69307	 => std_logic_vector(to_unsigned(46,8) ,
69308	 => std_logic_vector(to_unsigned(48,8) ,
69309	 => std_logic_vector(to_unsigned(37,8) ,
69310	 => std_logic_vector(to_unsigned(32,8) ,
69311	 => std_logic_vector(to_unsigned(34,8) ,
69312	 => std_logic_vector(to_unsigned(41,8) ,
69313	 => std_logic_vector(to_unsigned(48,8) ,
69314	 => std_logic_vector(to_unsigned(45,8) ,
69315	 => std_logic_vector(to_unsigned(38,8) ,
69316	 => std_logic_vector(to_unsigned(37,8) ,
69317	 => std_logic_vector(to_unsigned(46,8) ,
69318	 => std_logic_vector(to_unsigned(68,8) ,
69319	 => std_logic_vector(to_unsigned(68,8) ,
69320	 => std_logic_vector(to_unsigned(37,8) ,
69321	 => std_logic_vector(to_unsigned(29,8) ,
69322	 => std_logic_vector(to_unsigned(17,8) ,
69323	 => std_logic_vector(to_unsigned(17,8) ,
69324	 => std_logic_vector(to_unsigned(17,8) ,
69325	 => std_logic_vector(to_unsigned(19,8) ,
69326	 => std_logic_vector(to_unsigned(13,8) ,
69327	 => std_logic_vector(to_unsigned(9,8) ,
69328	 => std_logic_vector(to_unsigned(25,8) ,
69329	 => std_logic_vector(to_unsigned(35,8) ,
69330	 => std_logic_vector(to_unsigned(35,8) ,
69331	 => std_logic_vector(to_unsigned(27,8) ,
69332	 => std_logic_vector(to_unsigned(29,8) ,
69333	 => std_logic_vector(to_unsigned(34,8) ,
69334	 => std_logic_vector(to_unsigned(39,8) ,
69335	 => std_logic_vector(to_unsigned(36,8) ,
69336	 => std_logic_vector(to_unsigned(25,8) ,
69337	 => std_logic_vector(to_unsigned(25,8) ,
69338	 => std_logic_vector(to_unsigned(27,8) ,
69339	 => std_logic_vector(to_unsigned(29,8) ,
69340	 => std_logic_vector(to_unsigned(26,8) ,
69341	 => std_logic_vector(to_unsigned(26,8) ,
69342	 => std_logic_vector(to_unsigned(24,8) ,
69343	 => std_logic_vector(to_unsigned(28,8) ,
69344	 => std_logic_vector(to_unsigned(45,8) ,
69345	 => std_logic_vector(to_unsigned(40,8) ,
69346	 => std_logic_vector(to_unsigned(29,8) ,
69347	 => std_logic_vector(to_unsigned(32,8) ,
69348	 => std_logic_vector(to_unsigned(24,8) ,
69349	 => std_logic_vector(to_unsigned(3,8) ,
69350	 => std_logic_vector(to_unsigned(15,8) ,
69351	 => std_logic_vector(to_unsigned(38,8) ,
69352	 => std_logic_vector(to_unsigned(17,8) ,
69353	 => std_logic_vector(to_unsigned(24,8) ,
69354	 => std_logic_vector(to_unsigned(37,8) ,
69355	 => std_logic_vector(to_unsigned(71,8) ,
69356	 => std_logic_vector(to_unsigned(16,8) ,
69357	 => std_logic_vector(to_unsigned(4,8) ,
69358	 => std_logic_vector(to_unsigned(48,8) ,
69359	 => std_logic_vector(to_unsigned(67,8) ,
69360	 => std_logic_vector(to_unsigned(50,8) ,
69361	 => std_logic_vector(to_unsigned(58,8) ,
69362	 => std_logic_vector(to_unsigned(46,8) ,
69363	 => std_logic_vector(to_unsigned(71,8) ,
69364	 => std_logic_vector(to_unsigned(97,8) ,
69365	 => std_logic_vector(to_unsigned(109,8) ,
69366	 => std_logic_vector(to_unsigned(49,8) ,
69367	 => std_logic_vector(to_unsigned(67,8) ,
69368	 => std_logic_vector(to_unsigned(127,8) ,
69369	 => std_logic_vector(to_unsigned(109,8) ,
69370	 => std_logic_vector(to_unsigned(45,8) ,
69371	 => std_logic_vector(to_unsigned(27,8) ,
69372	 => std_logic_vector(to_unsigned(39,8) ,
69373	 => std_logic_vector(to_unsigned(36,8) ,
69374	 => std_logic_vector(to_unsigned(28,8) ,
69375	 => std_logic_vector(to_unsigned(14,8) ,
69376	 => std_logic_vector(to_unsigned(20,8) ,
69377	 => std_logic_vector(to_unsigned(47,8) ,
69378	 => std_logic_vector(to_unsigned(35,8) ,
69379	 => std_logic_vector(to_unsigned(26,8) ,
69380	 => std_logic_vector(to_unsigned(27,8) ,
69381	 => std_logic_vector(to_unsigned(18,8) ,
69382	 => std_logic_vector(to_unsigned(10,8) ,
69383	 => std_logic_vector(to_unsigned(7,8) ,
69384	 => std_logic_vector(to_unsigned(11,8) ,
69385	 => std_logic_vector(to_unsigned(9,8) ,
69386	 => std_logic_vector(to_unsigned(13,8) ,
69387	 => std_logic_vector(to_unsigned(16,8) ,
69388	 => std_logic_vector(to_unsigned(36,8) ,
69389	 => std_logic_vector(to_unsigned(45,8) ,
69390	 => std_logic_vector(to_unsigned(37,8) ,
69391	 => std_logic_vector(to_unsigned(29,8) ,
69392	 => std_logic_vector(to_unsigned(13,8) ,
69393	 => std_logic_vector(to_unsigned(14,8) ,
69394	 => std_logic_vector(to_unsigned(8,8) ,
69395	 => std_logic_vector(to_unsigned(0,8) ,
69396	 => std_logic_vector(to_unsigned(1,8) ,
69397	 => std_logic_vector(to_unsigned(10,8) ,
69398	 => std_logic_vector(to_unsigned(15,8) ,
69399	 => std_logic_vector(to_unsigned(13,8) ,
69400	 => std_logic_vector(to_unsigned(9,8) ,
69401	 => std_logic_vector(to_unsigned(11,8) ,
69402	 => std_logic_vector(to_unsigned(16,8) ,
69403	 => std_logic_vector(to_unsigned(13,8) ,
69404	 => std_logic_vector(to_unsigned(3,8) ,
69405	 => std_logic_vector(to_unsigned(6,8) ,
69406	 => std_logic_vector(to_unsigned(1,8) ,
69407	 => std_logic_vector(to_unsigned(0,8) ,
69408	 => std_logic_vector(to_unsigned(6,8) ,
69409	 => std_logic_vector(to_unsigned(25,8) ,
69410	 => std_logic_vector(to_unsigned(27,8) ,
69411	 => std_logic_vector(to_unsigned(19,8) ,
69412	 => std_logic_vector(to_unsigned(13,8) ,
69413	 => std_logic_vector(to_unsigned(11,8) ,
69414	 => std_logic_vector(to_unsigned(14,8) ,
69415	 => std_logic_vector(to_unsigned(20,8) ,
69416	 => std_logic_vector(to_unsigned(24,8) ,
69417	 => std_logic_vector(to_unsigned(27,8) ,
69418	 => std_logic_vector(to_unsigned(40,8) ,
69419	 => std_logic_vector(to_unsigned(64,8) ,
69420	 => std_logic_vector(to_unsigned(74,8) ,
69421	 => std_logic_vector(to_unsigned(6,8) ,
69422	 => std_logic_vector(to_unsigned(0,8) ,
69423	 => std_logic_vector(to_unsigned(5,8) ,
69424	 => std_logic_vector(to_unsigned(60,8) ,
69425	 => std_logic_vector(to_unsigned(92,8) ,
69426	 => std_logic_vector(to_unsigned(20,8) ,
69427	 => std_logic_vector(to_unsigned(54,8) ,
69428	 => std_logic_vector(to_unsigned(30,8) ,
69429	 => std_logic_vector(to_unsigned(8,8) ,
69430	 => std_logic_vector(to_unsigned(14,8) ,
69431	 => std_logic_vector(to_unsigned(12,8) ,
69432	 => std_logic_vector(to_unsigned(11,8) ,
69433	 => std_logic_vector(to_unsigned(13,8) ,
69434	 => std_logic_vector(to_unsigned(11,8) ,
69435	 => std_logic_vector(to_unsigned(9,8) ,
69436	 => std_logic_vector(to_unsigned(8,8) ,
69437	 => std_logic_vector(to_unsigned(7,8) ,
69438	 => std_logic_vector(to_unsigned(9,8) ,
69439	 => std_logic_vector(to_unsigned(13,8) ,
69440	 => std_logic_vector(to_unsigned(13,8) ,
69441	 => std_logic_vector(to_unsigned(70,8) ,
69442	 => std_logic_vector(to_unsigned(104,8) ,
69443	 => std_logic_vector(to_unsigned(116,8) ,
69444	 => std_logic_vector(to_unsigned(88,8) ,
69445	 => std_logic_vector(to_unsigned(108,8) ,
69446	 => std_logic_vector(to_unsigned(116,8) ,
69447	 => std_logic_vector(to_unsigned(118,8) ,
69448	 => std_logic_vector(to_unsigned(97,8) ,
69449	 => std_logic_vector(to_unsigned(87,8) ,
69450	 => std_logic_vector(to_unsigned(74,8) ,
69451	 => std_logic_vector(to_unsigned(76,8) ,
69452	 => std_logic_vector(to_unsigned(60,8) ,
69453	 => std_logic_vector(to_unsigned(47,8) ,
69454	 => std_logic_vector(to_unsigned(43,8) ,
69455	 => std_logic_vector(to_unsigned(31,8) ,
69456	 => std_logic_vector(to_unsigned(39,8) ,
69457	 => std_logic_vector(to_unsigned(76,8) ,
69458	 => std_logic_vector(to_unsigned(56,8) ,
69459	 => std_logic_vector(to_unsigned(45,8) ,
69460	 => std_logic_vector(to_unsigned(52,8) ,
69461	 => std_logic_vector(to_unsigned(51,8) ,
69462	 => std_logic_vector(to_unsigned(46,8) ,
69463	 => std_logic_vector(to_unsigned(47,8) ,
69464	 => std_logic_vector(to_unsigned(60,8) ,
69465	 => std_logic_vector(to_unsigned(38,8) ,
69466	 => std_logic_vector(to_unsigned(37,8) ,
69467	 => std_logic_vector(to_unsigned(48,8) ,
69468	 => std_logic_vector(to_unsigned(45,8) ,
69469	 => std_logic_vector(to_unsigned(37,8) ,
69470	 => std_logic_vector(to_unsigned(34,8) ,
69471	 => std_logic_vector(to_unsigned(27,8) ,
69472	 => std_logic_vector(to_unsigned(37,8) ,
69473	 => std_logic_vector(to_unsigned(73,8) ,
69474	 => std_logic_vector(to_unsigned(93,8) ,
69475	 => std_logic_vector(to_unsigned(87,8) ,
69476	 => std_logic_vector(to_unsigned(77,8) ,
69477	 => std_logic_vector(to_unsigned(70,8) ,
69478	 => std_logic_vector(to_unsigned(77,8) ,
69479	 => std_logic_vector(to_unsigned(60,8) ,
69480	 => std_logic_vector(to_unsigned(29,8) ,
69481	 => std_logic_vector(to_unsigned(28,8) ,
69482	 => std_logic_vector(to_unsigned(43,8) ,
69483	 => std_logic_vector(to_unsigned(60,8) ,
69484	 => std_logic_vector(to_unsigned(59,8) ,
69485	 => std_logic_vector(to_unsigned(53,8) ,
69486	 => std_logic_vector(to_unsigned(51,8) ,
69487	 => std_logic_vector(to_unsigned(39,8) ,
69488	 => std_logic_vector(to_unsigned(23,8) ,
69489	 => std_logic_vector(to_unsigned(23,8) ,
69490	 => std_logic_vector(to_unsigned(27,8) ,
69491	 => std_logic_vector(to_unsigned(28,8) ,
69492	 => std_logic_vector(to_unsigned(30,8) ,
69493	 => std_logic_vector(to_unsigned(30,8) ,
69494	 => std_logic_vector(to_unsigned(32,8) ,
69495	 => std_logic_vector(to_unsigned(45,8) ,
69496	 => std_logic_vector(to_unsigned(41,8) ,
69497	 => std_logic_vector(to_unsigned(40,8) ,
69498	 => std_logic_vector(to_unsigned(41,8) ,
69499	 => std_logic_vector(to_unsigned(38,8) ,
69500	 => std_logic_vector(to_unsigned(41,8) ,
69501	 => std_logic_vector(to_unsigned(40,8) ,
69502	 => std_logic_vector(to_unsigned(37,8) ,
69503	 => std_logic_vector(to_unsigned(47,8) ,
69504	 => std_logic_vector(to_unsigned(76,8) ,
69505	 => std_logic_vector(to_unsigned(90,8) ,
69506	 => std_logic_vector(to_unsigned(104,8) ,
69507	 => std_logic_vector(to_unsigned(99,8) ,
69508	 => std_logic_vector(to_unsigned(77,8) ,
69509	 => std_logic_vector(to_unsigned(57,8) ,
69510	 => std_logic_vector(to_unsigned(86,8) ,
69511	 => std_logic_vector(to_unsigned(118,8) ,
69512	 => std_logic_vector(to_unsigned(108,8) ,
69513	 => std_logic_vector(to_unsigned(109,8) ,
69514	 => std_logic_vector(to_unsigned(114,8) ,
69515	 => std_logic_vector(to_unsigned(86,8) ,
69516	 => std_logic_vector(to_unsigned(56,8) ,
69517	 => std_logic_vector(to_unsigned(60,8) ,
69518	 => std_logic_vector(to_unsigned(78,8) ,
69519	 => std_logic_vector(to_unsigned(84,8) ,
69520	 => std_logic_vector(to_unsigned(85,8) ,
69521	 => std_logic_vector(to_unsigned(101,8) ,
69522	 => std_logic_vector(to_unsigned(90,8) ,
69523	 => std_logic_vector(to_unsigned(87,8) ,
69524	 => std_logic_vector(to_unsigned(86,8) ,
69525	 => std_logic_vector(to_unsigned(82,8) ,
69526	 => std_logic_vector(to_unsigned(76,8) ,
69527	 => std_logic_vector(to_unsigned(69,8) ,
69528	 => std_logic_vector(to_unsigned(68,8) ,
69529	 => std_logic_vector(to_unsigned(52,8) ,
69530	 => std_logic_vector(to_unsigned(28,8) ,
69531	 => std_logic_vector(to_unsigned(14,8) ,
69532	 => std_logic_vector(to_unsigned(28,8) ,
69533	 => std_logic_vector(to_unsigned(32,8) ,
69534	 => std_logic_vector(to_unsigned(27,8) ,
69535	 => std_logic_vector(to_unsigned(35,8) ,
69536	 => std_logic_vector(to_unsigned(34,8) ,
69537	 => std_logic_vector(to_unsigned(33,8) ,
69538	 => std_logic_vector(to_unsigned(34,8) ,
69539	 => std_logic_vector(to_unsigned(33,8) ,
69540	 => std_logic_vector(to_unsigned(35,8) ,
69541	 => std_logic_vector(to_unsigned(38,8) ,
69542	 => std_logic_vector(to_unsigned(39,8) ,
69543	 => std_logic_vector(to_unsigned(27,8) ,
69544	 => std_logic_vector(to_unsigned(19,8) ,
69545	 => std_logic_vector(to_unsigned(17,8) ,
69546	 => std_logic_vector(to_unsigned(23,8) ,
69547	 => std_logic_vector(to_unsigned(28,8) ,
69548	 => std_logic_vector(to_unsigned(16,8) ,
69549	 => std_logic_vector(to_unsigned(24,8) ,
69550	 => std_logic_vector(to_unsigned(46,8) ,
69551	 => std_logic_vector(to_unsigned(43,8) ,
69552	 => std_logic_vector(to_unsigned(36,8) ,
69553	 => std_logic_vector(to_unsigned(33,8) ,
69554	 => std_logic_vector(to_unsigned(27,8) ,
69555	 => std_logic_vector(to_unsigned(50,8) ,
69556	 => std_logic_vector(to_unsigned(96,8) ,
69557	 => std_logic_vector(to_unsigned(116,8) ,
69558	 => std_logic_vector(to_unsigned(116,8) ,
69559	 => std_logic_vector(to_unsigned(133,8) ,
69560	 => std_logic_vector(to_unsigned(130,8) ,
69561	 => std_logic_vector(to_unsigned(134,8) ,
69562	 => std_logic_vector(to_unsigned(133,8) ,
69563	 => std_logic_vector(to_unsigned(116,8) ,
69564	 => std_logic_vector(to_unsigned(112,8) ,
69565	 => std_logic_vector(to_unsigned(104,8) ,
69566	 => std_logic_vector(to_unsigned(93,8) ,
69567	 => std_logic_vector(to_unsigned(84,8) ,
69568	 => std_logic_vector(to_unsigned(93,8) ,
69569	 => std_logic_vector(to_unsigned(107,8) ,
69570	 => std_logic_vector(to_unsigned(95,8) ,
69571	 => std_logic_vector(to_unsigned(96,8) ,
69572	 => std_logic_vector(to_unsigned(109,8) ,
69573	 => std_logic_vector(to_unsigned(88,8) ,
69574	 => std_logic_vector(to_unsigned(84,8) ,
69575	 => std_logic_vector(to_unsigned(86,8) ,
69576	 => std_logic_vector(to_unsigned(70,8) ,
69577	 => std_logic_vector(to_unsigned(55,8) ,
69578	 => std_logic_vector(to_unsigned(54,8) ,
69579	 => std_logic_vector(to_unsigned(29,8) ,
69580	 => std_logic_vector(to_unsigned(25,8) ,
69581	 => std_logic_vector(to_unsigned(49,8) ,
69582	 => std_logic_vector(to_unsigned(92,8) ,
69583	 => std_logic_vector(to_unsigned(85,8) ,
69584	 => std_logic_vector(to_unsigned(37,8) ,
69585	 => std_logic_vector(to_unsigned(38,8) ,
69586	 => std_logic_vector(to_unsigned(26,8) ,
69587	 => std_logic_vector(to_unsigned(8,8) ,
69588	 => std_logic_vector(to_unsigned(9,8) ,
69589	 => std_logic_vector(to_unsigned(12,8) ,
69590	 => std_logic_vector(to_unsigned(15,8) ,
69591	 => std_logic_vector(to_unsigned(16,8) ,
69592	 => std_logic_vector(to_unsigned(24,8) ,
69593	 => std_logic_vector(to_unsigned(29,8) ,
69594	 => std_logic_vector(to_unsigned(24,8) ,
69595	 => std_logic_vector(to_unsigned(29,8) ,
69596	 => std_logic_vector(to_unsigned(20,8) ,
69597	 => std_logic_vector(to_unsigned(8,8) ,
69598	 => std_logic_vector(to_unsigned(5,8) ,
69599	 => std_logic_vector(to_unsigned(4,8) ,
69600	 => std_logic_vector(to_unsigned(6,8) ,
69601	 => std_logic_vector(to_unsigned(7,8) ,
69602	 => std_logic_vector(to_unsigned(12,8) ,
69603	 => std_logic_vector(to_unsigned(8,8) ,
69604	 => std_logic_vector(to_unsigned(28,8) ,
69605	 => std_logic_vector(to_unsigned(58,8) ,
69606	 => std_logic_vector(to_unsigned(26,8) ,
69607	 => std_logic_vector(to_unsigned(7,8) ,
69608	 => std_logic_vector(to_unsigned(7,8) ,
69609	 => std_logic_vector(to_unsigned(22,8) ,
69610	 => std_logic_vector(to_unsigned(20,8) ,
69611	 => std_logic_vector(to_unsigned(22,8) ,
69612	 => std_logic_vector(to_unsigned(46,8) ,
69613	 => std_logic_vector(to_unsigned(23,8) ,
69614	 => std_logic_vector(to_unsigned(22,8) ,
69615	 => std_logic_vector(to_unsigned(25,8) ,
69616	 => std_logic_vector(to_unsigned(17,8) ,
69617	 => std_logic_vector(to_unsigned(32,8) ,
69618	 => std_logic_vector(to_unsigned(22,8) ,
69619	 => std_logic_vector(to_unsigned(25,8) ,
69620	 => std_logic_vector(to_unsigned(61,8) ,
69621	 => std_logic_vector(to_unsigned(20,8) ,
69622	 => std_logic_vector(to_unsigned(12,8) ,
69623	 => std_logic_vector(to_unsigned(20,8) ,
69624	 => std_logic_vector(to_unsigned(11,8) ,
69625	 => std_logic_vector(to_unsigned(10,8) ,
69626	 => std_logic_vector(to_unsigned(28,8) ,
69627	 => std_logic_vector(to_unsigned(45,8) ,
69628	 => std_logic_vector(to_unsigned(45,8) ,
69629	 => std_logic_vector(to_unsigned(41,8) ,
69630	 => std_logic_vector(to_unsigned(35,8) ,
69631	 => std_logic_vector(to_unsigned(37,8) ,
69632	 => std_logic_vector(to_unsigned(42,8) ,
69633	 => std_logic_vector(to_unsigned(40,8) ,
69634	 => std_logic_vector(to_unsigned(37,8) ,
69635	 => std_logic_vector(to_unsigned(36,8) ,
69636	 => std_logic_vector(to_unsigned(36,8) ,
69637	 => std_logic_vector(to_unsigned(37,8) ,
69638	 => std_logic_vector(to_unsigned(47,8) ,
69639	 => std_logic_vector(to_unsigned(45,8) ,
69640	 => std_logic_vector(to_unsigned(35,8) ,
69641	 => std_logic_vector(to_unsigned(19,8) ,
69642	 => std_logic_vector(to_unsigned(17,8) ,
69643	 => std_logic_vector(to_unsigned(28,8) ,
69644	 => std_logic_vector(to_unsigned(12,8) ,
69645	 => std_logic_vector(to_unsigned(16,8) ,
69646	 => std_logic_vector(to_unsigned(10,8) ,
69647	 => std_logic_vector(to_unsigned(12,8) ,
69648	 => std_logic_vector(to_unsigned(25,8) ,
69649	 => std_logic_vector(to_unsigned(56,8) ,
69650	 => std_logic_vector(to_unsigned(52,8) ,
69651	 => std_logic_vector(to_unsigned(16,8) ,
69652	 => std_logic_vector(to_unsigned(27,8) ,
69653	 => std_logic_vector(to_unsigned(34,8) ,
69654	 => std_logic_vector(to_unsigned(33,8) ,
69655	 => std_logic_vector(to_unsigned(40,8) ,
69656	 => std_logic_vector(to_unsigned(41,8) ,
69657	 => std_logic_vector(to_unsigned(26,8) ,
69658	 => std_logic_vector(to_unsigned(24,8) ,
69659	 => std_logic_vector(to_unsigned(29,8) ,
69660	 => std_logic_vector(to_unsigned(35,8) ,
69661	 => std_logic_vector(to_unsigned(37,8) ,
69662	 => std_logic_vector(to_unsigned(23,8) ,
69663	 => std_logic_vector(to_unsigned(24,8) ,
69664	 => std_logic_vector(to_unsigned(36,8) ,
69665	 => std_logic_vector(to_unsigned(37,8) ,
69666	 => std_logic_vector(to_unsigned(41,8) ,
69667	 => std_logic_vector(to_unsigned(27,8) ,
69668	 => std_logic_vector(to_unsigned(18,8) ,
69669	 => std_logic_vector(to_unsigned(4,8) ,
69670	 => std_logic_vector(to_unsigned(15,8) ,
69671	 => std_logic_vector(to_unsigned(46,8) ,
69672	 => std_logic_vector(to_unsigned(35,8) ,
69673	 => std_logic_vector(to_unsigned(34,8) ,
69674	 => std_logic_vector(to_unsigned(37,8) ,
69675	 => std_logic_vector(to_unsigned(62,8) ,
69676	 => std_logic_vector(to_unsigned(29,8) ,
69677	 => std_logic_vector(to_unsigned(22,8) ,
69678	 => std_logic_vector(to_unsigned(57,8) ,
69679	 => std_logic_vector(to_unsigned(68,8) ,
69680	 => std_logic_vector(to_unsigned(42,8) ,
69681	 => std_logic_vector(to_unsigned(29,8) ,
69682	 => std_logic_vector(to_unsigned(37,8) ,
69683	 => std_logic_vector(to_unsigned(76,8) ,
69684	 => std_logic_vector(to_unsigned(95,8) ,
69685	 => std_logic_vector(to_unsigned(99,8) ,
69686	 => std_logic_vector(to_unsigned(45,8) ,
69687	 => std_logic_vector(to_unsigned(70,8) ,
69688	 => std_logic_vector(to_unsigned(130,8) ,
69689	 => std_logic_vector(to_unsigned(100,8) ,
69690	 => std_logic_vector(to_unsigned(38,8) ,
69691	 => std_logic_vector(to_unsigned(27,8) ,
69692	 => std_logic_vector(to_unsigned(38,8) ,
69693	 => std_logic_vector(to_unsigned(37,8) ,
69694	 => std_logic_vector(to_unsigned(32,8) ,
69695	 => std_logic_vector(to_unsigned(23,8) ,
69696	 => std_logic_vector(to_unsigned(35,8) ,
69697	 => std_logic_vector(to_unsigned(43,8) ,
69698	 => std_logic_vector(to_unsigned(44,8) ,
69699	 => std_logic_vector(to_unsigned(26,8) ,
69700	 => std_logic_vector(to_unsigned(20,8) ,
69701	 => std_logic_vector(to_unsigned(32,8) ,
69702	 => std_logic_vector(to_unsigned(32,8) ,
69703	 => std_logic_vector(to_unsigned(40,8) ,
69704	 => std_logic_vector(to_unsigned(32,8) ,
69705	 => std_logic_vector(to_unsigned(8,8) ,
69706	 => std_logic_vector(to_unsigned(3,8) ,
69707	 => std_logic_vector(to_unsigned(8,8) ,
69708	 => std_logic_vector(to_unsigned(37,8) ,
69709	 => std_logic_vector(to_unsigned(28,8) ,
69710	 => std_logic_vector(to_unsigned(22,8) ,
69711	 => std_logic_vector(to_unsigned(26,8) ,
69712	 => std_logic_vector(to_unsigned(12,8) ,
69713	 => std_logic_vector(to_unsigned(17,8) ,
69714	 => std_logic_vector(to_unsigned(18,8) ,
69715	 => std_logic_vector(to_unsigned(0,8) ,
69716	 => std_logic_vector(to_unsigned(0,8) ,
69717	 => std_logic_vector(to_unsigned(16,8) ,
69718	 => std_logic_vector(to_unsigned(49,8) ,
69719	 => std_logic_vector(to_unsigned(43,8) ,
69720	 => std_logic_vector(to_unsigned(47,8) ,
69721	 => std_logic_vector(to_unsigned(25,8) ,
69722	 => std_logic_vector(to_unsigned(10,8) ,
69723	 => std_logic_vector(to_unsigned(7,8) ,
69724	 => std_logic_vector(to_unsigned(4,8) ,
69725	 => std_logic_vector(to_unsigned(8,8) ,
69726	 => std_logic_vector(to_unsigned(1,8) ,
69727	 => std_logic_vector(to_unsigned(0,8) ,
69728	 => std_logic_vector(to_unsigned(3,8) ,
69729	 => std_logic_vector(to_unsigned(44,8) ,
69730	 => std_logic_vector(to_unsigned(76,8) ,
69731	 => std_logic_vector(to_unsigned(11,8) ,
69732	 => std_logic_vector(to_unsigned(3,8) ,
69733	 => std_logic_vector(to_unsigned(1,8) ,
69734	 => std_logic_vector(to_unsigned(1,8) ,
69735	 => std_logic_vector(to_unsigned(1,8) ,
69736	 => std_logic_vector(to_unsigned(1,8) ,
69737	 => std_logic_vector(to_unsigned(1,8) ,
69738	 => std_logic_vector(to_unsigned(3,8) ,
69739	 => std_logic_vector(to_unsigned(6,8) ,
69740	 => std_logic_vector(to_unsigned(23,8) ,
69741	 => std_logic_vector(to_unsigned(13,8) ,
69742	 => std_logic_vector(to_unsigned(0,8) ,
69743	 => std_logic_vector(to_unsigned(1,8) ,
69744	 => std_logic_vector(to_unsigned(39,8) ,
69745	 => std_logic_vector(to_unsigned(99,8) ,
69746	 => std_logic_vector(to_unsigned(22,8) ,
69747	 => std_logic_vector(to_unsigned(26,8) ,
69748	 => std_logic_vector(to_unsigned(24,8) ,
69749	 => std_logic_vector(to_unsigned(10,8) ,
69750	 => std_logic_vector(to_unsigned(16,8) ,
69751	 => std_logic_vector(to_unsigned(15,8) ,
69752	 => std_logic_vector(to_unsigned(13,8) ,
69753	 => std_logic_vector(to_unsigned(14,8) ,
69754	 => std_logic_vector(to_unsigned(8,8) ,
69755	 => std_logic_vector(to_unsigned(7,8) ,
69756	 => std_logic_vector(to_unsigned(9,8) ,
69757	 => std_logic_vector(to_unsigned(9,8) ,
69758	 => std_logic_vector(to_unsigned(12,8) ,
69759	 => std_logic_vector(to_unsigned(12,8) ,
69760	 => std_logic_vector(to_unsigned(11,8) ,
69761	 => std_logic_vector(to_unsigned(54,8) ,
69762	 => std_logic_vector(to_unsigned(99,8) ,
69763	 => std_logic_vector(to_unsigned(119,8) ,
69764	 => std_logic_vector(to_unsigned(69,8) ,
69765	 => std_logic_vector(to_unsigned(86,8) ,
69766	 => std_logic_vector(to_unsigned(87,8) ,
69767	 => std_logic_vector(to_unsigned(97,8) ,
69768	 => std_logic_vector(to_unsigned(88,8) ,
69769	 => std_logic_vector(to_unsigned(87,8) ,
69770	 => std_logic_vector(to_unsigned(77,8) ,
69771	 => std_logic_vector(to_unsigned(80,8) ,
69772	 => std_logic_vector(to_unsigned(76,8) ,
69773	 => std_logic_vector(to_unsigned(51,8) ,
69774	 => std_logic_vector(to_unsigned(52,8) ,
69775	 => std_logic_vector(to_unsigned(45,8) ,
69776	 => std_logic_vector(to_unsigned(50,8) ,
69777	 => std_logic_vector(to_unsigned(73,8) ,
69778	 => std_logic_vector(to_unsigned(63,8) ,
69779	 => std_logic_vector(to_unsigned(38,8) ,
69780	 => std_logic_vector(to_unsigned(39,8) ,
69781	 => std_logic_vector(to_unsigned(45,8) ,
69782	 => std_logic_vector(to_unsigned(53,8) ,
69783	 => std_logic_vector(to_unsigned(51,8) ,
69784	 => std_logic_vector(to_unsigned(100,8) ,
69785	 => std_logic_vector(to_unsigned(82,8) ,
69786	 => std_logic_vector(to_unsigned(48,8) ,
69787	 => std_logic_vector(to_unsigned(39,8) ,
69788	 => std_logic_vector(to_unsigned(32,8) ,
69789	 => std_logic_vector(to_unsigned(27,8) ,
69790	 => std_logic_vector(to_unsigned(37,8) ,
69791	 => std_logic_vector(to_unsigned(41,8) ,
69792	 => std_logic_vector(to_unsigned(46,8) ,
69793	 => std_logic_vector(to_unsigned(41,8) ,
69794	 => std_logic_vector(to_unsigned(33,8) ,
69795	 => std_logic_vector(to_unsigned(49,8) ,
69796	 => std_logic_vector(to_unsigned(62,8) ,
69797	 => std_logic_vector(to_unsigned(70,8) ,
69798	 => std_logic_vector(to_unsigned(41,8) ,
69799	 => std_logic_vector(to_unsigned(26,8) ,
69800	 => std_logic_vector(to_unsigned(35,8) ,
69801	 => std_logic_vector(to_unsigned(50,8) ,
69802	 => std_logic_vector(to_unsigned(61,8) ,
69803	 => std_logic_vector(to_unsigned(60,8) ,
69804	 => std_logic_vector(to_unsigned(45,8) ,
69805	 => std_logic_vector(to_unsigned(28,8) ,
69806	 => std_logic_vector(to_unsigned(29,8) ,
69807	 => std_logic_vector(to_unsigned(19,8) ,
69808	 => std_logic_vector(to_unsigned(16,8) ,
69809	 => std_logic_vector(to_unsigned(27,8) ,
69810	 => std_logic_vector(to_unsigned(30,8) ,
69811	 => std_logic_vector(to_unsigned(31,8) ,
69812	 => std_logic_vector(to_unsigned(37,8) ,
69813	 => std_logic_vector(to_unsigned(38,8) ,
69814	 => std_logic_vector(to_unsigned(38,8) ,
69815	 => std_logic_vector(to_unsigned(46,8) ,
69816	 => std_logic_vector(to_unsigned(41,8) ,
69817	 => std_logic_vector(to_unsigned(41,8) ,
69818	 => std_logic_vector(to_unsigned(39,8) ,
69819	 => std_logic_vector(to_unsigned(34,8) ,
69820	 => std_logic_vector(to_unsigned(44,8) ,
69821	 => std_logic_vector(to_unsigned(48,8) ,
69822	 => std_logic_vector(to_unsigned(42,8) ,
69823	 => std_logic_vector(to_unsigned(46,8) ,
69824	 => std_logic_vector(to_unsigned(52,8) ,
69825	 => std_logic_vector(to_unsigned(54,8) ,
69826	 => std_logic_vector(to_unsigned(64,8) ,
69827	 => std_logic_vector(to_unsigned(71,8) ,
69828	 => std_logic_vector(to_unsigned(58,8) ,
69829	 => std_logic_vector(to_unsigned(41,8) ,
69830	 => std_logic_vector(to_unsigned(54,8) ,
69831	 => std_logic_vector(to_unsigned(79,8) ,
69832	 => std_logic_vector(to_unsigned(53,8) ,
69833	 => std_logic_vector(to_unsigned(66,8) ,
69834	 => std_logic_vector(to_unsigned(78,8) ,
69835	 => std_logic_vector(to_unsigned(60,8) ,
69836	 => std_logic_vector(to_unsigned(52,8) ,
69837	 => std_logic_vector(to_unsigned(59,8) ,
69838	 => std_logic_vector(to_unsigned(60,8) ,
69839	 => std_logic_vector(to_unsigned(60,8) ,
69840	 => std_logic_vector(to_unsigned(54,8) ,
69841	 => std_logic_vector(to_unsigned(70,8) ,
69842	 => std_logic_vector(to_unsigned(62,8) ,
69843	 => std_logic_vector(to_unsigned(93,8) ,
69844	 => std_logic_vector(to_unsigned(88,8) ,
69845	 => std_logic_vector(to_unsigned(84,8) ,
69846	 => std_logic_vector(to_unsigned(78,8) ,
69847	 => std_logic_vector(to_unsigned(67,8) ,
69848	 => std_logic_vector(to_unsigned(59,8) ,
69849	 => std_logic_vector(to_unsigned(51,8) ,
69850	 => std_logic_vector(to_unsigned(26,8) ,
69851	 => std_logic_vector(to_unsigned(16,8) ,
69852	 => std_logic_vector(to_unsigned(32,8) ,
69853	 => std_logic_vector(to_unsigned(36,8) ,
69854	 => std_logic_vector(to_unsigned(34,8) ,
69855	 => std_logic_vector(to_unsigned(34,8) ,
69856	 => std_logic_vector(to_unsigned(32,8) ,
69857	 => std_logic_vector(to_unsigned(32,8) ,
69858	 => std_logic_vector(to_unsigned(34,8) ,
69859	 => std_logic_vector(to_unsigned(32,8) ,
69860	 => std_logic_vector(to_unsigned(27,8) ,
69861	 => std_logic_vector(to_unsigned(31,8) ,
69862	 => std_logic_vector(to_unsigned(39,8) ,
69863	 => std_logic_vector(to_unsigned(21,8) ,
69864	 => std_logic_vector(to_unsigned(14,8) ,
69865	 => std_logic_vector(to_unsigned(24,8) ,
69866	 => std_logic_vector(to_unsigned(35,8) ,
69867	 => std_logic_vector(to_unsigned(26,8) ,
69868	 => std_logic_vector(to_unsigned(22,8) ,
69869	 => std_logic_vector(to_unsigned(32,8) ,
69870	 => std_logic_vector(to_unsigned(36,8) ,
69871	 => std_logic_vector(to_unsigned(41,8) ,
69872	 => std_logic_vector(to_unsigned(37,8) ,
69873	 => std_logic_vector(to_unsigned(32,8) ,
69874	 => std_logic_vector(to_unsigned(42,8) ,
69875	 => std_logic_vector(to_unsigned(68,8) ,
69876	 => std_logic_vector(to_unsigned(101,8) ,
69877	 => std_logic_vector(to_unsigned(114,8) ,
69878	 => std_logic_vector(to_unsigned(112,8) ,
69879	 => std_logic_vector(to_unsigned(118,8) ,
69880	 => std_logic_vector(to_unsigned(118,8) ,
69881	 => std_logic_vector(to_unsigned(125,8) ,
69882	 => std_logic_vector(to_unsigned(122,8) ,
69883	 => std_logic_vector(to_unsigned(115,8) ,
69884	 => std_logic_vector(to_unsigned(115,8) ,
69885	 => std_logic_vector(to_unsigned(118,8) ,
69886	 => std_logic_vector(to_unsigned(114,8) ,
69887	 => std_logic_vector(to_unsigned(101,8) ,
69888	 => std_logic_vector(to_unsigned(107,8) ,
69889	 => std_logic_vector(to_unsigned(104,8) ,
69890	 => std_logic_vector(to_unsigned(99,8) ,
69891	 => std_logic_vector(to_unsigned(103,8) ,
69892	 => std_logic_vector(to_unsigned(69,8) ,
69893	 => std_logic_vector(to_unsigned(27,8) ,
69894	 => std_logic_vector(to_unsigned(25,8) ,
69895	 => std_logic_vector(to_unsigned(27,8) ,
69896	 => std_logic_vector(to_unsigned(23,8) ,
69897	 => std_logic_vector(to_unsigned(41,8) ,
69898	 => std_logic_vector(to_unsigned(101,8) ,
69899	 => std_logic_vector(to_unsigned(84,8) ,
69900	 => std_logic_vector(to_unsigned(72,8) ,
69901	 => std_logic_vector(to_unsigned(92,8) ,
69902	 => std_logic_vector(to_unsigned(93,8) ,
69903	 => std_logic_vector(to_unsigned(81,8) ,
69904	 => std_logic_vector(to_unsigned(49,8) ,
69905	 => std_logic_vector(to_unsigned(42,8) ,
69906	 => std_logic_vector(to_unsigned(39,8) ,
69907	 => std_logic_vector(to_unsigned(24,8) ,
69908	 => std_logic_vector(to_unsigned(15,8) ,
69909	 => std_logic_vector(to_unsigned(7,8) ,
69910	 => std_logic_vector(to_unsigned(7,8) ,
69911	 => std_logic_vector(to_unsigned(8,8) ,
69912	 => std_logic_vector(to_unsigned(10,8) ,
69913	 => std_logic_vector(to_unsigned(17,8) ,
69914	 => std_logic_vector(to_unsigned(13,8) ,
69915	 => std_logic_vector(to_unsigned(10,8) ,
69916	 => std_logic_vector(to_unsigned(10,8) ,
69917	 => std_logic_vector(to_unsigned(6,8) ,
69918	 => std_logic_vector(to_unsigned(6,8) ,
69919	 => std_logic_vector(to_unsigned(4,8) ,
69920	 => std_logic_vector(to_unsigned(6,8) ,
69921	 => std_logic_vector(to_unsigned(16,8) ,
69922	 => std_logic_vector(to_unsigned(37,8) ,
69923	 => std_logic_vector(to_unsigned(53,8) ,
69924	 => std_logic_vector(to_unsigned(64,8) ,
69925	 => std_logic_vector(to_unsigned(71,8) ,
69926	 => std_logic_vector(to_unsigned(36,8) ,
69927	 => std_logic_vector(to_unsigned(8,8) ,
69928	 => std_logic_vector(to_unsigned(9,8) ,
69929	 => std_logic_vector(to_unsigned(20,8) ,
69930	 => std_logic_vector(to_unsigned(25,8) ,
69931	 => std_logic_vector(to_unsigned(37,8) ,
69932	 => std_logic_vector(to_unsigned(27,8) ,
69933	 => std_logic_vector(to_unsigned(17,8) ,
69934	 => std_logic_vector(to_unsigned(24,8) ,
69935	 => std_logic_vector(to_unsigned(21,8) ,
69936	 => std_logic_vector(to_unsigned(27,8) ,
69937	 => std_logic_vector(to_unsigned(20,8) ,
69938	 => std_logic_vector(to_unsigned(23,8) ,
69939	 => std_logic_vector(to_unsigned(50,8) ,
69940	 => std_logic_vector(to_unsigned(29,8) ,
69941	 => std_logic_vector(to_unsigned(11,8) ,
69942	 => std_logic_vector(to_unsigned(13,8) ,
69943	 => std_logic_vector(to_unsigned(17,8) ,
69944	 => std_logic_vector(to_unsigned(10,8) ,
69945	 => std_logic_vector(to_unsigned(10,8) ,
69946	 => std_logic_vector(to_unsigned(25,8) ,
69947	 => std_logic_vector(to_unsigned(30,8) ,
69948	 => std_logic_vector(to_unsigned(27,8) ,
69949	 => std_logic_vector(to_unsigned(35,8) ,
69950	 => std_logic_vector(to_unsigned(31,8) ,
69951	 => std_logic_vector(to_unsigned(32,8) ,
69952	 => std_logic_vector(to_unsigned(37,8) ,
69953	 => std_logic_vector(to_unsigned(51,8) ,
69954	 => std_logic_vector(to_unsigned(48,8) ,
69955	 => std_logic_vector(to_unsigned(32,8) ,
69956	 => std_logic_vector(to_unsigned(29,8) ,
69957	 => std_logic_vector(to_unsigned(41,8) ,
69958	 => std_logic_vector(to_unsigned(65,8) ,
69959	 => std_logic_vector(to_unsigned(45,8) ,
69960	 => std_logic_vector(to_unsigned(31,8) ,
69961	 => std_logic_vector(to_unsigned(25,8) ,
69962	 => std_logic_vector(to_unsigned(15,8) ,
69963	 => std_logic_vector(to_unsigned(8,8) ,
69964	 => std_logic_vector(to_unsigned(12,8) ,
69965	 => std_logic_vector(to_unsigned(15,8) ,
69966	 => std_logic_vector(to_unsigned(9,8) ,
69967	 => std_logic_vector(to_unsigned(10,8) ,
69968	 => std_logic_vector(to_unsigned(23,8) ,
69969	 => std_logic_vector(to_unsigned(51,8) ,
69970	 => std_logic_vector(to_unsigned(85,8) ,
69971	 => std_logic_vector(to_unsigned(58,8) ,
69972	 => std_logic_vector(to_unsigned(27,8) ,
69973	 => std_logic_vector(to_unsigned(29,8) ,
69974	 => std_logic_vector(to_unsigned(20,8) ,
69975	 => std_logic_vector(to_unsigned(12,8) ,
69976	 => std_logic_vector(to_unsigned(16,8) ,
69977	 => std_logic_vector(to_unsigned(19,8) ,
69978	 => std_logic_vector(to_unsigned(24,8) ,
69979	 => std_logic_vector(to_unsigned(20,8) ,
69980	 => std_logic_vector(to_unsigned(19,8) ,
69981	 => std_logic_vector(to_unsigned(28,8) ,
69982	 => std_logic_vector(to_unsigned(22,8) ,
69983	 => std_logic_vector(to_unsigned(27,8) ,
69984	 => std_logic_vector(to_unsigned(32,8) ,
69985	 => std_logic_vector(to_unsigned(30,8) ,
69986	 => std_logic_vector(to_unsigned(38,8) ,
69987	 => std_logic_vector(to_unsigned(32,8) ,
69988	 => std_logic_vector(to_unsigned(18,8) ,
69989	 => std_logic_vector(to_unsigned(3,8) ,
69990	 => std_logic_vector(to_unsigned(14,8) ,
69991	 => std_logic_vector(to_unsigned(46,8) ,
69992	 => std_logic_vector(to_unsigned(37,8) ,
69993	 => std_logic_vector(to_unsigned(30,8) ,
69994	 => std_logic_vector(to_unsigned(36,8) ,
69995	 => std_logic_vector(to_unsigned(52,8) ,
69996	 => std_logic_vector(to_unsigned(37,8) ,
69997	 => std_logic_vector(to_unsigned(41,8) ,
69998	 => std_logic_vector(to_unsigned(63,8) ,
69999	 => std_logic_vector(to_unsigned(65,8) ,
70000	 => std_logic_vector(to_unsigned(43,8) ,
70001	 => std_logic_vector(to_unsigned(39,8) ,
70002	 => std_logic_vector(to_unsigned(43,8) ,
70003	 => std_logic_vector(to_unsigned(78,8) ,
70004	 => std_logic_vector(to_unsigned(105,8) ,
70005	 => std_logic_vector(to_unsigned(100,8) ,
70006	 => std_logic_vector(to_unsigned(49,8) ,
70007	 => std_logic_vector(to_unsigned(73,8) ,
70008	 => std_logic_vector(to_unsigned(128,8) ,
70009	 => std_logic_vector(to_unsigned(119,8) ,
70010	 => std_logic_vector(to_unsigned(33,8) ,
70011	 => std_logic_vector(to_unsigned(11,8) ,
70012	 => std_logic_vector(to_unsigned(22,8) ,
70013	 => std_logic_vector(to_unsigned(30,8) ,
70014	 => std_logic_vector(to_unsigned(20,8) ,
70015	 => std_logic_vector(to_unsigned(23,8) ,
70016	 => std_logic_vector(to_unsigned(38,8) ,
70017	 => std_logic_vector(to_unsigned(41,8) ,
70018	 => std_logic_vector(to_unsigned(39,8) ,
70019	 => std_logic_vector(to_unsigned(37,8) ,
70020	 => std_logic_vector(to_unsigned(28,8) ,
70021	 => std_logic_vector(to_unsigned(36,8) ,
70022	 => std_logic_vector(to_unsigned(36,8) ,
70023	 => std_logic_vector(to_unsigned(42,8) ,
70024	 => std_logic_vector(to_unsigned(42,8) ,
70025	 => std_logic_vector(to_unsigned(32,8) ,
70026	 => std_logic_vector(to_unsigned(10,8) ,
70027	 => std_logic_vector(to_unsigned(9,8) ,
70028	 => std_logic_vector(to_unsigned(25,8) ,
70029	 => std_logic_vector(to_unsigned(13,8) ,
70030	 => std_logic_vector(to_unsigned(10,8) ,
70031	 => std_logic_vector(to_unsigned(16,8) ,
70032	 => std_logic_vector(to_unsigned(23,8) ,
70033	 => std_logic_vector(to_unsigned(29,8) ,
70034	 => std_logic_vector(to_unsigned(23,8) ,
70035	 => std_logic_vector(to_unsigned(2,8) ,
70036	 => std_logic_vector(to_unsigned(0,8) ,
70037	 => std_logic_vector(to_unsigned(5,8) ,
70038	 => std_logic_vector(to_unsigned(29,8) ,
70039	 => std_logic_vector(to_unsigned(47,8) ,
70040	 => std_logic_vector(to_unsigned(41,8) ,
70041	 => std_logic_vector(to_unsigned(20,8) ,
70042	 => std_logic_vector(to_unsigned(8,8) ,
70043	 => std_logic_vector(to_unsigned(5,8) ,
70044	 => std_logic_vector(to_unsigned(4,8) ,
70045	 => std_logic_vector(to_unsigned(12,8) ,
70046	 => std_logic_vector(to_unsigned(3,8) ,
70047	 => std_logic_vector(to_unsigned(0,8) ,
70048	 => std_logic_vector(to_unsigned(2,8) ,
70049	 => std_logic_vector(to_unsigned(24,8) ,
70050	 => std_logic_vector(to_unsigned(15,8) ,
70051	 => std_logic_vector(to_unsigned(0,8) ,
70052	 => std_logic_vector(to_unsigned(0,8) ,
70053	 => std_logic_vector(to_unsigned(0,8) ,
70054	 => std_logic_vector(to_unsigned(1,8) ,
70055	 => std_logic_vector(to_unsigned(0,8) ,
70056	 => std_logic_vector(to_unsigned(0,8) ,
70057	 => std_logic_vector(to_unsigned(1,8) ,
70058	 => std_logic_vector(to_unsigned(0,8) ,
70059	 => std_logic_vector(to_unsigned(0,8) ,
70060	 => std_logic_vector(to_unsigned(3,8) ,
70061	 => std_logic_vector(to_unsigned(11,8) ,
70062	 => std_logic_vector(to_unsigned(2,8) ,
70063	 => std_logic_vector(to_unsigned(0,8) ,
70064	 => std_logic_vector(to_unsigned(23,8) ,
70065	 => std_logic_vector(to_unsigned(104,8) ,
70066	 => std_logic_vector(to_unsigned(47,8) ,
70067	 => std_logic_vector(to_unsigned(33,8) ,
70068	 => std_logic_vector(to_unsigned(27,8) ,
70069	 => std_logic_vector(to_unsigned(13,8) ,
70070	 => std_logic_vector(to_unsigned(11,8) ,
70071	 => std_logic_vector(to_unsigned(12,8) ,
70072	 => std_logic_vector(to_unsigned(15,8) ,
70073	 => std_logic_vector(to_unsigned(15,8) ,
70074	 => std_logic_vector(to_unsigned(12,8) ,
70075	 => std_logic_vector(to_unsigned(12,8) ,
70076	 => std_logic_vector(to_unsigned(10,8) ,
70077	 => std_logic_vector(to_unsigned(8,8) ,
70078	 => std_logic_vector(to_unsigned(24,8) ,
70079	 => std_logic_vector(to_unsigned(18,8) ,
70080	 => std_logic_vector(to_unsigned(7,8) ,
70081	 => std_logic_vector(to_unsigned(87,8) ,
70082	 => std_logic_vector(to_unsigned(103,8) ,
70083	 => std_logic_vector(to_unsigned(112,8) ,
70084	 => std_logic_vector(to_unsigned(81,8) ,
70085	 => std_logic_vector(to_unsigned(85,8) ,
70086	 => std_logic_vector(to_unsigned(78,8) ,
70087	 => std_logic_vector(to_unsigned(69,8) ,
70088	 => std_logic_vector(to_unsigned(58,8) ,
70089	 => std_logic_vector(to_unsigned(62,8) ,
70090	 => std_logic_vector(to_unsigned(73,8) ,
70091	 => std_logic_vector(to_unsigned(77,8) ,
70092	 => std_logic_vector(to_unsigned(53,8) ,
70093	 => std_logic_vector(to_unsigned(44,8) ,
70094	 => std_logic_vector(to_unsigned(54,8) ,
70095	 => std_logic_vector(to_unsigned(50,8) ,
70096	 => std_logic_vector(to_unsigned(54,8) ,
70097	 => std_logic_vector(to_unsigned(59,8) ,
70098	 => std_logic_vector(to_unsigned(56,8) ,
70099	 => std_logic_vector(to_unsigned(37,8) ,
70100	 => std_logic_vector(to_unsigned(37,8) ,
70101	 => std_logic_vector(to_unsigned(41,8) ,
70102	 => std_logic_vector(to_unsigned(38,8) ,
70103	 => std_logic_vector(to_unsigned(56,8) ,
70104	 => std_logic_vector(to_unsigned(100,8) ,
70105	 => std_logic_vector(to_unsigned(96,8) ,
70106	 => std_logic_vector(to_unsigned(45,8) ,
70107	 => std_logic_vector(to_unsigned(35,8) ,
70108	 => std_logic_vector(to_unsigned(27,8) ,
70109	 => std_logic_vector(to_unsigned(37,8) ,
70110	 => std_logic_vector(to_unsigned(46,8) ,
70111	 => std_logic_vector(to_unsigned(45,8) ,
70112	 => std_logic_vector(to_unsigned(47,8) ,
70113	 => std_logic_vector(to_unsigned(32,8) ,
70114	 => std_logic_vector(to_unsigned(13,8) ,
70115	 => std_logic_vector(to_unsigned(15,8) ,
70116	 => std_logic_vector(to_unsigned(16,8) ,
70117	 => std_logic_vector(to_unsigned(23,8) ,
70118	 => std_logic_vector(to_unsigned(30,8) ,
70119	 => std_logic_vector(to_unsigned(20,8) ,
70120	 => std_logic_vector(to_unsigned(29,8) ,
70121	 => std_logic_vector(to_unsigned(32,8) ,
70122	 => std_logic_vector(to_unsigned(33,8) ,
70123	 => std_logic_vector(to_unsigned(38,8) ,
70124	 => std_logic_vector(to_unsigned(28,8) ,
70125	 => std_logic_vector(to_unsigned(19,8) ,
70126	 => std_logic_vector(to_unsigned(19,8) ,
70127	 => std_logic_vector(to_unsigned(19,8) ,
70128	 => std_logic_vector(to_unsigned(21,8) ,
70129	 => std_logic_vector(to_unsigned(27,8) ,
70130	 => std_logic_vector(to_unsigned(33,8) ,
70131	 => std_logic_vector(to_unsigned(30,8) ,
70132	 => std_logic_vector(to_unsigned(34,8) ,
70133	 => std_logic_vector(to_unsigned(43,8) ,
70134	 => std_logic_vector(to_unsigned(39,8) ,
70135	 => std_logic_vector(to_unsigned(34,8) ,
70136	 => std_logic_vector(to_unsigned(37,8) ,
70137	 => std_logic_vector(to_unsigned(46,8) ,
70138	 => std_logic_vector(to_unsigned(37,8) ,
70139	 => std_logic_vector(to_unsigned(40,8) ,
70140	 => std_logic_vector(to_unsigned(51,8) ,
70141	 => std_logic_vector(to_unsigned(60,8) ,
70142	 => std_logic_vector(to_unsigned(45,8) ,
70143	 => std_logic_vector(to_unsigned(46,8) ,
70144	 => std_logic_vector(to_unsigned(47,8) ,
70145	 => std_logic_vector(to_unsigned(51,8) ,
70146	 => std_logic_vector(to_unsigned(48,8) ,
70147	 => std_logic_vector(to_unsigned(45,8) ,
70148	 => std_logic_vector(to_unsigned(43,8) ,
70149	 => std_logic_vector(to_unsigned(44,8) ,
70150	 => std_logic_vector(to_unsigned(45,8) ,
70151	 => std_logic_vector(to_unsigned(54,8) ,
70152	 => std_logic_vector(to_unsigned(40,8) ,
70153	 => std_logic_vector(to_unsigned(48,8) ,
70154	 => std_logic_vector(to_unsigned(52,8) ,
70155	 => std_logic_vector(to_unsigned(45,8) ,
70156	 => std_logic_vector(to_unsigned(47,8) ,
70157	 => std_logic_vector(to_unsigned(59,8) ,
70158	 => std_logic_vector(to_unsigned(59,8) ,
70159	 => std_logic_vector(to_unsigned(55,8) ,
70160	 => std_logic_vector(to_unsigned(52,8) ,
70161	 => std_logic_vector(to_unsigned(63,8) ,
70162	 => std_logic_vector(to_unsigned(41,8) ,
70163	 => std_logic_vector(to_unsigned(88,8) ,
70164	 => std_logic_vector(to_unsigned(88,8) ,
70165	 => std_logic_vector(to_unsigned(79,8) ,
70166	 => std_logic_vector(to_unsigned(76,8) ,
70167	 => std_logic_vector(to_unsigned(66,8) ,
70168	 => std_logic_vector(to_unsigned(51,8) ,
70169	 => std_logic_vector(to_unsigned(37,8) ,
70170	 => std_logic_vector(to_unsigned(20,8) ,
70171	 => std_logic_vector(to_unsigned(23,8) ,
70172	 => std_logic_vector(to_unsigned(40,8) ,
70173	 => std_logic_vector(to_unsigned(29,8) ,
70174	 => std_logic_vector(to_unsigned(24,8) ,
70175	 => std_logic_vector(to_unsigned(30,8) ,
70176	 => std_logic_vector(to_unsigned(38,8) ,
70177	 => std_logic_vector(to_unsigned(35,8) ,
70178	 => std_logic_vector(to_unsigned(38,8) ,
70179	 => std_logic_vector(to_unsigned(43,8) ,
70180	 => std_logic_vector(to_unsigned(40,8) ,
70181	 => std_logic_vector(to_unsigned(45,8) ,
70182	 => std_logic_vector(to_unsigned(37,8) ,
70183	 => std_logic_vector(to_unsigned(24,8) ,
70184	 => std_logic_vector(to_unsigned(25,8) ,
70185	 => std_logic_vector(to_unsigned(39,8) ,
70186	 => std_logic_vector(to_unsigned(35,8) ,
70187	 => std_logic_vector(to_unsigned(34,8) ,
70188	 => std_logic_vector(to_unsigned(37,8) ,
70189	 => std_logic_vector(to_unsigned(66,8) ,
70190	 => std_logic_vector(to_unsigned(51,8) ,
70191	 => std_logic_vector(to_unsigned(51,8) ,
70192	 => std_logic_vector(to_unsigned(114,8) ,
70193	 => std_logic_vector(to_unsigned(115,8) ,
70194	 => std_logic_vector(to_unsigned(104,8) ,
70195	 => std_logic_vector(to_unsigned(74,8) ,
70196	 => std_logic_vector(to_unsigned(86,8) ,
70197	 => std_logic_vector(to_unsigned(116,8) ,
70198	 => std_logic_vector(to_unsigned(111,8) ,
70199	 => std_logic_vector(to_unsigned(114,8) ,
70200	 => std_logic_vector(to_unsigned(116,8) ,
70201	 => std_logic_vector(to_unsigned(116,8) ,
70202	 => std_logic_vector(to_unsigned(118,8) ,
70203	 => std_logic_vector(to_unsigned(114,8) ,
70204	 => std_logic_vector(to_unsigned(107,8) ,
70205	 => std_logic_vector(to_unsigned(105,8) ,
70206	 => std_logic_vector(to_unsigned(101,8) ,
70207	 => std_logic_vector(to_unsigned(93,8) ,
70208	 => std_logic_vector(to_unsigned(101,8) ,
70209	 => std_logic_vector(to_unsigned(104,8) ,
70210	 => std_logic_vector(to_unsigned(101,8) ,
70211	 => std_logic_vector(to_unsigned(104,8) ,
70212	 => std_logic_vector(to_unsigned(46,8) ,
70213	 => std_logic_vector(to_unsigned(19,8) ,
70214	 => std_logic_vector(to_unsigned(35,8) ,
70215	 => std_logic_vector(to_unsigned(17,8) ,
70216	 => std_logic_vector(to_unsigned(39,8) ,
70217	 => std_logic_vector(to_unsigned(101,8) ,
70218	 => std_logic_vector(to_unsigned(100,8) ,
70219	 => std_logic_vector(to_unsigned(95,8) ,
70220	 => std_logic_vector(to_unsigned(99,8) ,
70221	 => std_logic_vector(to_unsigned(96,8) ,
70222	 => std_logic_vector(to_unsigned(95,8) ,
70223	 => std_logic_vector(to_unsigned(96,8) ,
70224	 => std_logic_vector(to_unsigned(91,8) ,
70225	 => std_logic_vector(to_unsigned(82,8) ,
70226	 => std_logic_vector(to_unsigned(67,8) ,
70227	 => std_logic_vector(to_unsigned(47,8) ,
70228	 => std_logic_vector(to_unsigned(36,8) ,
70229	 => std_logic_vector(to_unsigned(30,8) ,
70230	 => std_logic_vector(to_unsigned(21,8) ,
70231	 => std_logic_vector(to_unsigned(14,8) ,
70232	 => std_logic_vector(to_unsigned(10,8) ,
70233	 => std_logic_vector(to_unsigned(10,8) ,
70234	 => std_logic_vector(to_unsigned(9,8) ,
70235	 => std_logic_vector(to_unsigned(10,8) ,
70236	 => std_logic_vector(to_unsigned(9,8) ,
70237	 => std_logic_vector(to_unsigned(5,8) ,
70238	 => std_logic_vector(to_unsigned(5,8) ,
70239	 => std_logic_vector(to_unsigned(3,8) ,
70240	 => std_logic_vector(to_unsigned(7,8) ,
70241	 => std_logic_vector(to_unsigned(25,8) ,
70242	 => std_logic_vector(to_unsigned(49,8) ,
70243	 => std_logic_vector(to_unsigned(65,8) ,
70244	 => std_logic_vector(to_unsigned(65,8) ,
70245	 => std_logic_vector(to_unsigned(68,8) ,
70246	 => std_logic_vector(to_unsigned(37,8) ,
70247	 => std_logic_vector(to_unsigned(5,8) ,
70248	 => std_logic_vector(to_unsigned(7,8) ,
70249	 => std_logic_vector(to_unsigned(14,8) ,
70250	 => std_logic_vector(to_unsigned(23,8) ,
70251	 => std_logic_vector(to_unsigned(22,8) ,
70252	 => std_logic_vector(to_unsigned(19,8) ,
70253	 => std_logic_vector(to_unsigned(29,8) ,
70254	 => std_logic_vector(to_unsigned(15,8) ,
70255	 => std_logic_vector(to_unsigned(23,8) ,
70256	 => std_logic_vector(to_unsigned(19,8) ,
70257	 => std_logic_vector(to_unsigned(20,8) ,
70258	 => std_logic_vector(to_unsigned(42,8) ,
70259	 => std_logic_vector(to_unsigned(23,8) ,
70260	 => std_logic_vector(to_unsigned(23,8) ,
70261	 => std_logic_vector(to_unsigned(18,8) ,
70262	 => std_logic_vector(to_unsigned(17,8) ,
70263	 => std_logic_vector(to_unsigned(18,8) ,
70264	 => std_logic_vector(to_unsigned(13,8) ,
70265	 => std_logic_vector(to_unsigned(14,8) ,
70266	 => std_logic_vector(to_unsigned(30,8) ,
70267	 => std_logic_vector(to_unsigned(22,8) ,
70268	 => std_logic_vector(to_unsigned(13,8) ,
70269	 => std_logic_vector(to_unsigned(19,8) ,
70270	 => std_logic_vector(to_unsigned(30,8) ,
70271	 => std_logic_vector(to_unsigned(32,8) ,
70272	 => std_logic_vector(to_unsigned(27,8) ,
70273	 => std_logic_vector(to_unsigned(34,8) ,
70274	 => std_logic_vector(to_unsigned(40,8) ,
70275	 => std_logic_vector(to_unsigned(30,8) ,
70276	 => std_logic_vector(to_unsigned(32,8) ,
70277	 => std_logic_vector(to_unsigned(42,8) ,
70278	 => std_logic_vector(to_unsigned(67,8) ,
70279	 => std_logic_vector(to_unsigned(61,8) ,
70280	 => std_logic_vector(to_unsigned(32,8) ,
70281	 => std_logic_vector(to_unsigned(28,8) ,
70282	 => std_logic_vector(to_unsigned(15,8) ,
70283	 => std_logic_vector(to_unsigned(9,8) ,
70284	 => std_logic_vector(to_unsigned(13,8) ,
70285	 => std_logic_vector(to_unsigned(16,8) ,
70286	 => std_logic_vector(to_unsigned(11,8) ,
70287	 => std_logic_vector(to_unsigned(9,8) ,
70288	 => std_logic_vector(to_unsigned(24,8) ,
70289	 => std_logic_vector(to_unsigned(33,8) ,
70290	 => std_logic_vector(to_unsigned(43,8) ,
70291	 => std_logic_vector(to_unsigned(38,8) ,
70292	 => std_logic_vector(to_unsigned(24,8) ,
70293	 => std_logic_vector(to_unsigned(28,8) ,
70294	 => std_logic_vector(to_unsigned(33,8) ,
70295	 => std_logic_vector(to_unsigned(25,8) ,
70296	 => std_logic_vector(to_unsigned(17,8) ,
70297	 => std_logic_vector(to_unsigned(17,8) ,
70298	 => std_logic_vector(to_unsigned(25,8) ,
70299	 => std_logic_vector(to_unsigned(22,8) ,
70300	 => std_logic_vector(to_unsigned(8,8) ,
70301	 => std_logic_vector(to_unsigned(6,8) ,
70302	 => std_logic_vector(to_unsigned(12,8) ,
70303	 => std_logic_vector(to_unsigned(34,8) ,
70304	 => std_logic_vector(to_unsigned(41,8) ,
70305	 => std_logic_vector(to_unsigned(33,8) ,
70306	 => std_logic_vector(to_unsigned(31,8) ,
70307	 => std_logic_vector(to_unsigned(35,8) ,
70308	 => std_logic_vector(to_unsigned(17,8) ,
70309	 => std_logic_vector(to_unsigned(3,8) ,
70310	 => std_logic_vector(to_unsigned(15,8) ,
70311	 => std_logic_vector(to_unsigned(35,8) ,
70312	 => std_logic_vector(to_unsigned(16,8) ,
70313	 => std_logic_vector(to_unsigned(25,8) ,
70314	 => std_logic_vector(to_unsigned(33,8) ,
70315	 => std_logic_vector(to_unsigned(49,8) ,
70316	 => std_logic_vector(to_unsigned(51,8) ,
70317	 => std_logic_vector(to_unsigned(48,8) ,
70318	 => std_logic_vector(to_unsigned(56,8) ,
70319	 => std_logic_vector(to_unsigned(58,8) ,
70320	 => std_logic_vector(to_unsigned(37,8) ,
70321	 => std_logic_vector(to_unsigned(36,8) ,
70322	 => std_logic_vector(to_unsigned(45,8) ,
70323	 => std_logic_vector(to_unsigned(74,8) ,
70324	 => std_logic_vector(to_unsigned(100,8) ,
70325	 => std_logic_vector(to_unsigned(101,8) ,
70326	 => std_logic_vector(to_unsigned(42,8) ,
70327	 => std_logic_vector(to_unsigned(70,8) ,
70328	 => std_logic_vector(to_unsigned(130,8) ,
70329	 => std_logic_vector(to_unsigned(121,8) ,
70330	 => std_logic_vector(to_unsigned(29,8) ,
70331	 => std_logic_vector(to_unsigned(5,8) ,
70332	 => std_logic_vector(to_unsigned(9,8) ,
70333	 => std_logic_vector(to_unsigned(8,8) ,
70334	 => std_logic_vector(to_unsigned(7,8) ,
70335	 => std_logic_vector(to_unsigned(10,8) ,
70336	 => std_logic_vector(to_unsigned(14,8) ,
70337	 => std_logic_vector(to_unsigned(20,8) ,
70338	 => std_logic_vector(to_unsigned(20,8) ,
70339	 => std_logic_vector(to_unsigned(27,8) ,
70340	 => std_logic_vector(to_unsigned(39,8) ,
70341	 => std_logic_vector(to_unsigned(52,8) ,
70342	 => std_logic_vector(to_unsigned(51,8) ,
70343	 => std_logic_vector(to_unsigned(40,8) ,
70344	 => std_logic_vector(to_unsigned(37,8) ,
70345	 => std_logic_vector(to_unsigned(51,8) ,
70346	 => std_logic_vector(to_unsigned(45,8) ,
70347	 => std_logic_vector(to_unsigned(37,8) ,
70348	 => std_logic_vector(to_unsigned(32,8) ,
70349	 => std_logic_vector(to_unsigned(17,8) ,
70350	 => std_logic_vector(to_unsigned(22,8) ,
70351	 => std_logic_vector(to_unsigned(13,8) ,
70352	 => std_logic_vector(to_unsigned(10,8) ,
70353	 => std_logic_vector(to_unsigned(20,8) ,
70354	 => std_logic_vector(to_unsigned(23,8) ,
70355	 => std_logic_vector(to_unsigned(3,8) ,
70356	 => std_logic_vector(to_unsigned(0,8) ,
70357	 => std_logic_vector(to_unsigned(2,8) ,
70358	 => std_logic_vector(to_unsigned(19,8) ,
70359	 => std_logic_vector(to_unsigned(13,8) ,
70360	 => std_logic_vector(to_unsigned(8,8) ,
70361	 => std_logic_vector(to_unsigned(7,8) ,
70362	 => std_logic_vector(to_unsigned(6,8) ,
70363	 => std_logic_vector(to_unsigned(4,8) ,
70364	 => std_logic_vector(to_unsigned(4,8) ,
70365	 => std_logic_vector(to_unsigned(12,8) ,
70366	 => std_logic_vector(to_unsigned(5,8) ,
70367	 => std_logic_vector(to_unsigned(0,8) ,
70368	 => std_logic_vector(to_unsigned(1,8) ,
70369	 => std_logic_vector(to_unsigned(3,8) ,
70370	 => std_logic_vector(to_unsigned(0,8) ,
70371	 => std_logic_vector(to_unsigned(0,8) ,
70372	 => std_logic_vector(to_unsigned(1,8) ,
70373	 => std_logic_vector(to_unsigned(1,8) ,
70374	 => std_logic_vector(to_unsigned(2,8) ,
70375	 => std_logic_vector(to_unsigned(3,8) ,
70376	 => std_logic_vector(to_unsigned(3,8) ,
70377	 => std_logic_vector(to_unsigned(3,8) ,
70378	 => std_logic_vector(to_unsigned(2,8) ,
70379	 => std_logic_vector(to_unsigned(0,8) ,
70380	 => std_logic_vector(to_unsigned(0,8) ,
70381	 => std_logic_vector(to_unsigned(1,8) ,
70382	 => std_logic_vector(to_unsigned(1,8) ,
70383	 => std_logic_vector(to_unsigned(0,8) ,
70384	 => std_logic_vector(to_unsigned(7,8) ,
70385	 => std_logic_vector(to_unsigned(86,8) ,
70386	 => std_logic_vector(to_unsigned(56,8) ,
70387	 => std_logic_vector(to_unsigned(64,8) ,
70388	 => std_logic_vector(to_unsigned(62,8) ,
70389	 => std_logic_vector(to_unsigned(23,8) ,
70390	 => std_logic_vector(to_unsigned(13,8) ,
70391	 => std_logic_vector(to_unsigned(23,8) ,
70392	 => std_logic_vector(to_unsigned(12,8) ,
70393	 => std_logic_vector(to_unsigned(16,8) ,
70394	 => std_logic_vector(to_unsigned(12,8) ,
70395	 => std_logic_vector(to_unsigned(6,8) ,
70396	 => std_logic_vector(to_unsigned(6,8) ,
70397	 => std_logic_vector(to_unsigned(6,8) ,
70398	 => std_logic_vector(to_unsigned(10,8) ,
70399	 => std_logic_vector(to_unsigned(12,8) ,
70400	 => std_logic_vector(to_unsigned(11,8) ,
70401	 => std_logic_vector(to_unsigned(115,8) ,
70402	 => std_logic_vector(to_unsigned(104,8) ,
70403	 => std_logic_vector(to_unsigned(100,8) ,
70404	 => std_logic_vector(to_unsigned(103,8) ,
70405	 => std_logic_vector(to_unsigned(96,8) ,
70406	 => std_logic_vector(to_unsigned(91,8) ,
70407	 => std_logic_vector(to_unsigned(81,8) ,
70408	 => std_logic_vector(to_unsigned(86,8) ,
70409	 => std_logic_vector(to_unsigned(79,8) ,
70410	 => std_logic_vector(to_unsigned(70,8) ,
70411	 => std_logic_vector(to_unsigned(63,8) ,
70412	 => std_logic_vector(to_unsigned(46,8) ,
70413	 => std_logic_vector(to_unsigned(34,8) ,
70414	 => std_logic_vector(to_unsigned(32,8) ,
70415	 => std_logic_vector(to_unsigned(39,8) ,
70416	 => std_logic_vector(to_unsigned(41,8) ,
70417	 => std_logic_vector(to_unsigned(66,8) ,
70418	 => std_logic_vector(to_unsigned(74,8) ,
70419	 => std_logic_vector(to_unsigned(66,8) ,
70420	 => std_logic_vector(to_unsigned(77,8) ,
70421	 => std_logic_vector(to_unsigned(58,8) ,
70422	 => std_logic_vector(to_unsigned(24,8) ,
70423	 => std_logic_vector(to_unsigned(27,8) ,
70424	 => std_logic_vector(to_unsigned(32,8) ,
70425	 => std_logic_vector(to_unsigned(42,8) ,
70426	 => std_logic_vector(to_unsigned(39,8) ,
70427	 => std_logic_vector(to_unsigned(38,8) ,
70428	 => std_logic_vector(to_unsigned(33,8) ,
70429	 => std_logic_vector(to_unsigned(35,8) ,
70430	 => std_logic_vector(to_unsigned(37,8) ,
70431	 => std_logic_vector(to_unsigned(33,8) ,
70432	 => std_logic_vector(to_unsigned(35,8) ,
70433	 => std_logic_vector(to_unsigned(49,8) ,
70434	 => std_logic_vector(to_unsigned(40,8) ,
70435	 => std_logic_vector(to_unsigned(24,8) ,
70436	 => std_logic_vector(to_unsigned(12,8) ,
70437	 => std_logic_vector(to_unsigned(13,8) ,
70438	 => std_logic_vector(to_unsigned(37,8) ,
70439	 => std_logic_vector(to_unsigned(17,8) ,
70440	 => std_logic_vector(to_unsigned(19,8) ,
70441	 => std_logic_vector(to_unsigned(20,8) ,
70442	 => std_logic_vector(to_unsigned(18,8) ,
70443	 => std_logic_vector(to_unsigned(21,8) ,
70444	 => std_logic_vector(to_unsigned(21,8) ,
70445	 => std_logic_vector(to_unsigned(24,8) ,
70446	 => std_logic_vector(to_unsigned(23,8) ,
70447	 => std_logic_vector(to_unsigned(22,8) ,
70448	 => std_logic_vector(to_unsigned(22,8) ,
70449	 => std_logic_vector(to_unsigned(25,8) ,
70450	 => std_logic_vector(to_unsigned(32,8) ,
70451	 => std_logic_vector(to_unsigned(33,8) ,
70452	 => std_logic_vector(to_unsigned(35,8) ,
70453	 => std_logic_vector(to_unsigned(41,8) ,
70454	 => std_logic_vector(to_unsigned(37,8) ,
70455	 => std_logic_vector(to_unsigned(28,8) ,
70456	 => std_logic_vector(to_unsigned(33,8) ,
70457	 => std_logic_vector(to_unsigned(45,8) ,
70458	 => std_logic_vector(to_unsigned(40,8) ,
70459	 => std_logic_vector(to_unsigned(48,8) ,
70460	 => std_logic_vector(to_unsigned(54,8) ,
70461	 => std_logic_vector(to_unsigned(61,8) ,
70462	 => std_logic_vector(to_unsigned(51,8) ,
70463	 => std_logic_vector(to_unsigned(50,8) ,
70464	 => std_logic_vector(to_unsigned(68,8) ,
70465	 => std_logic_vector(to_unsigned(57,8) ,
70466	 => std_logic_vector(to_unsigned(50,8) ,
70467	 => std_logic_vector(to_unsigned(42,8) ,
70468	 => std_logic_vector(to_unsigned(37,8) ,
70469	 => std_logic_vector(to_unsigned(41,8) ,
70470	 => std_logic_vector(to_unsigned(42,8) ,
70471	 => std_logic_vector(to_unsigned(41,8) ,
70472	 => std_logic_vector(to_unsigned(39,8) ,
70473	 => std_logic_vector(to_unsigned(42,8) ,
70474	 => std_logic_vector(to_unsigned(51,8) ,
70475	 => std_logic_vector(to_unsigned(48,8) ,
70476	 => std_logic_vector(to_unsigned(44,8) ,
70477	 => std_logic_vector(to_unsigned(58,8) ,
70478	 => std_logic_vector(to_unsigned(68,8) ,
70479	 => std_logic_vector(to_unsigned(68,8) ,
70480	 => std_logic_vector(to_unsigned(71,8) ,
70481	 => std_logic_vector(to_unsigned(79,8) ,
70482	 => std_logic_vector(to_unsigned(51,8) ,
70483	 => std_logic_vector(to_unsigned(77,8) ,
70484	 => std_logic_vector(to_unsigned(88,8) ,
70485	 => std_logic_vector(to_unsigned(80,8) ,
70486	 => std_logic_vector(to_unsigned(74,8) ,
70487	 => std_logic_vector(to_unsigned(68,8) ,
70488	 => std_logic_vector(to_unsigned(49,8) ,
70489	 => std_logic_vector(to_unsigned(32,8) ,
70490	 => std_logic_vector(to_unsigned(24,8) ,
70491	 => std_logic_vector(to_unsigned(40,8) ,
70492	 => std_logic_vector(to_unsigned(42,8) ,
70493	 => std_logic_vector(to_unsigned(27,8) ,
70494	 => std_logic_vector(to_unsigned(21,8) ,
70495	 => std_logic_vector(to_unsigned(32,8) ,
70496	 => std_logic_vector(to_unsigned(25,8) ,
70497	 => std_logic_vector(to_unsigned(21,8) ,
70498	 => std_logic_vector(to_unsigned(32,8) ,
70499	 => std_logic_vector(to_unsigned(34,8) ,
70500	 => std_logic_vector(to_unsigned(37,8) ,
70501	 => std_logic_vector(to_unsigned(35,8) ,
70502	 => std_logic_vector(to_unsigned(32,8) ,
70503	 => std_logic_vector(to_unsigned(32,8) ,
70504	 => std_logic_vector(to_unsigned(30,8) ,
70505	 => std_logic_vector(to_unsigned(35,8) ,
70506	 => std_logic_vector(to_unsigned(35,8) ,
70507	 => std_logic_vector(to_unsigned(53,8) ,
70508	 => std_logic_vector(to_unsigned(53,8) ,
70509	 => std_logic_vector(to_unsigned(51,8) ,
70510	 => std_logic_vector(to_unsigned(35,8) ,
70511	 => std_logic_vector(to_unsigned(35,8) ,
70512	 => std_logic_vector(to_unsigned(99,8) ,
70513	 => std_logic_vector(to_unsigned(141,8) ,
70514	 => std_logic_vector(to_unsigned(114,8) ,
70515	 => std_logic_vector(to_unsigned(46,8) ,
70516	 => std_logic_vector(to_unsigned(74,8) ,
70517	 => std_logic_vector(to_unsigned(119,8) ,
70518	 => std_logic_vector(to_unsigned(105,8) ,
70519	 => std_logic_vector(to_unsigned(115,8) ,
70520	 => std_logic_vector(to_unsigned(119,8) ,
70521	 => std_logic_vector(to_unsigned(115,8) ,
70522	 => std_logic_vector(to_unsigned(119,8) ,
70523	 => std_logic_vector(to_unsigned(119,8) ,
70524	 => std_logic_vector(to_unsigned(111,8) ,
70525	 => std_logic_vector(to_unsigned(105,8) ,
70526	 => std_logic_vector(to_unsigned(101,8) ,
70527	 => std_logic_vector(to_unsigned(93,8) ,
70528	 => std_logic_vector(to_unsigned(101,8) ,
70529	 => std_logic_vector(to_unsigned(107,8) ,
70530	 => std_logic_vector(to_unsigned(93,8) ,
70531	 => std_logic_vector(to_unsigned(93,8) ,
70532	 => std_logic_vector(to_unsigned(67,8) ,
70533	 => std_logic_vector(to_unsigned(49,8) ,
70534	 => std_logic_vector(to_unsigned(64,8) ,
70535	 => std_logic_vector(to_unsigned(60,8) ,
70536	 => std_logic_vector(to_unsigned(91,8) ,
70537	 => std_logic_vector(to_unsigned(95,8) ,
70538	 => std_logic_vector(to_unsigned(93,8) ,
70539	 => std_logic_vector(to_unsigned(99,8) ,
70540	 => std_logic_vector(to_unsigned(103,8) ,
70541	 => std_logic_vector(to_unsigned(99,8) ,
70542	 => std_logic_vector(to_unsigned(101,8) ,
70543	 => std_logic_vector(to_unsigned(101,8) ,
70544	 => std_logic_vector(to_unsigned(97,8) ,
70545	 => std_logic_vector(to_unsigned(95,8) ,
70546	 => std_logic_vector(to_unsigned(99,8) ,
70547	 => std_logic_vector(to_unsigned(95,8) ,
70548	 => std_logic_vector(to_unsigned(81,8) ,
70549	 => std_logic_vector(to_unsigned(74,8) ,
70550	 => std_logic_vector(to_unsigned(71,8) ,
70551	 => std_logic_vector(to_unsigned(64,8) ,
70552	 => std_logic_vector(to_unsigned(47,8) ,
70553	 => std_logic_vector(to_unsigned(37,8) ,
70554	 => std_logic_vector(to_unsigned(23,8) ,
70555	 => std_logic_vector(to_unsigned(12,8) ,
70556	 => std_logic_vector(to_unsigned(10,8) ,
70557	 => std_logic_vector(to_unsigned(7,8) ,
70558	 => std_logic_vector(to_unsigned(6,8) ,
70559	 => std_logic_vector(to_unsigned(7,8) ,
70560	 => std_logic_vector(to_unsigned(11,8) ,
70561	 => std_logic_vector(to_unsigned(29,8) ,
70562	 => std_logic_vector(to_unsigned(44,8) ,
70563	 => std_logic_vector(to_unsigned(64,8) ,
70564	 => std_logic_vector(to_unsigned(72,8) ,
70565	 => std_logic_vector(to_unsigned(68,8) ,
70566	 => std_logic_vector(to_unsigned(35,8) ,
70567	 => std_logic_vector(to_unsigned(5,8) ,
70568	 => std_logic_vector(to_unsigned(5,8) ,
70569	 => std_logic_vector(to_unsigned(13,8) ,
70570	 => std_logic_vector(to_unsigned(14,8) ,
70571	 => std_logic_vector(to_unsigned(23,8) ,
70572	 => std_logic_vector(to_unsigned(28,8) ,
70573	 => std_logic_vector(to_unsigned(14,8) ,
70574	 => std_logic_vector(to_unsigned(22,8) ,
70575	 => std_logic_vector(to_unsigned(23,8) ,
70576	 => std_logic_vector(to_unsigned(16,8) ,
70577	 => std_logic_vector(to_unsigned(43,8) ,
70578	 => std_logic_vector(to_unsigned(25,8) ,
70579	 => std_logic_vector(to_unsigned(15,8) ,
70580	 => std_logic_vector(to_unsigned(27,8) ,
70581	 => std_logic_vector(to_unsigned(19,8) ,
70582	 => std_logic_vector(to_unsigned(28,8) ,
70583	 => std_logic_vector(to_unsigned(37,8) ,
70584	 => std_logic_vector(to_unsigned(17,8) ,
70585	 => std_logic_vector(to_unsigned(15,8) ,
70586	 => std_logic_vector(to_unsigned(31,8) ,
70587	 => std_logic_vector(to_unsigned(25,8) ,
70588	 => std_logic_vector(to_unsigned(14,8) ,
70589	 => std_logic_vector(to_unsigned(14,8) ,
70590	 => std_logic_vector(to_unsigned(28,8) ,
70591	 => std_logic_vector(to_unsigned(37,8) ,
70592	 => std_logic_vector(to_unsigned(17,8) ,
70593	 => std_logic_vector(to_unsigned(12,8) ,
70594	 => std_logic_vector(to_unsigned(18,8) ,
70595	 => std_logic_vector(to_unsigned(32,8) ,
70596	 => std_logic_vector(to_unsigned(34,8) ,
70597	 => std_logic_vector(to_unsigned(40,8) ,
70598	 => std_logic_vector(to_unsigned(47,8) ,
70599	 => std_logic_vector(to_unsigned(32,8) ,
70600	 => std_logic_vector(to_unsigned(26,8) ,
70601	 => std_logic_vector(to_unsigned(20,8) ,
70602	 => std_logic_vector(to_unsigned(15,8) ,
70603	 => std_logic_vector(to_unsigned(18,8) ,
70604	 => std_logic_vector(to_unsigned(15,8) ,
70605	 => std_logic_vector(to_unsigned(17,8) ,
70606	 => std_logic_vector(to_unsigned(11,8) ,
70607	 => std_logic_vector(to_unsigned(10,8) ,
70608	 => std_logic_vector(to_unsigned(22,8) ,
70609	 => std_logic_vector(to_unsigned(43,8) ,
70610	 => std_logic_vector(to_unsigned(59,8) ,
70611	 => std_logic_vector(to_unsigned(38,8) ,
70612	 => std_logic_vector(to_unsigned(23,8) ,
70613	 => std_logic_vector(to_unsigned(24,8) ,
70614	 => std_logic_vector(to_unsigned(28,8) ,
70615	 => std_logic_vector(to_unsigned(37,8) ,
70616	 => std_logic_vector(to_unsigned(31,8) ,
70617	 => std_logic_vector(to_unsigned(21,8) ,
70618	 => std_logic_vector(to_unsigned(20,8) ,
70619	 => std_logic_vector(to_unsigned(23,8) ,
70620	 => std_logic_vector(to_unsigned(32,8) ,
70621	 => std_logic_vector(to_unsigned(28,8) ,
70622	 => std_logic_vector(to_unsigned(15,8) ,
70623	 => std_logic_vector(to_unsigned(24,8) ,
70624	 => std_logic_vector(to_unsigned(45,8) ,
70625	 => std_logic_vector(to_unsigned(37,8) ,
70626	 => std_logic_vector(to_unsigned(31,8) ,
70627	 => std_logic_vector(to_unsigned(24,8) ,
70628	 => std_logic_vector(to_unsigned(16,8) ,
70629	 => std_logic_vector(to_unsigned(4,8) ,
70630	 => std_logic_vector(to_unsigned(13,8) ,
70631	 => std_logic_vector(to_unsigned(29,8) ,
70632	 => std_logic_vector(to_unsigned(16,8) ,
70633	 => std_logic_vector(to_unsigned(29,8) ,
70634	 => std_logic_vector(to_unsigned(33,8) ,
70635	 => std_logic_vector(to_unsigned(50,8) ,
70636	 => std_logic_vector(to_unsigned(45,8) ,
70637	 => std_logic_vector(to_unsigned(41,8) ,
70638	 => std_logic_vector(to_unsigned(54,8) ,
70639	 => std_logic_vector(to_unsigned(59,8) ,
70640	 => std_logic_vector(to_unsigned(32,8) ,
70641	 => std_logic_vector(to_unsigned(19,8) ,
70642	 => std_logic_vector(to_unsigned(34,8) ,
70643	 => std_logic_vector(to_unsigned(65,8) ,
70644	 => std_logic_vector(to_unsigned(87,8) ,
70645	 => std_logic_vector(to_unsigned(100,8) ,
70646	 => std_logic_vector(to_unsigned(44,8) ,
70647	 => std_logic_vector(to_unsigned(70,8) ,
70648	 => std_logic_vector(to_unsigned(131,8) ,
70649	 => std_logic_vector(to_unsigned(107,8) ,
70650	 => std_logic_vector(to_unsigned(19,8) ,
70651	 => std_logic_vector(to_unsigned(8,8) ,
70652	 => std_logic_vector(to_unsigned(11,8) ,
70653	 => std_logic_vector(to_unsigned(7,8) ,
70654	 => std_logic_vector(to_unsigned(8,8) ,
70655	 => std_logic_vector(to_unsigned(7,8) ,
70656	 => std_logic_vector(to_unsigned(7,8) ,
70657	 => std_logic_vector(to_unsigned(7,8) ,
70658	 => std_logic_vector(to_unsigned(8,8) ,
70659	 => std_logic_vector(to_unsigned(6,8) ,
70660	 => std_logic_vector(to_unsigned(11,8) ,
70661	 => std_logic_vector(to_unsigned(18,8) ,
70662	 => std_logic_vector(to_unsigned(23,8) ,
70663	 => std_logic_vector(to_unsigned(26,8) ,
70664	 => std_logic_vector(to_unsigned(24,8) ,
70665	 => std_logic_vector(to_unsigned(27,8) ,
70666	 => std_logic_vector(to_unsigned(45,8) ,
70667	 => std_logic_vector(to_unsigned(41,8) ,
70668	 => std_logic_vector(to_unsigned(31,8) ,
70669	 => std_logic_vector(to_unsigned(24,8) ,
70670	 => std_logic_vector(to_unsigned(28,8) ,
70671	 => std_logic_vector(to_unsigned(11,8) ,
70672	 => std_logic_vector(to_unsigned(3,8) ,
70673	 => std_logic_vector(to_unsigned(5,8) ,
70674	 => std_logic_vector(to_unsigned(7,8) ,
70675	 => std_logic_vector(to_unsigned(6,8) ,
70676	 => std_logic_vector(to_unsigned(0,8) ,
70677	 => std_logic_vector(to_unsigned(1,8) ,
70678	 => std_logic_vector(to_unsigned(10,8) ,
70679	 => std_logic_vector(to_unsigned(10,8) ,
70680	 => std_logic_vector(to_unsigned(11,8) ,
70681	 => std_logic_vector(to_unsigned(11,8) ,
70682	 => std_logic_vector(to_unsigned(10,8) ,
70683	 => std_logic_vector(to_unsigned(6,8) ,
70684	 => std_logic_vector(to_unsigned(4,8) ,
70685	 => std_logic_vector(to_unsigned(12,8) ,
70686	 => std_logic_vector(to_unsigned(5,8) ,
70687	 => std_logic_vector(to_unsigned(1,8) ,
70688	 => std_logic_vector(to_unsigned(1,8) ,
70689	 => std_logic_vector(to_unsigned(0,8) ,
70690	 => std_logic_vector(to_unsigned(1,8) ,
70691	 => std_logic_vector(to_unsigned(1,8) ,
70692	 => std_logic_vector(to_unsigned(1,8) ,
70693	 => std_logic_vector(to_unsigned(0,8) ,
70694	 => std_logic_vector(to_unsigned(1,8) ,
70695	 => std_logic_vector(to_unsigned(1,8) ,
70696	 => std_logic_vector(to_unsigned(1,8) ,
70697	 => std_logic_vector(to_unsigned(3,8) ,
70698	 => std_logic_vector(to_unsigned(6,8) ,
70699	 => std_logic_vector(to_unsigned(4,8) ,
70700	 => std_logic_vector(to_unsigned(1,8) ,
70701	 => std_logic_vector(to_unsigned(0,8) ,
70702	 => std_logic_vector(to_unsigned(0,8) ,
70703	 => std_logic_vector(to_unsigned(0,8) ,
70704	 => std_logic_vector(to_unsigned(1,8) ,
70705	 => std_logic_vector(to_unsigned(49,8) ,
70706	 => std_logic_vector(to_unsigned(73,8) ,
70707	 => std_logic_vector(to_unsigned(95,8) ,
70708	 => std_logic_vector(to_unsigned(65,8) ,
70709	 => std_logic_vector(to_unsigned(21,8) ,
70710	 => std_logic_vector(to_unsigned(19,8) ,
70711	 => std_logic_vector(to_unsigned(44,8) ,
70712	 => std_logic_vector(to_unsigned(14,8) ,
70713	 => std_logic_vector(to_unsigned(38,8) ,
70714	 => std_logic_vector(to_unsigned(14,8) ,
70715	 => std_logic_vector(to_unsigned(12,8) ,
70716	 => std_logic_vector(to_unsigned(19,8) ,
70717	 => std_logic_vector(to_unsigned(11,8) ,
70718	 => std_logic_vector(to_unsigned(8,8) ,
70719	 => std_logic_vector(to_unsigned(9,8) ,
70720	 => std_logic_vector(to_unsigned(14,8) ,
70721	 => std_logic_vector(to_unsigned(116,8) ,
70722	 => std_logic_vector(to_unsigned(115,8) ,
70723	 => std_logic_vector(to_unsigned(114,8) ,
70724	 => std_logic_vector(to_unsigned(103,8) ,
70725	 => std_logic_vector(to_unsigned(84,8) ,
70726	 => std_logic_vector(to_unsigned(96,8) ,
70727	 => std_logic_vector(to_unsigned(116,8) ,
70728	 => std_logic_vector(to_unsigned(128,8) ,
70729	 => std_logic_vector(to_unsigned(130,8) ,
70730	 => std_logic_vector(to_unsigned(122,8) ,
70731	 => std_logic_vector(to_unsigned(90,8) ,
70732	 => std_logic_vector(to_unsigned(61,8) ,
70733	 => std_logic_vector(to_unsigned(50,8) ,
70734	 => std_logic_vector(to_unsigned(29,8) ,
70735	 => std_logic_vector(to_unsigned(35,8) ,
70736	 => std_logic_vector(to_unsigned(39,8) ,
70737	 => std_logic_vector(to_unsigned(55,8) ,
70738	 => std_logic_vector(to_unsigned(97,8) ,
70739	 => std_logic_vector(to_unsigned(108,8) ,
70740	 => std_logic_vector(to_unsigned(91,8) ,
70741	 => std_logic_vector(to_unsigned(62,8) ,
70742	 => std_logic_vector(to_unsigned(54,8) ,
70743	 => std_logic_vector(to_unsigned(46,8) ,
70744	 => std_logic_vector(to_unsigned(36,8) ,
70745	 => std_logic_vector(to_unsigned(27,8) ,
70746	 => std_logic_vector(to_unsigned(24,8) ,
70747	 => std_logic_vector(to_unsigned(25,8) ,
70748	 => std_logic_vector(to_unsigned(28,8) ,
70749	 => std_logic_vector(to_unsigned(29,8) ,
70750	 => std_logic_vector(to_unsigned(37,8) ,
70751	 => std_logic_vector(to_unsigned(37,8) ,
70752	 => std_logic_vector(to_unsigned(37,8) ,
70753	 => std_logic_vector(to_unsigned(56,8) ,
70754	 => std_logic_vector(to_unsigned(45,8) ,
70755	 => std_logic_vector(to_unsigned(47,8) ,
70756	 => std_logic_vector(to_unsigned(44,8) ,
70757	 => std_logic_vector(to_unsigned(46,8) ,
70758	 => std_logic_vector(to_unsigned(45,8) ,
70759	 => std_logic_vector(to_unsigned(18,8) ,
70760	 => std_logic_vector(to_unsigned(19,8) ,
70761	 => std_logic_vector(to_unsigned(24,8) ,
70762	 => std_logic_vector(to_unsigned(20,8) ,
70763	 => std_logic_vector(to_unsigned(23,8) ,
70764	 => std_logic_vector(to_unsigned(26,8) ,
70765	 => std_logic_vector(to_unsigned(23,8) ,
70766	 => std_logic_vector(to_unsigned(20,8) ,
70767	 => std_logic_vector(to_unsigned(20,8) ,
70768	 => std_logic_vector(to_unsigned(23,8) ,
70769	 => std_logic_vector(to_unsigned(26,8) ,
70770	 => std_logic_vector(to_unsigned(34,8) ,
70771	 => std_logic_vector(to_unsigned(37,8) ,
70772	 => std_logic_vector(to_unsigned(35,8) ,
70773	 => std_logic_vector(to_unsigned(33,8) ,
70774	 => std_logic_vector(to_unsigned(41,8) ,
70775	 => std_logic_vector(to_unsigned(39,8) ,
70776	 => std_logic_vector(to_unsigned(40,8) ,
70777	 => std_logic_vector(to_unsigned(42,8) ,
70778	 => std_logic_vector(to_unsigned(44,8) ,
70779	 => std_logic_vector(to_unsigned(45,8) ,
70780	 => std_logic_vector(to_unsigned(57,8) ,
70781	 => std_logic_vector(to_unsigned(54,8) ,
70782	 => std_logic_vector(to_unsigned(53,8) ,
70783	 => std_logic_vector(to_unsigned(53,8) ,
70784	 => std_logic_vector(to_unsigned(49,8) ,
70785	 => std_logic_vector(to_unsigned(46,8) ,
70786	 => std_logic_vector(to_unsigned(51,8) ,
70787	 => std_logic_vector(to_unsigned(41,8) ,
70788	 => std_logic_vector(to_unsigned(41,8) ,
70789	 => std_logic_vector(to_unsigned(41,8) ,
70790	 => std_logic_vector(to_unsigned(42,8) ,
70791	 => std_logic_vector(to_unsigned(42,8) ,
70792	 => std_logic_vector(to_unsigned(39,8) ,
70793	 => std_logic_vector(to_unsigned(45,8) ,
70794	 => std_logic_vector(to_unsigned(52,8) ,
70795	 => std_logic_vector(to_unsigned(51,8) ,
70796	 => std_logic_vector(to_unsigned(45,8) ,
70797	 => std_logic_vector(to_unsigned(54,8) ,
70798	 => std_logic_vector(to_unsigned(59,8) ,
70799	 => std_logic_vector(to_unsigned(66,8) ,
70800	 => std_logic_vector(to_unsigned(70,8) ,
70801	 => std_logic_vector(to_unsigned(82,8) ,
70802	 => std_logic_vector(to_unsigned(73,8) ,
70803	 => std_logic_vector(to_unsigned(79,8) ,
70804	 => std_logic_vector(to_unsigned(87,8) ,
70805	 => std_logic_vector(to_unsigned(84,8) ,
70806	 => std_logic_vector(to_unsigned(77,8) ,
70807	 => std_logic_vector(to_unsigned(52,8) ,
70808	 => std_logic_vector(to_unsigned(47,8) ,
70809	 => std_logic_vector(to_unsigned(31,8) ,
70810	 => std_logic_vector(to_unsigned(35,8) ,
70811	 => std_logic_vector(to_unsigned(54,8) ,
70812	 => std_logic_vector(to_unsigned(35,8) ,
70813	 => std_logic_vector(to_unsigned(28,8) ,
70814	 => std_logic_vector(to_unsigned(33,8) ,
70815	 => std_logic_vector(to_unsigned(36,8) ,
70816	 => std_logic_vector(to_unsigned(30,8) ,
70817	 => std_logic_vector(to_unsigned(29,8) ,
70818	 => std_logic_vector(to_unsigned(28,8) ,
70819	 => std_logic_vector(to_unsigned(27,8) ,
70820	 => std_logic_vector(to_unsigned(22,8) ,
70821	 => std_logic_vector(to_unsigned(18,8) ,
70822	 => std_logic_vector(to_unsigned(32,8) ,
70823	 => std_logic_vector(to_unsigned(22,8) ,
70824	 => std_logic_vector(to_unsigned(19,8) ,
70825	 => std_logic_vector(to_unsigned(25,8) ,
70826	 => std_logic_vector(to_unsigned(20,8) ,
70827	 => std_logic_vector(to_unsigned(45,8) ,
70828	 => std_logic_vector(to_unsigned(41,8) ,
70829	 => std_logic_vector(to_unsigned(19,8) ,
70830	 => std_logic_vector(to_unsigned(15,8) ,
70831	 => std_logic_vector(to_unsigned(34,8) ,
70832	 => std_logic_vector(to_unsigned(40,8) ,
70833	 => std_logic_vector(to_unsigned(39,8) ,
70834	 => std_logic_vector(to_unsigned(37,8) ,
70835	 => std_logic_vector(to_unsigned(43,8) ,
70836	 => std_logic_vector(to_unsigned(88,8) ,
70837	 => std_logic_vector(to_unsigned(119,8) ,
70838	 => std_logic_vector(to_unsigned(115,8) ,
70839	 => std_logic_vector(to_unsigned(115,8) ,
70840	 => std_logic_vector(to_unsigned(116,8) ,
70841	 => std_logic_vector(to_unsigned(122,8) ,
70842	 => std_logic_vector(to_unsigned(125,8) ,
70843	 => std_logic_vector(to_unsigned(116,8) ,
70844	 => std_logic_vector(to_unsigned(114,8) ,
70845	 => std_logic_vector(to_unsigned(105,8) ,
70846	 => std_logic_vector(to_unsigned(100,8) ,
70847	 => std_logic_vector(to_unsigned(96,8) ,
70848	 => std_logic_vector(to_unsigned(100,8) ,
70849	 => std_logic_vector(to_unsigned(104,8) ,
70850	 => std_logic_vector(to_unsigned(90,8) ,
70851	 => std_logic_vector(to_unsigned(74,8) ,
70852	 => std_logic_vector(to_unsigned(72,8) ,
70853	 => std_logic_vector(to_unsigned(81,8) ,
70854	 => std_logic_vector(to_unsigned(87,8) ,
70855	 => std_logic_vector(to_unsigned(96,8) ,
70856	 => std_logic_vector(to_unsigned(88,8) ,
70857	 => std_logic_vector(to_unsigned(49,8) ,
70858	 => std_logic_vector(to_unsigned(79,8) ,
70859	 => std_logic_vector(to_unsigned(104,8) ,
70860	 => std_logic_vector(to_unsigned(90,8) ,
70861	 => std_logic_vector(to_unsigned(96,8) ,
70862	 => std_logic_vector(to_unsigned(97,8) ,
70863	 => std_logic_vector(to_unsigned(97,8) ,
70864	 => std_logic_vector(to_unsigned(87,8) ,
70865	 => std_logic_vector(to_unsigned(87,8) ,
70866	 => std_logic_vector(to_unsigned(90,8) ,
70867	 => std_logic_vector(to_unsigned(88,8) ,
70868	 => std_logic_vector(to_unsigned(79,8) ,
70869	 => std_logic_vector(to_unsigned(77,8) ,
70870	 => std_logic_vector(to_unsigned(79,8) ,
70871	 => std_logic_vector(to_unsigned(77,8) ,
70872	 => std_logic_vector(to_unsigned(70,8) ,
70873	 => std_logic_vector(to_unsigned(59,8) ,
70874	 => std_logic_vector(to_unsigned(37,8) ,
70875	 => std_logic_vector(to_unsigned(20,8) ,
70876	 => std_logic_vector(to_unsigned(24,8) ,
70877	 => std_logic_vector(to_unsigned(12,8) ,
70878	 => std_logic_vector(to_unsigned(8,8) ,
70879	 => std_logic_vector(to_unsigned(12,8) ,
70880	 => std_logic_vector(to_unsigned(12,8) ,
70881	 => std_logic_vector(to_unsigned(13,8) ,
70882	 => std_logic_vector(to_unsigned(17,8) ,
70883	 => std_logic_vector(to_unsigned(58,8) ,
70884	 => std_logic_vector(to_unsigned(67,8) ,
70885	 => std_logic_vector(to_unsigned(55,8) ,
70886	 => std_logic_vector(to_unsigned(33,8) ,
70887	 => std_logic_vector(to_unsigned(6,8) ,
70888	 => std_logic_vector(to_unsigned(6,8) ,
70889	 => std_logic_vector(to_unsigned(15,8) ,
70890	 => std_logic_vector(to_unsigned(16,8) ,
70891	 => std_logic_vector(to_unsigned(24,8) ,
70892	 => std_logic_vector(to_unsigned(16,8) ,
70893	 => std_logic_vector(to_unsigned(17,8) ,
70894	 => std_logic_vector(to_unsigned(17,8) ,
70895	 => std_logic_vector(to_unsigned(14,8) ,
70896	 => std_logic_vector(to_unsigned(41,8) ,
70897	 => std_logic_vector(to_unsigned(24,8) ,
70898	 => std_logic_vector(to_unsigned(16,8) ,
70899	 => std_logic_vector(to_unsigned(21,8) ,
70900	 => std_logic_vector(to_unsigned(15,8) ,
70901	 => std_logic_vector(to_unsigned(19,8) ,
70902	 => std_logic_vector(to_unsigned(27,8) ,
70903	 => std_logic_vector(to_unsigned(45,8) ,
70904	 => std_logic_vector(to_unsigned(18,8) ,
70905	 => std_logic_vector(to_unsigned(6,8) ,
70906	 => std_logic_vector(to_unsigned(22,8) ,
70907	 => std_logic_vector(to_unsigned(41,8) ,
70908	 => std_logic_vector(to_unsigned(50,8) ,
70909	 => std_logic_vector(to_unsigned(36,8) ,
70910	 => std_logic_vector(to_unsigned(28,8) ,
70911	 => std_logic_vector(to_unsigned(30,8) ,
70912	 => std_logic_vector(to_unsigned(21,8) ,
70913	 => std_logic_vector(to_unsigned(12,8) ,
70914	 => std_logic_vector(to_unsigned(16,8) ,
70915	 => std_logic_vector(to_unsigned(36,8) ,
70916	 => std_logic_vector(to_unsigned(33,8) ,
70917	 => std_logic_vector(to_unsigned(42,8) ,
70918	 => std_logic_vector(to_unsigned(68,8) ,
70919	 => std_logic_vector(to_unsigned(45,8) ,
70920	 => std_logic_vector(to_unsigned(29,8) ,
70921	 => std_logic_vector(to_unsigned(22,8) ,
70922	 => std_logic_vector(to_unsigned(17,8) ,
70923	 => std_logic_vector(to_unsigned(12,8) ,
70924	 => std_logic_vector(to_unsigned(13,8) ,
70925	 => std_logic_vector(to_unsigned(15,8) ,
70926	 => std_logic_vector(to_unsigned(8,8) ,
70927	 => std_logic_vector(to_unsigned(9,8) ,
70928	 => std_logic_vector(to_unsigned(19,8) ,
70929	 => std_logic_vector(to_unsigned(51,8) ,
70930	 => std_logic_vector(to_unsigned(84,8) ,
70931	 => std_logic_vector(to_unsigned(59,8) ,
70932	 => std_logic_vector(to_unsigned(23,8) ,
70933	 => std_logic_vector(to_unsigned(22,8) ,
70934	 => std_logic_vector(to_unsigned(31,8) ,
70935	 => std_logic_vector(to_unsigned(35,8) ,
70936	 => std_logic_vector(to_unsigned(27,8) ,
70937	 => std_logic_vector(to_unsigned(23,8) ,
70938	 => std_logic_vector(to_unsigned(20,8) ,
70939	 => std_logic_vector(to_unsigned(18,8) ,
70940	 => std_logic_vector(to_unsigned(29,8) ,
70941	 => std_logic_vector(to_unsigned(33,8) ,
70942	 => std_logic_vector(to_unsigned(23,8) ,
70943	 => std_logic_vector(to_unsigned(23,8) ,
70944	 => std_logic_vector(to_unsigned(42,8) ,
70945	 => std_logic_vector(to_unsigned(39,8) ,
70946	 => std_logic_vector(to_unsigned(30,8) ,
70947	 => std_logic_vector(to_unsigned(32,8) ,
70948	 => std_logic_vector(to_unsigned(23,8) ,
70949	 => std_logic_vector(to_unsigned(5,8) ,
70950	 => std_logic_vector(to_unsigned(12,8) ,
70951	 => std_logic_vector(to_unsigned(35,8) ,
70952	 => std_logic_vector(to_unsigned(28,8) ,
70953	 => std_logic_vector(to_unsigned(27,8) ,
70954	 => std_logic_vector(to_unsigned(32,8) ,
70955	 => std_logic_vector(to_unsigned(45,8) ,
70956	 => std_logic_vector(to_unsigned(31,8) ,
70957	 => std_logic_vector(to_unsigned(25,8) ,
70958	 => std_logic_vector(to_unsigned(54,8) ,
70959	 => std_logic_vector(to_unsigned(63,8) ,
70960	 => std_logic_vector(to_unsigned(40,8) ,
70961	 => std_logic_vector(to_unsigned(29,8) ,
70962	 => std_logic_vector(to_unsigned(33,8) ,
70963	 => std_logic_vector(to_unsigned(71,8) ,
70964	 => std_logic_vector(to_unsigned(99,8) ,
70965	 => std_logic_vector(to_unsigned(105,8) ,
70966	 => std_logic_vector(to_unsigned(47,8) ,
70967	 => std_logic_vector(to_unsigned(72,8) ,
70968	 => std_logic_vector(to_unsigned(128,8) ,
70969	 => std_logic_vector(to_unsigned(99,8) ,
70970	 => std_logic_vector(to_unsigned(15,8) ,
70971	 => std_logic_vector(to_unsigned(8,8) ,
70972	 => std_logic_vector(to_unsigned(9,8) ,
70973	 => std_logic_vector(to_unsigned(6,8) ,
70974	 => std_logic_vector(to_unsigned(11,8) ,
70975	 => std_logic_vector(to_unsigned(7,8) ,
70976	 => std_logic_vector(to_unsigned(12,8) ,
70977	 => std_logic_vector(to_unsigned(10,8) ,
70978	 => std_logic_vector(to_unsigned(8,8) ,
70979	 => std_logic_vector(to_unsigned(9,8) ,
70980	 => std_logic_vector(to_unsigned(9,8) ,
70981	 => std_logic_vector(to_unsigned(9,8) ,
70982	 => std_logic_vector(to_unsigned(8,8) ,
70983	 => std_logic_vector(to_unsigned(8,8) ,
70984	 => std_logic_vector(to_unsigned(6,8) ,
70985	 => std_logic_vector(to_unsigned(8,8) ,
70986	 => std_logic_vector(to_unsigned(9,8) ,
70987	 => std_logic_vector(to_unsigned(10,8) ,
70988	 => std_logic_vector(to_unsigned(14,8) ,
70989	 => std_logic_vector(to_unsigned(24,8) ,
70990	 => std_logic_vector(to_unsigned(28,8) ,
70991	 => std_logic_vector(to_unsigned(10,8) ,
70992	 => std_logic_vector(to_unsigned(5,8) ,
70993	 => std_logic_vector(to_unsigned(4,8) ,
70994	 => std_logic_vector(to_unsigned(8,8) ,
70995	 => std_logic_vector(to_unsigned(14,8) ,
70996	 => std_logic_vector(to_unsigned(1,8) ,
70997	 => std_logic_vector(to_unsigned(0,8) ,
70998	 => std_logic_vector(to_unsigned(6,8) ,
70999	 => std_logic_vector(to_unsigned(13,8) ,
71000	 => std_logic_vector(to_unsigned(13,8) ,
71001	 => std_logic_vector(to_unsigned(14,8) ,
71002	 => std_logic_vector(to_unsigned(13,8) ,
71003	 => std_logic_vector(to_unsigned(6,8) ,
71004	 => std_logic_vector(to_unsigned(5,8) ,
71005	 => std_logic_vector(to_unsigned(13,8) ,
71006	 => std_logic_vector(to_unsigned(8,8) ,
71007	 => std_logic_vector(to_unsigned(1,8) ,
71008	 => std_logic_vector(to_unsigned(0,8) ,
71009	 => std_logic_vector(to_unsigned(0,8) ,
71010	 => std_logic_vector(to_unsigned(1,8) ,
71011	 => std_logic_vector(to_unsigned(1,8) ,
71012	 => std_logic_vector(to_unsigned(0,8) ,
71013	 => std_logic_vector(to_unsigned(0,8) ,
71014	 => std_logic_vector(to_unsigned(0,8) ,
71015	 => std_logic_vector(to_unsigned(0,8) ,
71016	 => std_logic_vector(to_unsigned(0,8) ,
71017	 => std_logic_vector(to_unsigned(0,8) ,
71018	 => std_logic_vector(to_unsigned(1,8) ,
71019	 => std_logic_vector(to_unsigned(2,8) ,
71020	 => std_logic_vector(to_unsigned(3,8) ,
71021	 => std_logic_vector(to_unsigned(1,8) ,
71022	 => std_logic_vector(to_unsigned(0,8) ,
71023	 => std_logic_vector(to_unsigned(0,8) ,
71024	 => std_logic_vector(to_unsigned(0,8) ,
71025	 => std_logic_vector(to_unsigned(19,8) ,
71026	 => std_logic_vector(to_unsigned(116,8) ,
71027	 => std_logic_vector(to_unsigned(142,8) ,
71028	 => std_logic_vector(to_unsigned(34,8) ,
71029	 => std_logic_vector(to_unsigned(13,8) ,
71030	 => std_logic_vector(to_unsigned(17,8) ,
71031	 => std_logic_vector(to_unsigned(22,8) ,
71032	 => std_logic_vector(to_unsigned(11,8) ,
71033	 => std_logic_vector(to_unsigned(29,8) ,
71034	 => std_logic_vector(to_unsigned(15,8) ,
71035	 => std_logic_vector(to_unsigned(35,8) ,
71036	 => std_logic_vector(to_unsigned(44,8) ,
71037	 => std_logic_vector(to_unsigned(24,8) ,
71038	 => std_logic_vector(to_unsigned(22,8) ,
71039	 => std_logic_vector(to_unsigned(12,8) ,
71040	 => std_logic_vector(to_unsigned(22,8) ,
71041	 => std_logic_vector(to_unsigned(118,8) ,
71042	 => std_logic_vector(to_unsigned(119,8) ,
71043	 => std_logic_vector(to_unsigned(122,8) ,
71044	 => std_logic_vector(to_unsigned(95,8) ,
71045	 => std_logic_vector(to_unsigned(80,8) ,
71046	 => std_logic_vector(to_unsigned(121,8) ,
71047	 => std_logic_vector(to_unsigned(133,8) ,
71048	 => std_logic_vector(to_unsigned(119,8) ,
71049	 => std_logic_vector(to_unsigned(112,8) ,
71050	 => std_logic_vector(to_unsigned(122,8) ,
71051	 => std_logic_vector(to_unsigned(93,8) ,
71052	 => std_logic_vector(to_unsigned(86,8) ,
71053	 => std_logic_vector(to_unsigned(84,8) ,
71054	 => std_logic_vector(to_unsigned(77,8) ,
71055	 => std_logic_vector(to_unsigned(57,8) ,
71056	 => std_logic_vector(to_unsigned(40,8) ,
71057	 => std_logic_vector(to_unsigned(49,8) ,
71058	 => std_logic_vector(to_unsigned(81,8) ,
71059	 => std_logic_vector(to_unsigned(87,8) ,
71060	 => std_logic_vector(to_unsigned(59,8) ,
71061	 => std_logic_vector(to_unsigned(57,8) ,
71062	 => std_logic_vector(to_unsigned(61,8) ,
71063	 => std_logic_vector(to_unsigned(55,8) ,
71064	 => std_logic_vector(to_unsigned(54,8) ,
71065	 => std_logic_vector(to_unsigned(45,8) ,
71066	 => std_logic_vector(to_unsigned(44,8) ,
71067	 => std_logic_vector(to_unsigned(47,8) ,
71068	 => std_logic_vector(to_unsigned(40,8) ,
71069	 => std_logic_vector(to_unsigned(34,8) ,
71070	 => std_logic_vector(to_unsigned(36,8) ,
71071	 => std_logic_vector(to_unsigned(37,8) ,
71072	 => std_logic_vector(to_unsigned(42,8) ,
71073	 => std_logic_vector(to_unsigned(45,8) ,
71074	 => std_logic_vector(to_unsigned(17,8) ,
71075	 => std_logic_vector(to_unsigned(18,8) ,
71076	 => std_logic_vector(to_unsigned(25,8) ,
71077	 => std_logic_vector(to_unsigned(42,8) ,
71078	 => std_logic_vector(to_unsigned(45,8) ,
71079	 => std_logic_vector(to_unsigned(23,8) ,
71080	 => std_logic_vector(to_unsigned(19,8) ,
71081	 => std_logic_vector(to_unsigned(24,8) ,
71082	 => std_logic_vector(to_unsigned(22,8) ,
71083	 => std_logic_vector(to_unsigned(25,8) ,
71084	 => std_logic_vector(to_unsigned(24,8) ,
71085	 => std_logic_vector(to_unsigned(20,8) ,
71086	 => std_logic_vector(to_unsigned(21,8) ,
71087	 => std_logic_vector(to_unsigned(21,8) ,
71088	 => std_logic_vector(to_unsigned(21,8) ,
71089	 => std_logic_vector(to_unsigned(25,8) ,
71090	 => std_logic_vector(to_unsigned(35,8) ,
71091	 => std_logic_vector(to_unsigned(37,8) ,
71092	 => std_logic_vector(to_unsigned(29,8) ,
71093	 => std_logic_vector(to_unsigned(29,8) ,
71094	 => std_logic_vector(to_unsigned(35,8) ,
71095	 => std_logic_vector(to_unsigned(40,8) ,
71096	 => std_logic_vector(to_unsigned(37,8) ,
71097	 => std_logic_vector(to_unsigned(43,8) ,
71098	 => std_logic_vector(to_unsigned(44,8) ,
71099	 => std_logic_vector(to_unsigned(43,8) ,
71100	 => std_logic_vector(to_unsigned(56,8) ,
71101	 => std_logic_vector(to_unsigned(53,8) ,
71102	 => std_logic_vector(to_unsigned(48,8) ,
71103	 => std_logic_vector(to_unsigned(48,8) ,
71104	 => std_logic_vector(to_unsigned(45,8) ,
71105	 => std_logic_vector(to_unsigned(46,8) ,
71106	 => std_logic_vector(to_unsigned(51,8) ,
71107	 => std_logic_vector(to_unsigned(42,8) ,
71108	 => std_logic_vector(to_unsigned(41,8) ,
71109	 => std_logic_vector(to_unsigned(35,8) ,
71110	 => std_logic_vector(to_unsigned(36,8) ,
71111	 => std_logic_vector(to_unsigned(41,8) ,
71112	 => std_logic_vector(to_unsigned(41,8) ,
71113	 => std_logic_vector(to_unsigned(46,8) ,
71114	 => std_logic_vector(to_unsigned(51,8) ,
71115	 => std_logic_vector(to_unsigned(52,8) ,
71116	 => std_logic_vector(to_unsigned(55,8) ,
71117	 => std_logic_vector(to_unsigned(56,8) ,
71118	 => std_logic_vector(to_unsigned(49,8) ,
71119	 => std_logic_vector(to_unsigned(53,8) ,
71120	 => std_logic_vector(to_unsigned(46,8) ,
71121	 => std_logic_vector(to_unsigned(65,8) ,
71122	 => std_logic_vector(to_unsigned(48,8) ,
71123	 => std_logic_vector(to_unsigned(72,8) ,
71124	 => std_logic_vector(to_unsigned(87,8) ,
71125	 => std_logic_vector(to_unsigned(82,8) ,
71126	 => std_logic_vector(to_unsigned(62,8) ,
71127	 => std_logic_vector(to_unsigned(29,8) ,
71128	 => std_logic_vector(to_unsigned(41,8) ,
71129	 => std_logic_vector(to_unsigned(34,8) ,
71130	 => std_logic_vector(to_unsigned(29,8) ,
71131	 => std_logic_vector(to_unsigned(35,8) ,
71132	 => std_logic_vector(to_unsigned(45,8) ,
71133	 => std_logic_vector(to_unsigned(52,8) ,
71134	 => std_logic_vector(to_unsigned(46,8) ,
71135	 => std_logic_vector(to_unsigned(52,8) ,
71136	 => std_logic_vector(to_unsigned(48,8) ,
71137	 => std_logic_vector(to_unsigned(49,8) ,
71138	 => std_logic_vector(to_unsigned(35,8) ,
71139	 => std_logic_vector(to_unsigned(32,8) ,
71140	 => std_logic_vector(to_unsigned(29,8) ,
71141	 => std_logic_vector(to_unsigned(23,8) ,
71142	 => std_logic_vector(to_unsigned(29,8) ,
71143	 => std_logic_vector(to_unsigned(30,8) ,
71144	 => std_logic_vector(to_unsigned(32,8) ,
71145	 => std_logic_vector(to_unsigned(35,8) ,
71146	 => std_logic_vector(to_unsigned(25,8) ,
71147	 => std_logic_vector(to_unsigned(21,8) ,
71148	 => std_logic_vector(to_unsigned(15,8) ,
71149	 => std_logic_vector(to_unsigned(14,8) ,
71150	 => std_logic_vector(to_unsigned(31,8) ,
71151	 => std_logic_vector(to_unsigned(67,8) ,
71152	 => std_logic_vector(to_unsigned(73,8) ,
71153	 => std_logic_vector(to_unsigned(54,8) ,
71154	 => std_logic_vector(to_unsigned(50,8) ,
71155	 => std_logic_vector(to_unsigned(49,8) ,
71156	 => std_logic_vector(to_unsigned(87,8) ,
71157	 => std_logic_vector(to_unsigned(125,8) ,
71158	 => std_logic_vector(to_unsigned(121,8) ,
71159	 => std_logic_vector(to_unsigned(119,8) ,
71160	 => std_logic_vector(to_unsigned(116,8) ,
71161	 => std_logic_vector(to_unsigned(122,8) ,
71162	 => std_logic_vector(to_unsigned(128,8) ,
71163	 => std_logic_vector(to_unsigned(118,8) ,
71164	 => std_logic_vector(to_unsigned(116,8) ,
71165	 => std_logic_vector(to_unsigned(109,8) ,
71166	 => std_logic_vector(to_unsigned(103,8) ,
71167	 => std_logic_vector(to_unsigned(99,8) ,
71168	 => std_logic_vector(to_unsigned(93,8) ,
71169	 => std_logic_vector(to_unsigned(97,8) ,
71170	 => std_logic_vector(to_unsigned(86,8) ,
71171	 => std_logic_vector(to_unsigned(51,8) ,
71172	 => std_logic_vector(to_unsigned(63,8) ,
71173	 => std_logic_vector(to_unsigned(80,8) ,
71174	 => std_logic_vector(to_unsigned(87,8) ,
71175	 => std_logic_vector(to_unsigned(93,8) ,
71176	 => std_logic_vector(to_unsigned(86,8) ,
71177	 => std_logic_vector(to_unsigned(74,8) ,
71178	 => std_logic_vector(to_unsigned(87,8) ,
71179	 => std_logic_vector(to_unsigned(97,8) ,
71180	 => std_logic_vector(to_unsigned(92,8) ,
71181	 => std_logic_vector(to_unsigned(93,8) ,
71182	 => std_logic_vector(to_unsigned(93,8) ,
71183	 => std_logic_vector(to_unsigned(91,8) ,
71184	 => std_logic_vector(to_unsigned(90,8) ,
71185	 => std_logic_vector(to_unsigned(86,8) ,
71186	 => std_logic_vector(to_unsigned(87,8) ,
71187	 => std_logic_vector(to_unsigned(85,8) ,
71188	 => std_logic_vector(to_unsigned(74,8) ,
71189	 => std_logic_vector(to_unsigned(74,8) ,
71190	 => std_logic_vector(to_unsigned(71,8) ,
71191	 => std_logic_vector(to_unsigned(66,8) ,
71192	 => std_logic_vector(to_unsigned(55,8) ,
71193	 => std_logic_vector(to_unsigned(51,8) ,
71194	 => std_logic_vector(to_unsigned(36,8) ,
71195	 => std_logic_vector(to_unsigned(17,8) ,
71196	 => std_logic_vector(to_unsigned(23,8) ,
71197	 => std_logic_vector(to_unsigned(10,8) ,
71198	 => std_logic_vector(to_unsigned(6,8) ,
71199	 => std_logic_vector(to_unsigned(7,8) ,
71200	 => std_logic_vector(to_unsigned(10,8) ,
71201	 => std_logic_vector(to_unsigned(17,8) ,
71202	 => std_logic_vector(to_unsigned(24,8) ,
71203	 => std_logic_vector(to_unsigned(45,8) ,
71204	 => std_logic_vector(to_unsigned(54,8) ,
71205	 => std_logic_vector(to_unsigned(50,8) ,
71206	 => std_logic_vector(to_unsigned(38,8) ,
71207	 => std_logic_vector(to_unsigned(5,8) ,
71208	 => std_logic_vector(to_unsigned(5,8) ,
71209	 => std_logic_vector(to_unsigned(13,8) ,
71210	 => std_logic_vector(to_unsigned(13,8) ,
71211	 => std_logic_vector(to_unsigned(15,8) ,
71212	 => std_logic_vector(to_unsigned(19,8) ,
71213	 => std_logic_vector(to_unsigned(24,8) ,
71214	 => std_logic_vector(to_unsigned(17,8) ,
71215	 => std_logic_vector(to_unsigned(34,8) ,
71216	 => std_logic_vector(to_unsigned(32,8) ,
71217	 => std_logic_vector(to_unsigned(17,8) ,
71218	 => std_logic_vector(to_unsigned(19,8) ,
71219	 => std_logic_vector(to_unsigned(14,8) ,
71220	 => std_logic_vector(to_unsigned(29,8) ,
71221	 => std_logic_vector(to_unsigned(24,8) ,
71222	 => std_logic_vector(to_unsigned(25,8) ,
71223	 => std_logic_vector(to_unsigned(23,8) ,
71224	 => std_logic_vector(to_unsigned(9,8) ,
71225	 => std_logic_vector(to_unsigned(9,8) ,
71226	 => std_logic_vector(to_unsigned(23,8) ,
71227	 => std_logic_vector(to_unsigned(41,8) ,
71228	 => std_logic_vector(to_unsigned(58,8) ,
71229	 => std_logic_vector(to_unsigned(44,8) ,
71230	 => std_logic_vector(to_unsigned(28,8) ,
71231	 => std_logic_vector(to_unsigned(30,8) ,
71232	 => std_logic_vector(to_unsigned(37,8) ,
71233	 => std_logic_vector(to_unsigned(38,8) ,
71234	 => std_logic_vector(to_unsigned(35,8) ,
71235	 => std_logic_vector(to_unsigned(34,8) ,
71236	 => std_logic_vector(to_unsigned(30,8) ,
71237	 => std_logic_vector(to_unsigned(41,8) ,
71238	 => std_logic_vector(to_unsigned(72,8) ,
71239	 => std_logic_vector(to_unsigned(70,8) ,
71240	 => std_logic_vector(to_unsigned(32,8) ,
71241	 => std_logic_vector(to_unsigned(32,8) ,
71242	 => std_logic_vector(to_unsigned(16,8) ,
71243	 => std_logic_vector(to_unsigned(8,8) ,
71244	 => std_logic_vector(to_unsigned(17,8) ,
71245	 => std_logic_vector(to_unsigned(17,8) ,
71246	 => std_logic_vector(to_unsigned(10,8) ,
71247	 => std_logic_vector(to_unsigned(9,8) ,
71248	 => std_logic_vector(to_unsigned(20,8) ,
71249	 => std_logic_vector(to_unsigned(36,8) ,
71250	 => std_logic_vector(to_unsigned(47,8) ,
71251	 => std_logic_vector(to_unsigned(41,8) ,
71252	 => std_logic_vector(to_unsigned(20,8) ,
71253	 => std_logic_vector(to_unsigned(20,8) ,
71254	 => std_logic_vector(to_unsigned(37,8) ,
71255	 => std_logic_vector(to_unsigned(49,8) ,
71256	 => std_logic_vector(to_unsigned(38,8) ,
71257	 => std_logic_vector(to_unsigned(21,8) ,
71258	 => std_logic_vector(to_unsigned(22,8) ,
71259	 => std_logic_vector(to_unsigned(27,8) ,
71260	 => std_logic_vector(to_unsigned(31,8) ,
71261	 => std_logic_vector(to_unsigned(25,8) ,
71262	 => std_logic_vector(to_unsigned(20,8) ,
71263	 => std_logic_vector(to_unsigned(27,8) ,
71264	 => std_logic_vector(to_unsigned(30,8) ,
71265	 => std_logic_vector(to_unsigned(29,8) ,
71266	 => std_logic_vector(to_unsigned(24,8) ,
71267	 => std_logic_vector(to_unsigned(29,8) ,
71268	 => std_logic_vector(to_unsigned(19,8) ,
71269	 => std_logic_vector(to_unsigned(5,8) ,
71270	 => std_logic_vector(to_unsigned(13,8) ,
71271	 => std_logic_vector(to_unsigned(20,8) ,
71272	 => std_logic_vector(to_unsigned(10,8) ,
71273	 => std_logic_vector(to_unsigned(21,8) ,
71274	 => std_logic_vector(to_unsigned(31,8) ,
71275	 => std_logic_vector(to_unsigned(47,8) ,
71276	 => std_logic_vector(to_unsigned(33,8) ,
71277	 => std_logic_vector(to_unsigned(31,8) ,
71278	 => std_logic_vector(to_unsigned(53,8) ,
71279	 => std_logic_vector(to_unsigned(59,8) ,
71280	 => std_logic_vector(to_unsigned(39,8) ,
71281	 => std_logic_vector(to_unsigned(36,8) ,
71282	 => std_logic_vector(to_unsigned(45,8) ,
71283	 => std_logic_vector(to_unsigned(78,8) ,
71284	 => std_logic_vector(to_unsigned(108,8) ,
71285	 => std_logic_vector(to_unsigned(104,8) ,
71286	 => std_logic_vector(to_unsigned(47,8) ,
71287	 => std_logic_vector(to_unsigned(78,8) ,
71288	 => std_logic_vector(to_unsigned(128,8) ,
71289	 => std_logic_vector(to_unsigned(105,8) ,
71290	 => std_logic_vector(to_unsigned(22,8) ,
71291	 => std_logic_vector(to_unsigned(8,8) ,
71292	 => std_logic_vector(to_unsigned(10,8) ,
71293	 => std_logic_vector(to_unsigned(8,8) ,
71294	 => std_logic_vector(to_unsigned(10,8) ,
71295	 => std_logic_vector(to_unsigned(12,8) ,
71296	 => std_logic_vector(to_unsigned(15,8) ,
71297	 => std_logic_vector(to_unsigned(11,8) ,
71298	 => std_logic_vector(to_unsigned(10,8) ,
71299	 => std_logic_vector(to_unsigned(13,8) ,
71300	 => std_logic_vector(to_unsigned(8,8) ,
71301	 => std_logic_vector(to_unsigned(10,8) ,
71302	 => std_logic_vector(to_unsigned(9,8) ,
71303	 => std_logic_vector(to_unsigned(10,8) ,
71304	 => std_logic_vector(to_unsigned(8,8) ,
71305	 => std_logic_vector(to_unsigned(8,8) ,
71306	 => std_logic_vector(to_unsigned(8,8) ,
71307	 => std_logic_vector(to_unsigned(8,8) ,
71308	 => std_logic_vector(to_unsigned(8,8) ,
71309	 => std_logic_vector(to_unsigned(25,8) ,
71310	 => std_logic_vector(to_unsigned(41,8) ,
71311	 => std_logic_vector(to_unsigned(25,8) ,
71312	 => std_logic_vector(to_unsigned(8,8) ,
71313	 => std_logic_vector(to_unsigned(16,8) ,
71314	 => std_logic_vector(to_unsigned(24,8) ,
71315	 => std_logic_vector(to_unsigned(23,8) ,
71316	 => std_logic_vector(to_unsigned(2,8) ,
71317	 => std_logic_vector(to_unsigned(0,8) ,
71318	 => std_logic_vector(to_unsigned(4,8) ,
71319	 => std_logic_vector(to_unsigned(12,8) ,
71320	 => std_logic_vector(to_unsigned(13,8) ,
71321	 => std_logic_vector(to_unsigned(12,8) ,
71322	 => std_logic_vector(to_unsigned(12,8) ,
71323	 => std_logic_vector(to_unsigned(4,8) ,
71324	 => std_logic_vector(to_unsigned(8,8) ,
71325	 => std_logic_vector(to_unsigned(17,8) ,
71326	 => std_logic_vector(to_unsigned(15,8) ,
71327	 => std_logic_vector(to_unsigned(4,8) ,
71328	 => std_logic_vector(to_unsigned(0,8) ,
71329	 => std_logic_vector(to_unsigned(0,8) ,
71330	 => std_logic_vector(to_unsigned(0,8) ,
71331	 => std_logic_vector(to_unsigned(0,8) ,
71332	 => std_logic_vector(to_unsigned(0,8) ,
71333	 => std_logic_vector(to_unsigned(0,8) ,
71334	 => std_logic_vector(to_unsigned(0,8) ,
71335	 => std_logic_vector(to_unsigned(0,8) ,
71336	 => std_logic_vector(to_unsigned(0,8) ,
71337	 => std_logic_vector(to_unsigned(1,8) ,
71338	 => std_logic_vector(to_unsigned(1,8) ,
71339	 => std_logic_vector(to_unsigned(0,8) ,
71340	 => std_logic_vector(to_unsigned(1,8) ,
71341	 => std_logic_vector(to_unsigned(1,8) ,
71342	 => std_logic_vector(to_unsigned(0,8) ,
71343	 => std_logic_vector(to_unsigned(0,8) ,
71344	 => std_logic_vector(to_unsigned(0,8) ,
71345	 => std_logic_vector(to_unsigned(7,8) ,
71346	 => std_logic_vector(to_unsigned(107,8) ,
71347	 => std_logic_vector(to_unsigned(115,8) ,
71348	 => std_logic_vector(to_unsigned(21,8) ,
71349	 => std_logic_vector(to_unsigned(10,8) ,
71350	 => std_logic_vector(to_unsigned(19,8) ,
71351	 => std_logic_vector(to_unsigned(22,8) ,
71352	 => std_logic_vector(to_unsigned(24,8) ,
71353	 => std_logic_vector(to_unsigned(21,8) ,
71354	 => std_logic_vector(to_unsigned(11,8) ,
71355	 => std_logic_vector(to_unsigned(14,8) ,
71356	 => std_logic_vector(to_unsigned(24,8) ,
71357	 => std_logic_vector(to_unsigned(41,8) ,
71358	 => std_logic_vector(to_unsigned(36,8) ,
71359	 => std_logic_vector(to_unsigned(17,8) ,
71360	 => std_logic_vector(to_unsigned(10,8) ,
71361	 => std_logic_vector(to_unsigned(125,8) ,
71362	 => std_logic_vector(to_unsigned(124,8) ,
71363	 => std_logic_vector(to_unsigned(122,8) ,
71364	 => std_logic_vector(to_unsigned(119,8) ,
71365	 => std_logic_vector(to_unsigned(125,8) ,
71366	 => std_logic_vector(to_unsigned(136,8) ,
71367	 => std_logic_vector(to_unsigned(141,8) ,
71368	 => std_logic_vector(to_unsigned(112,8) ,
71369	 => std_logic_vector(to_unsigned(74,8) ,
71370	 => std_logic_vector(to_unsigned(84,8) ,
71371	 => std_logic_vector(to_unsigned(88,8) ,
71372	 => std_logic_vector(to_unsigned(88,8) ,
71373	 => std_logic_vector(to_unsigned(78,8) ,
71374	 => std_logic_vector(to_unsigned(62,8) ,
71375	 => std_logic_vector(to_unsigned(57,8) ,
71376	 => std_logic_vector(to_unsigned(61,8) ,
71377	 => std_logic_vector(to_unsigned(68,8) ,
71378	 => std_logic_vector(to_unsigned(72,8) ,
71379	 => std_logic_vector(to_unsigned(69,8) ,
71380	 => std_logic_vector(to_unsigned(60,8) ,
71381	 => std_logic_vector(to_unsigned(58,8) ,
71382	 => std_logic_vector(to_unsigned(51,8) ,
71383	 => std_logic_vector(to_unsigned(46,8) ,
71384	 => std_logic_vector(to_unsigned(48,8) ,
71385	 => std_logic_vector(to_unsigned(46,8) ,
71386	 => std_logic_vector(to_unsigned(47,8) ,
71387	 => std_logic_vector(to_unsigned(48,8) ,
71388	 => std_logic_vector(to_unsigned(51,8) ,
71389	 => std_logic_vector(to_unsigned(51,8) ,
71390	 => std_logic_vector(to_unsigned(49,8) ,
71391	 => std_logic_vector(to_unsigned(37,8) ,
71392	 => std_logic_vector(to_unsigned(39,8) ,
71393	 => std_logic_vector(to_unsigned(59,8) ,
71394	 => std_logic_vector(to_unsigned(30,8) ,
71395	 => std_logic_vector(to_unsigned(25,8) ,
71396	 => std_logic_vector(to_unsigned(20,8) ,
71397	 => std_logic_vector(to_unsigned(16,8) ,
71398	 => std_logic_vector(to_unsigned(31,8) ,
71399	 => std_logic_vector(to_unsigned(22,8) ,
71400	 => std_logic_vector(to_unsigned(20,8) ,
71401	 => std_logic_vector(to_unsigned(27,8) ,
71402	 => std_logic_vector(to_unsigned(29,8) ,
71403	 => std_logic_vector(to_unsigned(28,8) ,
71404	 => std_logic_vector(to_unsigned(23,8) ,
71405	 => std_logic_vector(to_unsigned(23,8) ,
71406	 => std_logic_vector(to_unsigned(29,8) ,
71407	 => std_logic_vector(to_unsigned(23,8) ,
71408	 => std_logic_vector(to_unsigned(23,8) ,
71409	 => std_logic_vector(to_unsigned(24,8) ,
71410	 => std_logic_vector(to_unsigned(33,8) ,
71411	 => std_logic_vector(to_unsigned(35,8) ,
71412	 => std_logic_vector(to_unsigned(26,8) ,
71413	 => std_logic_vector(to_unsigned(27,8) ,
71414	 => std_logic_vector(to_unsigned(35,8) ,
71415	 => std_logic_vector(to_unsigned(41,8) ,
71416	 => std_logic_vector(to_unsigned(36,8) ,
71417	 => std_logic_vector(to_unsigned(44,8) ,
71418	 => std_logic_vector(to_unsigned(40,8) ,
71419	 => std_logic_vector(to_unsigned(46,8) ,
71420	 => std_logic_vector(to_unsigned(52,8) ,
71421	 => std_logic_vector(to_unsigned(54,8) ,
71422	 => std_logic_vector(to_unsigned(53,8) ,
71423	 => std_logic_vector(to_unsigned(46,8) ,
71424	 => std_logic_vector(to_unsigned(50,8) ,
71425	 => std_logic_vector(to_unsigned(51,8) ,
71426	 => std_logic_vector(to_unsigned(45,8) ,
71427	 => std_logic_vector(to_unsigned(45,8) ,
71428	 => std_logic_vector(to_unsigned(44,8) ,
71429	 => std_logic_vector(to_unsigned(45,8) ,
71430	 => std_logic_vector(to_unsigned(44,8) ,
71431	 => std_logic_vector(to_unsigned(38,8) ,
71432	 => std_logic_vector(to_unsigned(43,8) ,
71433	 => std_logic_vector(to_unsigned(51,8) ,
71434	 => std_logic_vector(to_unsigned(59,8) ,
71435	 => std_logic_vector(to_unsigned(56,8) ,
71436	 => std_logic_vector(to_unsigned(53,8) ,
71437	 => std_logic_vector(to_unsigned(58,8) ,
71438	 => std_logic_vector(to_unsigned(48,8) ,
71439	 => std_logic_vector(to_unsigned(47,8) ,
71440	 => std_logic_vector(to_unsigned(43,8) ,
71441	 => std_logic_vector(to_unsigned(67,8) ,
71442	 => std_logic_vector(to_unsigned(43,8) ,
71443	 => std_logic_vector(to_unsigned(63,8) ,
71444	 => std_logic_vector(to_unsigned(85,8) ,
71445	 => std_logic_vector(to_unsigned(77,8) ,
71446	 => std_logic_vector(to_unsigned(45,8) ,
71447	 => std_logic_vector(to_unsigned(28,8) ,
71448	 => std_logic_vector(to_unsigned(33,8) ,
71449	 => std_logic_vector(to_unsigned(28,8) ,
71450	 => std_logic_vector(to_unsigned(31,8) ,
71451	 => std_logic_vector(to_unsigned(41,8) ,
71452	 => std_logic_vector(to_unsigned(51,8) ,
71453	 => std_logic_vector(to_unsigned(51,8) ,
71454	 => std_logic_vector(to_unsigned(33,8) ,
71455	 => std_logic_vector(to_unsigned(37,8) ,
71456	 => std_logic_vector(to_unsigned(54,8) ,
71457	 => std_logic_vector(to_unsigned(43,8) ,
71458	 => std_logic_vector(to_unsigned(46,8) ,
71459	 => std_logic_vector(to_unsigned(54,8) ,
71460	 => std_logic_vector(to_unsigned(47,8) ,
71461	 => std_logic_vector(to_unsigned(41,8) ,
71462	 => std_logic_vector(to_unsigned(41,8) ,
71463	 => std_logic_vector(to_unsigned(41,8) ,
71464	 => std_logic_vector(to_unsigned(37,8) ,
71465	 => std_logic_vector(to_unsigned(29,8) ,
71466	 => std_logic_vector(to_unsigned(22,8) ,
71467	 => std_logic_vector(to_unsigned(30,8) ,
71468	 => std_logic_vector(to_unsigned(29,8) ,
71469	 => std_logic_vector(to_unsigned(32,8) ,
71470	 => std_logic_vector(to_unsigned(61,8) ,
71471	 => std_logic_vector(to_unsigned(69,8) ,
71472	 => std_logic_vector(to_unsigned(69,8) ,
71473	 => std_logic_vector(to_unsigned(70,8) ,
71474	 => std_logic_vector(to_unsigned(59,8) ,
71475	 => std_logic_vector(to_unsigned(41,8) ,
71476	 => std_logic_vector(to_unsigned(90,8) ,
71477	 => std_logic_vector(to_unsigned(131,8) ,
71478	 => std_logic_vector(to_unsigned(118,8) ,
71479	 => std_logic_vector(to_unsigned(127,8) ,
71480	 => std_logic_vector(to_unsigned(125,8) ,
71481	 => std_logic_vector(to_unsigned(121,8) ,
71482	 => std_logic_vector(to_unsigned(122,8) ,
71483	 => std_logic_vector(to_unsigned(115,8) ,
71484	 => std_logic_vector(to_unsigned(119,8) ,
71485	 => std_logic_vector(to_unsigned(111,8) ,
71486	 => std_logic_vector(to_unsigned(105,8) ,
71487	 => std_logic_vector(to_unsigned(101,8) ,
71488	 => std_logic_vector(to_unsigned(91,8) ,
71489	 => std_logic_vector(to_unsigned(93,8) ,
71490	 => std_logic_vector(to_unsigned(78,8) ,
71491	 => std_logic_vector(to_unsigned(33,8) ,
71492	 => std_logic_vector(to_unsigned(36,8) ,
71493	 => std_logic_vector(to_unsigned(54,8) ,
71494	 => std_logic_vector(to_unsigned(57,8) ,
71495	 => std_logic_vector(to_unsigned(50,8) ,
71496	 => std_logic_vector(to_unsigned(71,8) ,
71497	 => std_logic_vector(to_unsigned(84,8) ,
71498	 => std_logic_vector(to_unsigned(82,8) ,
71499	 => std_logic_vector(to_unsigned(90,8) ,
71500	 => std_logic_vector(to_unsigned(87,8) ,
71501	 => std_logic_vector(to_unsigned(90,8) ,
71502	 => std_logic_vector(to_unsigned(97,8) ,
71503	 => std_logic_vector(to_unsigned(95,8) ,
71504	 => std_logic_vector(to_unsigned(93,8) ,
71505	 => std_logic_vector(to_unsigned(88,8) ,
71506	 => std_logic_vector(to_unsigned(82,8) ,
71507	 => std_logic_vector(to_unsigned(73,8) ,
71508	 => std_logic_vector(to_unsigned(65,8) ,
71509	 => std_logic_vector(to_unsigned(65,8) ,
71510	 => std_logic_vector(to_unsigned(60,8) ,
71511	 => std_logic_vector(to_unsigned(51,8) ,
71512	 => std_logic_vector(to_unsigned(45,8) ,
71513	 => std_logic_vector(to_unsigned(47,8) ,
71514	 => std_logic_vector(to_unsigned(35,8) ,
71515	 => std_logic_vector(to_unsigned(16,8) ,
71516	 => std_logic_vector(to_unsigned(17,8) ,
71517	 => std_logic_vector(to_unsigned(9,8) ,
71518	 => std_logic_vector(to_unsigned(19,8) ,
71519	 => std_logic_vector(to_unsigned(31,8) ,
71520	 => std_logic_vector(to_unsigned(11,8) ,
71521	 => std_logic_vector(to_unsigned(12,8) ,
71522	 => std_logic_vector(to_unsigned(16,8) ,
71523	 => std_logic_vector(to_unsigned(45,8) ,
71524	 => std_logic_vector(to_unsigned(62,8) ,
71525	 => std_logic_vector(to_unsigned(61,8) ,
71526	 => std_logic_vector(to_unsigned(35,8) ,
71527	 => std_logic_vector(to_unsigned(4,8) ,
71528	 => std_logic_vector(to_unsigned(6,8) ,
71529	 => std_logic_vector(to_unsigned(13,8) ,
71530	 => std_logic_vector(to_unsigned(11,8) ,
71531	 => std_logic_vector(to_unsigned(20,8) ,
71532	 => std_logic_vector(to_unsigned(28,8) ,
71533	 => std_logic_vector(to_unsigned(12,8) ,
71534	 => std_logic_vector(to_unsigned(36,8) ,
71535	 => std_logic_vector(to_unsigned(33,8) ,
71536	 => std_logic_vector(to_unsigned(12,8) ,
71537	 => std_logic_vector(to_unsigned(20,8) ,
71538	 => std_logic_vector(to_unsigned(13,8) ,
71539	 => std_logic_vector(to_unsigned(21,8) ,
71540	 => std_logic_vector(to_unsigned(40,8) ,
71541	 => std_logic_vector(to_unsigned(27,8) ,
71542	 => std_logic_vector(to_unsigned(44,8) ,
71543	 => std_logic_vector(to_unsigned(46,8) ,
71544	 => std_logic_vector(to_unsigned(32,8) ,
71545	 => std_logic_vector(to_unsigned(27,8) ,
71546	 => std_logic_vector(to_unsigned(26,8) ,
71547	 => std_logic_vector(to_unsigned(41,8) ,
71548	 => std_logic_vector(to_unsigned(62,8) ,
71549	 => std_logic_vector(to_unsigned(58,8) ,
71550	 => std_logic_vector(to_unsigned(29,8) ,
71551	 => std_logic_vector(to_unsigned(29,8) ,
71552	 => std_logic_vector(to_unsigned(39,8) ,
71553	 => std_logic_vector(to_unsigned(49,8) ,
71554	 => std_logic_vector(to_unsigned(38,8) ,
71555	 => std_logic_vector(to_unsigned(31,8) ,
71556	 => std_logic_vector(to_unsigned(28,8) ,
71557	 => std_logic_vector(to_unsigned(30,8) ,
71558	 => std_logic_vector(to_unsigned(40,8) ,
71559	 => std_logic_vector(to_unsigned(41,8) ,
71560	 => std_logic_vector(to_unsigned(30,8) ,
71561	 => std_logic_vector(to_unsigned(22,8) ,
71562	 => std_logic_vector(to_unsigned(11,8) ,
71563	 => std_logic_vector(to_unsigned(12,8) ,
71564	 => std_logic_vector(to_unsigned(15,8) ,
71565	 => std_logic_vector(to_unsigned(22,8) ,
71566	 => std_logic_vector(to_unsigned(13,8) ,
71567	 => std_logic_vector(to_unsigned(9,8) ,
71568	 => std_logic_vector(to_unsigned(18,8) ,
71569	 => std_logic_vector(to_unsigned(33,8) ,
71570	 => std_logic_vector(to_unsigned(52,8) ,
71571	 => std_logic_vector(to_unsigned(37,8) ,
71572	 => std_logic_vector(to_unsigned(20,8) ,
71573	 => std_logic_vector(to_unsigned(24,8) ,
71574	 => std_logic_vector(to_unsigned(20,8) ,
71575	 => std_logic_vector(to_unsigned(22,8) ,
71576	 => std_logic_vector(to_unsigned(29,8) ,
71577	 => std_logic_vector(to_unsigned(20,8) ,
71578	 => std_logic_vector(to_unsigned(19,8) ,
71579	 => std_logic_vector(to_unsigned(26,8) ,
71580	 => std_logic_vector(to_unsigned(36,8) ,
71581	 => std_logic_vector(to_unsigned(38,8) ,
71582	 => std_logic_vector(to_unsigned(15,8) ,
71583	 => std_logic_vector(to_unsigned(22,8) ,
71584	 => std_logic_vector(to_unsigned(33,8) ,
71585	 => std_logic_vector(to_unsigned(29,8) ,
71586	 => std_logic_vector(to_unsigned(26,8) ,
71587	 => std_logic_vector(to_unsigned(20,8) ,
71588	 => std_logic_vector(to_unsigned(11,8) ,
71589	 => std_logic_vector(to_unsigned(3,8) ,
71590	 => std_logic_vector(to_unsigned(13,8) ,
71591	 => std_logic_vector(to_unsigned(13,8) ,
71592	 => std_logic_vector(to_unsigned(5,8) ,
71593	 => std_logic_vector(to_unsigned(22,8) ,
71594	 => std_logic_vector(to_unsigned(39,8) ,
71595	 => std_logic_vector(to_unsigned(41,8) ,
71596	 => std_logic_vector(to_unsigned(10,8) ,
71597	 => std_logic_vector(to_unsigned(13,8) ,
71598	 => std_logic_vector(to_unsigned(51,8) ,
71599	 => std_logic_vector(to_unsigned(53,8) ,
71600	 => std_logic_vector(to_unsigned(19,8) ,
71601	 => std_logic_vector(to_unsigned(10,8) ,
71602	 => std_logic_vector(to_unsigned(33,8) ,
71603	 => std_logic_vector(to_unsigned(73,8) ,
71604	 => std_logic_vector(to_unsigned(104,8) ,
71605	 => std_logic_vector(to_unsigned(96,8) ,
71606	 => std_logic_vector(to_unsigned(45,8) ,
71607	 => std_logic_vector(to_unsigned(79,8) ,
71608	 => std_logic_vector(to_unsigned(128,8) ,
71609	 => std_logic_vector(to_unsigned(87,8) ,
71610	 => std_logic_vector(to_unsigned(13,8) ,
71611	 => std_logic_vector(to_unsigned(7,8) ,
71612	 => std_logic_vector(to_unsigned(9,8) ,
71613	 => std_logic_vector(to_unsigned(6,8) ,
71614	 => std_logic_vector(to_unsigned(9,8) ,
71615	 => std_logic_vector(to_unsigned(9,8) ,
71616	 => std_logic_vector(to_unsigned(9,8) ,
71617	 => std_logic_vector(to_unsigned(11,8) ,
71618	 => std_logic_vector(to_unsigned(12,8) ,
71619	 => std_logic_vector(to_unsigned(13,8) ,
71620	 => std_logic_vector(to_unsigned(11,8) ,
71621	 => std_logic_vector(to_unsigned(9,8) ,
71622	 => std_logic_vector(to_unsigned(7,8) ,
71623	 => std_logic_vector(to_unsigned(7,8) ,
71624	 => std_logic_vector(to_unsigned(12,8) ,
71625	 => std_logic_vector(to_unsigned(11,8) ,
71626	 => std_logic_vector(to_unsigned(9,8) ,
71627	 => std_logic_vector(to_unsigned(10,8) ,
71628	 => std_logic_vector(to_unsigned(12,8) ,
71629	 => std_logic_vector(to_unsigned(30,8) ,
71630	 => std_logic_vector(to_unsigned(35,8) ,
71631	 => std_logic_vector(to_unsigned(44,8) ,
71632	 => std_logic_vector(to_unsigned(27,8) ,
71633	 => std_logic_vector(to_unsigned(16,8) ,
71634	 => std_logic_vector(to_unsigned(17,8) ,
71635	 => std_logic_vector(to_unsigned(18,8) ,
71636	 => std_logic_vector(to_unsigned(5,8) ,
71637	 => std_logic_vector(to_unsigned(0,8) ,
71638	 => std_logic_vector(to_unsigned(2,8) ,
71639	 => std_logic_vector(to_unsigned(13,8) ,
71640	 => std_logic_vector(to_unsigned(13,8) ,
71641	 => std_logic_vector(to_unsigned(11,8) ,
71642	 => std_logic_vector(to_unsigned(9,8) ,
71643	 => std_logic_vector(to_unsigned(3,8) ,
71644	 => std_logic_vector(to_unsigned(8,8) ,
71645	 => std_logic_vector(to_unsigned(16,8) ,
71646	 => std_logic_vector(to_unsigned(15,8) ,
71647	 => std_logic_vector(to_unsigned(9,8) ,
71648	 => std_logic_vector(to_unsigned(1,8) ,
71649	 => std_logic_vector(to_unsigned(0,8) ,
71650	 => std_logic_vector(to_unsigned(0,8) ,
71651	 => std_logic_vector(to_unsigned(0,8) ,
71652	 => std_logic_vector(to_unsigned(0,8) ,
71653	 => std_logic_vector(to_unsigned(0,8) ,
71654	 => std_logic_vector(to_unsigned(2,8) ,
71655	 => std_logic_vector(to_unsigned(2,8) ,
71656	 => std_logic_vector(to_unsigned(1,8) ,
71657	 => std_logic_vector(to_unsigned(0,8) ,
71658	 => std_logic_vector(to_unsigned(1,8) ,
71659	 => std_logic_vector(to_unsigned(1,8) ,
71660	 => std_logic_vector(to_unsigned(1,8) ,
71661	 => std_logic_vector(to_unsigned(1,8) ,
71662	 => std_logic_vector(to_unsigned(1,8) ,
71663	 => std_logic_vector(to_unsigned(1,8) ,
71664	 => std_logic_vector(to_unsigned(0,8) ,
71665	 => std_logic_vector(to_unsigned(3,8) ,
71666	 => std_logic_vector(to_unsigned(52,8) ,
71667	 => std_logic_vector(to_unsigned(56,8) ,
71668	 => std_logic_vector(to_unsigned(41,8) ,
71669	 => std_logic_vector(to_unsigned(32,8) ,
71670	 => std_logic_vector(to_unsigned(68,8) ,
71671	 => std_logic_vector(to_unsigned(78,8) ,
71672	 => std_logic_vector(to_unsigned(59,8) ,
71673	 => std_logic_vector(to_unsigned(29,8) ,
71674	 => std_logic_vector(to_unsigned(15,8) ,
71675	 => std_logic_vector(to_unsigned(9,8) ,
71676	 => std_logic_vector(to_unsigned(26,8) ,
71677	 => std_logic_vector(to_unsigned(61,8) ,
71678	 => std_logic_vector(to_unsigned(51,8) ,
71679	 => std_logic_vector(to_unsigned(45,8) ,
71680	 => std_logic_vector(to_unsigned(14,8) ,
71681	 => std_logic_vector(to_unsigned(121,8) ,
71682	 => std_logic_vector(to_unsigned(125,8) ,
71683	 => std_logic_vector(to_unsigned(136,8) ,
71684	 => std_logic_vector(to_unsigned(142,8) ,
71685	 => std_logic_vector(to_unsigned(149,8) ,
71686	 => std_logic_vector(to_unsigned(136,8) ,
71687	 => std_logic_vector(to_unsigned(130,8) ,
71688	 => std_logic_vector(to_unsigned(100,8) ,
71689	 => std_logic_vector(to_unsigned(87,8) ,
71690	 => std_logic_vector(to_unsigned(97,8) ,
71691	 => std_logic_vector(to_unsigned(91,8) ,
71692	 => std_logic_vector(to_unsigned(68,8) ,
71693	 => std_logic_vector(to_unsigned(63,8) ,
71694	 => std_logic_vector(to_unsigned(61,8) ,
71695	 => std_logic_vector(to_unsigned(70,8) ,
71696	 => std_logic_vector(to_unsigned(80,8) ,
71697	 => std_logic_vector(to_unsigned(79,8) ,
71698	 => std_logic_vector(to_unsigned(81,8) ,
71699	 => std_logic_vector(to_unsigned(74,8) ,
71700	 => std_logic_vector(to_unsigned(67,8) ,
71701	 => std_logic_vector(to_unsigned(60,8) ,
71702	 => std_logic_vector(to_unsigned(55,8) ,
71703	 => std_logic_vector(to_unsigned(51,8) ,
71704	 => std_logic_vector(to_unsigned(47,8) ,
71705	 => std_logic_vector(to_unsigned(45,8) ,
71706	 => std_logic_vector(to_unsigned(48,8) ,
71707	 => std_logic_vector(to_unsigned(47,8) ,
71708	 => std_logic_vector(to_unsigned(39,8) ,
71709	 => std_logic_vector(to_unsigned(44,8) ,
71710	 => std_logic_vector(to_unsigned(51,8) ,
71711	 => std_logic_vector(to_unsigned(36,8) ,
71712	 => std_logic_vector(to_unsigned(37,8) ,
71713	 => std_logic_vector(to_unsigned(69,8) ,
71714	 => std_logic_vector(to_unsigned(92,8) ,
71715	 => std_logic_vector(to_unsigned(99,8) ,
71716	 => std_logic_vector(to_unsigned(81,8) ,
71717	 => std_logic_vector(to_unsigned(51,8) ,
71718	 => std_logic_vector(to_unsigned(47,8) ,
71719	 => std_logic_vector(to_unsigned(21,8) ,
71720	 => std_logic_vector(to_unsigned(19,8) ,
71721	 => std_logic_vector(to_unsigned(23,8) ,
71722	 => std_logic_vector(to_unsigned(24,8) ,
71723	 => std_logic_vector(to_unsigned(25,8) ,
71724	 => std_logic_vector(to_unsigned(27,8) ,
71725	 => std_logic_vector(to_unsigned(29,8) ,
71726	 => std_logic_vector(to_unsigned(26,8) ,
71727	 => std_logic_vector(to_unsigned(25,8) ,
71728	 => std_logic_vector(to_unsigned(29,8) ,
71729	 => std_logic_vector(to_unsigned(28,8) ,
71730	 => std_logic_vector(to_unsigned(29,8) ,
71731	 => std_logic_vector(to_unsigned(37,8) ,
71732	 => std_logic_vector(to_unsigned(36,8) ,
71733	 => std_logic_vector(to_unsigned(34,8) ,
71734	 => std_logic_vector(to_unsigned(38,8) ,
71735	 => std_logic_vector(to_unsigned(40,8) ,
71736	 => std_logic_vector(to_unsigned(41,8) ,
71737	 => std_logic_vector(to_unsigned(47,8) ,
71738	 => std_logic_vector(to_unsigned(44,8) ,
71739	 => std_logic_vector(to_unsigned(46,8) ,
71740	 => std_logic_vector(to_unsigned(51,8) ,
71741	 => std_logic_vector(to_unsigned(55,8) ,
71742	 => std_logic_vector(to_unsigned(55,8) ,
71743	 => std_logic_vector(to_unsigned(49,8) ,
71744	 => std_logic_vector(to_unsigned(44,8) ,
71745	 => std_logic_vector(to_unsigned(41,8) ,
71746	 => std_logic_vector(to_unsigned(45,8) ,
71747	 => std_logic_vector(to_unsigned(45,8) ,
71748	 => std_logic_vector(to_unsigned(43,8) ,
71749	 => std_logic_vector(to_unsigned(51,8) ,
71750	 => std_logic_vector(to_unsigned(51,8) ,
71751	 => std_logic_vector(to_unsigned(45,8) ,
71752	 => std_logic_vector(to_unsigned(44,8) ,
71753	 => std_logic_vector(to_unsigned(51,8) ,
71754	 => std_logic_vector(to_unsigned(61,8) ,
71755	 => std_logic_vector(to_unsigned(58,8) ,
71756	 => std_logic_vector(to_unsigned(59,8) ,
71757	 => std_logic_vector(to_unsigned(58,8) ,
71758	 => std_logic_vector(to_unsigned(48,8) ,
71759	 => std_logic_vector(to_unsigned(52,8) ,
71760	 => std_logic_vector(to_unsigned(45,8) ,
71761	 => std_logic_vector(to_unsigned(62,8) ,
71762	 => std_logic_vector(to_unsigned(45,8) ,
71763	 => std_logic_vector(to_unsigned(80,8) ,
71764	 => std_logic_vector(to_unsigned(91,8) ,
71765	 => std_logic_vector(to_unsigned(60,8) ,
71766	 => std_logic_vector(to_unsigned(54,8) ,
71767	 => std_logic_vector(to_unsigned(56,8) ,
71768	 => std_logic_vector(to_unsigned(54,8) ,
71769	 => std_logic_vector(to_unsigned(46,8) ,
71770	 => std_logic_vector(to_unsigned(55,8) ,
71771	 => std_logic_vector(to_unsigned(52,8) ,
71772	 => std_logic_vector(to_unsigned(39,8) ,
71773	 => std_logic_vector(to_unsigned(38,8) ,
71774	 => std_logic_vector(to_unsigned(25,8) ,
71775	 => std_logic_vector(to_unsigned(30,8) ,
71776	 => std_logic_vector(to_unsigned(52,8) ,
71777	 => std_logic_vector(to_unsigned(50,8) ,
71778	 => std_logic_vector(to_unsigned(62,8) ,
71779	 => std_logic_vector(to_unsigned(52,8) ,
71780	 => std_logic_vector(to_unsigned(37,8) ,
71781	 => std_logic_vector(to_unsigned(40,8) ,
71782	 => std_logic_vector(to_unsigned(41,8) ,
71783	 => std_logic_vector(to_unsigned(33,8) ,
71784	 => std_logic_vector(to_unsigned(33,8) ,
71785	 => std_logic_vector(to_unsigned(39,8) ,
71786	 => std_logic_vector(to_unsigned(43,8) ,
71787	 => std_logic_vector(to_unsigned(52,8) ,
71788	 => std_logic_vector(to_unsigned(76,8) ,
71789	 => std_logic_vector(to_unsigned(105,8) ,
71790	 => std_logic_vector(to_unsigned(88,8) ,
71791	 => std_logic_vector(to_unsigned(65,8) ,
71792	 => std_logic_vector(to_unsigned(70,8) ,
71793	 => std_logic_vector(to_unsigned(66,8) ,
71794	 => std_logic_vector(to_unsigned(63,8) ,
71795	 => std_logic_vector(to_unsigned(47,8) ,
71796	 => std_logic_vector(to_unsigned(84,8) ,
71797	 => std_logic_vector(to_unsigned(133,8) ,
71798	 => std_logic_vector(to_unsigned(122,8) ,
71799	 => std_logic_vector(to_unsigned(125,8) ,
71800	 => std_logic_vector(to_unsigned(127,8) ,
71801	 => std_logic_vector(to_unsigned(125,8) ,
71802	 => std_logic_vector(to_unsigned(121,8) ,
71803	 => std_logic_vector(to_unsigned(119,8) ,
71804	 => std_logic_vector(to_unsigned(122,8) ,
71805	 => std_logic_vector(to_unsigned(115,8) ,
71806	 => std_logic_vector(to_unsigned(109,8) ,
71807	 => std_logic_vector(to_unsigned(100,8) ,
71808	 => std_logic_vector(to_unsigned(92,8) ,
71809	 => std_logic_vector(to_unsigned(108,8) ,
71810	 => std_logic_vector(to_unsigned(81,8) ,
71811	 => std_logic_vector(to_unsigned(22,8) ,
71812	 => std_logic_vector(to_unsigned(15,8) ,
71813	 => std_logic_vector(to_unsigned(46,8) ,
71814	 => std_logic_vector(to_unsigned(53,8) ,
71815	 => std_logic_vector(to_unsigned(52,8) ,
71816	 => std_logic_vector(to_unsigned(100,8) ,
71817	 => std_logic_vector(to_unsigned(68,8) ,
71818	 => std_logic_vector(to_unsigned(61,8) ,
71819	 => std_logic_vector(to_unsigned(73,8) ,
71820	 => std_logic_vector(to_unsigned(67,8) ,
71821	 => std_logic_vector(to_unsigned(63,8) ,
71822	 => std_logic_vector(to_unsigned(72,8) ,
71823	 => std_logic_vector(to_unsigned(82,8) ,
71824	 => std_logic_vector(to_unsigned(71,8) ,
71825	 => std_logic_vector(to_unsigned(70,8) ,
71826	 => std_logic_vector(to_unsigned(74,8) ,
71827	 => std_logic_vector(to_unsigned(73,8) ,
71828	 => std_logic_vector(to_unsigned(70,8) ,
71829	 => std_logic_vector(to_unsigned(62,8) ,
71830	 => std_logic_vector(to_unsigned(55,8) ,
71831	 => std_logic_vector(to_unsigned(51,8) ,
71832	 => std_logic_vector(to_unsigned(47,8) ,
71833	 => std_logic_vector(to_unsigned(42,8) ,
71834	 => std_logic_vector(to_unsigned(50,8) ,
71835	 => std_logic_vector(to_unsigned(41,8) ,
71836	 => std_logic_vector(to_unsigned(38,8) ,
71837	 => std_logic_vector(to_unsigned(23,8) ,
71838	 => std_logic_vector(to_unsigned(51,8) ,
71839	 => std_logic_vector(to_unsigned(74,8) ,
71840	 => std_logic_vector(to_unsigned(13,8) ,
71841	 => std_logic_vector(to_unsigned(9,8) ,
71842	 => std_logic_vector(to_unsigned(17,8) ,
71843	 => std_logic_vector(to_unsigned(65,8) ,
71844	 => std_logic_vector(to_unsigned(58,8) ,
71845	 => std_logic_vector(to_unsigned(48,8) ,
71846	 => std_logic_vector(to_unsigned(30,8) ,
71847	 => std_logic_vector(to_unsigned(5,8) ,
71848	 => std_logic_vector(to_unsigned(6,8) ,
71849	 => std_logic_vector(to_unsigned(13,8) ,
71850	 => std_logic_vector(to_unsigned(11,8) ,
71851	 => std_logic_vector(to_unsigned(15,8) ,
71852	 => std_logic_vector(to_unsigned(13,8) ,
71853	 => std_logic_vector(to_unsigned(29,8) ,
71854	 => std_logic_vector(to_unsigned(33,8) ,
71855	 => std_logic_vector(to_unsigned(11,8) ,
71856	 => std_logic_vector(to_unsigned(20,8) ,
71857	 => std_logic_vector(to_unsigned(14,8) ,
71858	 => std_logic_vector(to_unsigned(17,8) ,
71859	 => std_logic_vector(to_unsigned(37,8) ,
71860	 => std_logic_vector(to_unsigned(39,8) ,
71861	 => std_logic_vector(to_unsigned(27,8) ,
71862	 => std_logic_vector(to_unsigned(22,8) ,
71863	 => std_logic_vector(to_unsigned(39,8) ,
71864	 => std_logic_vector(to_unsigned(46,8) ,
71865	 => std_logic_vector(to_unsigned(30,8) ,
71866	 => std_logic_vector(to_unsigned(30,8) ,
71867	 => std_logic_vector(to_unsigned(37,8) ,
71868	 => std_logic_vector(to_unsigned(44,8) ,
71869	 => std_logic_vector(to_unsigned(47,8) ,
71870	 => std_logic_vector(to_unsigned(24,8) ,
71871	 => std_logic_vector(to_unsigned(20,8) ,
71872	 => std_logic_vector(to_unsigned(46,8) ,
71873	 => std_logic_vector(to_unsigned(88,8) ,
71874	 => std_logic_vector(to_unsigned(60,8) ,
71875	 => std_logic_vector(to_unsigned(31,8) ,
71876	 => std_logic_vector(to_unsigned(25,8) ,
71877	 => std_logic_vector(to_unsigned(30,8) ,
71878	 => std_logic_vector(to_unsigned(41,8) ,
71879	 => std_logic_vector(to_unsigned(34,8) ,
71880	 => std_logic_vector(to_unsigned(32,8) ,
71881	 => std_logic_vector(to_unsigned(17,8) ,
71882	 => std_logic_vector(to_unsigned(10,8) ,
71883	 => std_logic_vector(to_unsigned(9,8) ,
71884	 => std_logic_vector(to_unsigned(10,8) ,
71885	 => std_logic_vector(to_unsigned(14,8) ,
71886	 => std_logic_vector(to_unsigned(9,8) ,
71887	 => std_logic_vector(to_unsigned(9,8) ,
71888	 => std_logic_vector(to_unsigned(16,8) ,
71889	 => std_logic_vector(to_unsigned(50,8) ,
71890	 => std_logic_vector(to_unsigned(96,8) ,
71891	 => std_logic_vector(to_unsigned(60,8) ,
71892	 => std_logic_vector(to_unsigned(19,8) ,
71893	 => std_logic_vector(to_unsigned(20,8) ,
71894	 => std_logic_vector(to_unsigned(20,8) ,
71895	 => std_logic_vector(to_unsigned(12,8) ,
71896	 => std_logic_vector(to_unsigned(16,8) ,
71897	 => std_logic_vector(to_unsigned(24,8) ,
71898	 => std_logic_vector(to_unsigned(21,8) ,
71899	 => std_logic_vector(to_unsigned(17,8) ,
71900	 => std_logic_vector(to_unsigned(19,8) ,
71901	 => std_logic_vector(to_unsigned(24,8) ,
71902	 => std_logic_vector(to_unsigned(15,8) ,
71903	 => std_logic_vector(to_unsigned(22,8) ,
71904	 => std_logic_vector(to_unsigned(29,8) ,
71905	 => std_logic_vector(to_unsigned(23,8) ,
71906	 => std_logic_vector(to_unsigned(27,8) ,
71907	 => std_logic_vector(to_unsigned(28,8) ,
71908	 => std_logic_vector(to_unsigned(13,8) ,
71909	 => std_logic_vector(to_unsigned(3,8) ,
71910	 => std_logic_vector(to_unsigned(13,8) ,
71911	 => std_logic_vector(to_unsigned(23,8) ,
71912	 => std_logic_vector(to_unsigned(18,8) ,
71913	 => std_logic_vector(to_unsigned(26,8) ,
71914	 => std_logic_vector(to_unsigned(35,8) ,
71915	 => std_logic_vector(to_unsigned(40,8) ,
71916	 => std_logic_vector(to_unsigned(8,8) ,
71917	 => std_logic_vector(to_unsigned(5,8) ,
71918	 => std_logic_vector(to_unsigned(45,8) ,
71919	 => std_logic_vector(to_unsigned(56,8) ,
71920	 => std_logic_vector(to_unsigned(15,8) ,
71921	 => std_logic_vector(to_unsigned(3,8) ,
71922	 => std_logic_vector(to_unsigned(24,8) ,
71923	 => std_logic_vector(to_unsigned(69,8) ,
71924	 => std_logic_vector(to_unsigned(100,8) ,
71925	 => std_logic_vector(to_unsigned(100,8) ,
71926	 => std_logic_vector(to_unsigned(41,8) ,
71927	 => std_logic_vector(to_unsigned(71,8) ,
71928	 => std_logic_vector(to_unsigned(130,8) ,
71929	 => std_logic_vector(to_unsigned(85,8) ,
71930	 => std_logic_vector(to_unsigned(15,8) ,
71931	 => std_logic_vector(to_unsigned(7,8) ,
71932	 => std_logic_vector(to_unsigned(8,8) ,
71933	 => std_logic_vector(to_unsigned(7,8) ,
71934	 => std_logic_vector(to_unsigned(8,8) ,
71935	 => std_logic_vector(to_unsigned(5,8) ,
71936	 => std_logic_vector(to_unsigned(8,8) ,
71937	 => std_logic_vector(to_unsigned(10,8) ,
71938	 => std_logic_vector(to_unsigned(8,8) ,
71939	 => std_logic_vector(to_unsigned(9,8) ,
71940	 => std_logic_vector(to_unsigned(11,8) ,
71941	 => std_logic_vector(to_unsigned(10,8) ,
71942	 => std_logic_vector(to_unsigned(9,8) ,
71943	 => std_logic_vector(to_unsigned(10,8) ,
71944	 => std_logic_vector(to_unsigned(14,8) ,
71945	 => std_logic_vector(to_unsigned(17,8) ,
71946	 => std_logic_vector(to_unsigned(16,8) ,
71947	 => std_logic_vector(to_unsigned(10,8) ,
71948	 => std_logic_vector(to_unsigned(13,8) ,
71949	 => std_logic_vector(to_unsigned(30,8) ,
71950	 => std_logic_vector(to_unsigned(22,8) ,
71951	 => std_logic_vector(to_unsigned(15,8) ,
71952	 => std_logic_vector(to_unsigned(24,8) ,
71953	 => std_logic_vector(to_unsigned(8,8) ,
71954	 => std_logic_vector(to_unsigned(4,8) ,
71955	 => std_logic_vector(to_unsigned(10,8) ,
71956	 => std_logic_vector(to_unsigned(6,8) ,
71957	 => std_logic_vector(to_unsigned(0,8) ,
71958	 => std_logic_vector(to_unsigned(0,8) ,
71959	 => std_logic_vector(to_unsigned(12,8) ,
71960	 => std_logic_vector(to_unsigned(23,8) ,
71961	 => std_logic_vector(to_unsigned(15,8) ,
71962	 => std_logic_vector(to_unsigned(13,8) ,
71963	 => std_logic_vector(to_unsigned(4,8) ,
71964	 => std_logic_vector(to_unsigned(10,8) ,
71965	 => std_logic_vector(to_unsigned(11,8) ,
71966	 => std_logic_vector(to_unsigned(12,8) ,
71967	 => std_logic_vector(to_unsigned(13,8) ,
71968	 => std_logic_vector(to_unsigned(2,8) ,
71969	 => std_logic_vector(to_unsigned(0,8) ,
71970	 => std_logic_vector(to_unsigned(0,8) ,
71971	 => std_logic_vector(to_unsigned(0,8) ,
71972	 => std_logic_vector(to_unsigned(1,8) ,
71973	 => std_logic_vector(to_unsigned(2,8) ,
71974	 => std_logic_vector(to_unsigned(3,8) ,
71975	 => std_logic_vector(to_unsigned(6,8) ,
71976	 => std_logic_vector(to_unsigned(5,8) ,
71977	 => std_logic_vector(to_unsigned(3,8) ,
71978	 => std_logic_vector(to_unsigned(0,8) ,
71979	 => std_logic_vector(to_unsigned(0,8) ,
71980	 => std_logic_vector(to_unsigned(0,8) ,
71981	 => std_logic_vector(to_unsigned(0,8) ,
71982	 => std_logic_vector(to_unsigned(1,8) ,
71983	 => std_logic_vector(to_unsigned(1,8) ,
71984	 => std_logic_vector(to_unsigned(0,8) ,
71985	 => std_logic_vector(to_unsigned(3,8) ,
71986	 => std_logic_vector(to_unsigned(40,8) ,
71987	 => std_logic_vector(to_unsigned(45,8) ,
71988	 => std_logic_vector(to_unsigned(41,8) ,
71989	 => std_logic_vector(to_unsigned(32,8) ,
71990	 => std_logic_vector(to_unsigned(95,8) ,
71991	 => std_logic_vector(to_unsigned(125,8) ,
71992	 => std_logic_vector(to_unsigned(69,8) ,
71993	 => std_logic_vector(to_unsigned(37,8) ,
71994	 => std_logic_vector(to_unsigned(39,8) ,
71995	 => std_logic_vector(to_unsigned(24,8) ,
71996	 => std_logic_vector(to_unsigned(37,8) ,
71997	 => std_logic_vector(to_unsigned(76,8) ,
71998	 => std_logic_vector(to_unsigned(64,8) ,
71999	 => std_logic_vector(to_unsigned(56,8) ,
72000	 => std_logic_vector(to_unsigned(39,8) ,
72001	 => std_logic_vector(to_unsigned(122,8) ,
72002	 => std_logic_vector(to_unsigned(127,8) ,
72003	 => std_logic_vector(to_unsigned(142,8) ,
72004	 => std_logic_vector(to_unsigned(138,8) ,
72005	 => std_logic_vector(to_unsigned(144,8) ,
72006	 => std_logic_vector(to_unsigned(128,8) ,
72007	 => std_logic_vector(to_unsigned(104,8) ,
72008	 => std_logic_vector(to_unsigned(104,8) ,
72009	 => std_logic_vector(to_unsigned(104,8) ,
72010	 => std_logic_vector(to_unsigned(93,8) ,
72011	 => std_logic_vector(to_unsigned(77,8) ,
72012	 => std_logic_vector(to_unsigned(68,8) ,
72013	 => std_logic_vector(to_unsigned(77,8) ,
72014	 => std_logic_vector(to_unsigned(80,8) ,
72015	 => std_logic_vector(to_unsigned(85,8) ,
72016	 => std_logic_vector(to_unsigned(78,8) ,
72017	 => std_logic_vector(to_unsigned(76,8) ,
72018	 => std_logic_vector(to_unsigned(85,8) ,
72019	 => std_logic_vector(to_unsigned(76,8) ,
72020	 => std_logic_vector(to_unsigned(63,8) ,
72021	 => std_logic_vector(to_unsigned(57,8) ,
72022	 => std_logic_vector(to_unsigned(54,8) ,
72023	 => std_logic_vector(to_unsigned(52,8) ,
72024	 => std_logic_vector(to_unsigned(50,8) ,
72025	 => std_logic_vector(to_unsigned(46,8) ,
72026	 => std_logic_vector(to_unsigned(44,8) ,
72027	 => std_logic_vector(to_unsigned(41,8) ,
72028	 => std_logic_vector(to_unsigned(37,8) ,
72029	 => std_logic_vector(to_unsigned(45,8) ,
72030	 => std_logic_vector(to_unsigned(47,8) ,
72031	 => std_logic_vector(to_unsigned(32,8) ,
72032	 => std_logic_vector(to_unsigned(27,8) ,
72033	 => std_logic_vector(to_unsigned(45,8) ,
72034	 => std_logic_vector(to_unsigned(38,8) ,
72035	 => std_logic_vector(to_unsigned(46,8) ,
72036	 => std_logic_vector(to_unsigned(62,8) ,
72037	 => std_logic_vector(to_unsigned(92,8) ,
72038	 => std_logic_vector(to_unsigned(92,8) ,
72039	 => std_logic_vector(to_unsigned(32,8) ,
72040	 => std_logic_vector(to_unsigned(20,8) ,
72041	 => std_logic_vector(to_unsigned(26,8) ,
72042	 => std_logic_vector(to_unsigned(22,8) ,
72043	 => std_logic_vector(to_unsigned(19,8) ,
72044	 => std_logic_vector(to_unsigned(28,8) ,
72045	 => std_logic_vector(to_unsigned(30,8) ,
72046	 => std_logic_vector(to_unsigned(28,8) ,
72047	 => std_logic_vector(to_unsigned(26,8) ,
72048	 => std_logic_vector(to_unsigned(30,8) ,
72049	 => std_logic_vector(to_unsigned(23,8) ,
72050	 => std_logic_vector(to_unsigned(25,8) ,
72051	 => std_logic_vector(to_unsigned(39,8) ,
72052	 => std_logic_vector(to_unsigned(37,8) ,
72053	 => std_logic_vector(to_unsigned(40,8) ,
72054	 => std_logic_vector(to_unsigned(37,8) ,
72055	 => std_logic_vector(to_unsigned(37,8) ,
72056	 => std_logic_vector(to_unsigned(43,8) ,
72057	 => std_logic_vector(to_unsigned(50,8) ,
72058	 => std_logic_vector(to_unsigned(50,8) ,
72059	 => std_logic_vector(to_unsigned(46,8) ,
72060	 => std_logic_vector(to_unsigned(50,8) ,
72061	 => std_logic_vector(to_unsigned(53,8) ,
72062	 => std_logic_vector(to_unsigned(51,8) ,
72063	 => std_logic_vector(to_unsigned(49,8) ,
72064	 => std_logic_vector(to_unsigned(40,8) ,
72065	 => std_logic_vector(to_unsigned(43,8) ,
72066	 => std_logic_vector(to_unsigned(44,8) ,
72067	 => std_logic_vector(to_unsigned(36,8) ,
72068	 => std_logic_vector(to_unsigned(44,8) ,
72069	 => std_logic_vector(to_unsigned(37,8) ,
72070	 => std_logic_vector(to_unsigned(40,8) ,
72071	 => std_logic_vector(to_unsigned(45,8) ,
72072	 => std_logic_vector(to_unsigned(39,8) ,
72073	 => std_logic_vector(to_unsigned(49,8) ,
72074	 => std_logic_vector(to_unsigned(64,8) ,
72075	 => std_logic_vector(to_unsigned(59,8) ,
72076	 => std_logic_vector(to_unsigned(71,8) ,
72077	 => std_logic_vector(to_unsigned(64,8) ,
72078	 => std_logic_vector(to_unsigned(62,8) ,
72079	 => std_logic_vector(to_unsigned(80,8) ,
72080	 => std_logic_vector(to_unsigned(77,8) ,
72081	 => std_logic_vector(to_unsigned(71,8) ,
72082	 => std_logic_vector(to_unsigned(67,8) ,
72083	 => std_logic_vector(to_unsigned(81,8) ,
72084	 => std_logic_vector(to_unsigned(67,8) ,
72085	 => std_logic_vector(to_unsigned(64,8) ,
72086	 => std_logic_vector(to_unsigned(82,8) ,
72087	 => std_logic_vector(to_unsigned(90,8) ,
72088	 => std_logic_vector(to_unsigned(87,8) ,
72089	 => std_logic_vector(to_unsigned(86,8) ,
72090	 => std_logic_vector(to_unsigned(69,8) ,
72091	 => std_logic_vector(to_unsigned(49,8) ,
72092	 => std_logic_vector(to_unsigned(48,8) ,
72093	 => std_logic_vector(to_unsigned(51,8) ,
72094	 => std_logic_vector(to_unsigned(42,8) ,
72095	 => std_logic_vector(to_unsigned(45,8) ,
72096	 => std_logic_vector(to_unsigned(51,8) ,
72097	 => std_logic_vector(to_unsigned(50,8) ,
72098	 => std_logic_vector(to_unsigned(41,8) ,
72099	 => std_logic_vector(to_unsigned(37,8) ,
72100	 => std_logic_vector(to_unsigned(27,8) ,
72101	 => std_logic_vector(to_unsigned(24,8) ,
72102	 => std_logic_vector(to_unsigned(27,8) ,
72103	 => std_logic_vector(to_unsigned(45,8) ,
72104	 => std_logic_vector(to_unsigned(57,8) ,
72105	 => std_logic_vector(to_unsigned(64,8) ,
72106	 => std_logic_vector(to_unsigned(82,8) ,
72107	 => std_logic_vector(to_unsigned(99,8) ,
72108	 => std_logic_vector(to_unsigned(147,8) ,
72109	 => std_logic_vector(to_unsigned(170,8) ,
72110	 => std_logic_vector(to_unsigned(146,8) ,
72111	 => std_logic_vector(to_unsigned(86,8) ,
72112	 => std_logic_vector(to_unsigned(64,8) ,
72113	 => std_logic_vector(to_unsigned(68,8) ,
72114	 => std_logic_vector(to_unsigned(66,8) ,
72115	 => std_logic_vector(to_unsigned(49,8) ,
72116	 => std_logic_vector(to_unsigned(69,8) ,
72117	 => std_logic_vector(to_unsigned(115,8) ,
72118	 => std_logic_vector(to_unsigned(111,8) ,
72119	 => std_logic_vector(to_unsigned(114,8) ,
72120	 => std_logic_vector(to_unsigned(118,8) ,
72121	 => std_logic_vector(to_unsigned(122,8) ,
72122	 => std_logic_vector(to_unsigned(119,8) ,
72123	 => std_logic_vector(to_unsigned(119,8) ,
72124	 => std_logic_vector(to_unsigned(118,8) ,
72125	 => std_logic_vector(to_unsigned(108,8) ,
72126	 => std_logic_vector(to_unsigned(100,8) ,
72127	 => std_logic_vector(to_unsigned(90,8) ,
72128	 => std_logic_vector(to_unsigned(78,8) ,
72129	 => std_logic_vector(to_unsigned(88,8) ,
72130	 => std_logic_vector(to_unsigned(74,8) ,
72131	 => std_logic_vector(to_unsigned(56,8) ,
72132	 => std_logic_vector(to_unsigned(57,8) ,
72133	 => std_logic_vector(to_unsigned(77,8) ,
72134	 => std_logic_vector(to_unsigned(90,8) ,
72135	 => std_logic_vector(to_unsigned(121,8) ,
72136	 => std_logic_vector(to_unsigned(112,8) ,
72137	 => std_logic_vector(to_unsigned(42,8) ,
72138	 => std_logic_vector(to_unsigned(36,8) ,
72139	 => std_logic_vector(to_unsigned(58,8) ,
72140	 => std_logic_vector(to_unsigned(64,8) ,
72141	 => std_logic_vector(to_unsigned(69,8) ,
72142	 => std_logic_vector(to_unsigned(63,8) ,
72143	 => std_logic_vector(to_unsigned(73,8) ,
72144	 => std_logic_vector(to_unsigned(60,8) ,
72145	 => std_logic_vector(to_unsigned(58,8) ,
72146	 => std_logic_vector(to_unsigned(65,8) ,
72147	 => std_logic_vector(to_unsigned(62,8) ,
72148	 => std_logic_vector(to_unsigned(59,8) ,
72149	 => std_logic_vector(to_unsigned(64,8) ,
72150	 => std_logic_vector(to_unsigned(61,8) ,
72151	 => std_logic_vector(to_unsigned(60,8) ,
72152	 => std_logic_vector(to_unsigned(51,8) ,
72153	 => std_logic_vector(to_unsigned(35,8) ,
72154	 => std_logic_vector(to_unsigned(27,8) ,
72155	 => std_logic_vector(to_unsigned(27,8) ,
72156	 => std_logic_vector(to_unsigned(73,8) ,
72157	 => std_logic_vector(to_unsigned(54,8) ,
72158	 => std_logic_vector(to_unsigned(40,8) ,
72159	 => std_logic_vector(to_unsigned(69,8) ,
72160	 => std_logic_vector(to_unsigned(38,8) ,
72161	 => std_logic_vector(to_unsigned(37,8) ,
72162	 => std_logic_vector(to_unsigned(63,8) ,
72163	 => std_logic_vector(to_unsigned(53,8) ,
72164	 => std_logic_vector(to_unsigned(35,8) ,
72165	 => std_logic_vector(to_unsigned(46,8) ,
72166	 => std_logic_vector(to_unsigned(32,8) ,
72167	 => std_logic_vector(to_unsigned(6,8) ,
72168	 => std_logic_vector(to_unsigned(6,8) ,
72169	 => std_logic_vector(to_unsigned(13,8) ,
72170	 => std_logic_vector(to_unsigned(13,8) ,
72171	 => std_logic_vector(to_unsigned(12,8) ,
72172	 => std_logic_vector(to_unsigned(23,8) ,
72173	 => std_logic_vector(to_unsigned(37,8) ,
72174	 => std_logic_vector(to_unsigned(18,8) ,
72175	 => std_logic_vector(to_unsigned(17,8) ,
72176	 => std_logic_vector(to_unsigned(15,8) ,
72177	 => std_logic_vector(to_unsigned(18,8) ,
72178	 => std_logic_vector(to_unsigned(33,8) ,
72179	 => std_logic_vector(to_unsigned(36,8) ,
72180	 => std_logic_vector(to_unsigned(49,8) ,
72181	 => std_logic_vector(to_unsigned(20,8) ,
72182	 => std_logic_vector(to_unsigned(5,8) ,
72183	 => std_logic_vector(to_unsigned(10,8) ,
72184	 => std_logic_vector(to_unsigned(12,8) ,
72185	 => std_logic_vector(to_unsigned(11,8) ,
72186	 => std_logic_vector(to_unsigned(23,8) ,
72187	 => std_logic_vector(to_unsigned(39,8) ,
72188	 => std_logic_vector(to_unsigned(57,8) ,
72189	 => std_logic_vector(to_unsigned(41,8) ,
72190	 => std_logic_vector(to_unsigned(25,8) ,
72191	 => std_logic_vector(to_unsigned(23,8) ,
72192	 => std_logic_vector(to_unsigned(32,8) ,
72193	 => std_logic_vector(to_unsigned(50,8) ,
72194	 => std_logic_vector(to_unsigned(46,8) ,
72195	 => std_logic_vector(to_unsigned(23,8) ,
72196	 => std_logic_vector(to_unsigned(22,8) ,
72197	 => std_logic_vector(to_unsigned(40,8) ,
72198	 => std_logic_vector(to_unsigned(53,8) ,
72199	 => std_logic_vector(to_unsigned(51,8) ,
72200	 => std_logic_vector(to_unsigned(32,8) ,
72201	 => std_logic_vector(to_unsigned(25,8) ,
72202	 => std_logic_vector(to_unsigned(12,8) ,
72203	 => std_logic_vector(to_unsigned(6,8) ,
72204	 => std_logic_vector(to_unsigned(11,8) ,
72205	 => std_logic_vector(to_unsigned(12,8) ,
72206	 => std_logic_vector(to_unsigned(7,8) ,
72207	 => std_logic_vector(to_unsigned(9,8) ,
72208	 => std_logic_vector(to_unsigned(21,8) ,
72209	 => std_logic_vector(to_unsigned(40,8) ,
72210	 => std_logic_vector(to_unsigned(64,8) ,
72211	 => std_logic_vector(to_unsigned(47,8) ,
72212	 => std_logic_vector(to_unsigned(18,8) ,
72213	 => std_logic_vector(to_unsigned(20,8) ,
72214	 => std_logic_vector(to_unsigned(27,8) ,
72215	 => std_logic_vector(to_unsigned(17,8) ,
72216	 => std_logic_vector(to_unsigned(10,8) ,
72217	 => std_logic_vector(to_unsigned(19,8) ,
72218	 => std_logic_vector(to_unsigned(24,8) ,
72219	 => std_logic_vector(to_unsigned(21,8) ,
72220	 => std_logic_vector(to_unsigned(13,8) ,
72221	 => std_logic_vector(to_unsigned(13,8) ,
72222	 => std_logic_vector(to_unsigned(16,8) ,
72223	 => std_logic_vector(to_unsigned(24,8) ,
72224	 => std_logic_vector(to_unsigned(32,8) ,
72225	 => std_logic_vector(to_unsigned(22,8) ,
72226	 => std_logic_vector(to_unsigned(27,8) ,
72227	 => std_logic_vector(to_unsigned(34,8) ,
72228	 => std_logic_vector(to_unsigned(17,8) ,
72229	 => std_logic_vector(to_unsigned(4,8) ,
72230	 => std_logic_vector(to_unsigned(14,8) ,
72231	 => std_logic_vector(to_unsigned(35,8) ,
72232	 => std_logic_vector(to_unsigned(31,8) ,
72233	 => std_logic_vector(to_unsigned(25,8) ,
72234	 => std_logic_vector(to_unsigned(34,8) ,
72235	 => std_logic_vector(to_unsigned(42,8) ,
72236	 => std_logic_vector(to_unsigned(27,8) ,
72237	 => std_logic_vector(to_unsigned(19,8) ,
72238	 => std_logic_vector(to_unsigned(45,8) ,
72239	 => std_logic_vector(to_unsigned(54,8) ,
72240	 => std_logic_vector(to_unsigned(29,8) ,
72241	 => std_logic_vector(to_unsigned(20,8) ,
72242	 => std_logic_vector(to_unsigned(30,8) ,
72243	 => std_logic_vector(to_unsigned(67,8) ,
72244	 => std_logic_vector(to_unsigned(93,8) ,
72245	 => std_logic_vector(to_unsigned(87,8) ,
72246	 => std_logic_vector(to_unsigned(38,8) ,
72247	 => std_logic_vector(to_unsigned(74,8) ,
72248	 => std_logic_vector(to_unsigned(134,8) ,
72249	 => std_logic_vector(to_unsigned(95,8) ,
72250	 => std_logic_vector(to_unsigned(19,8) ,
72251	 => std_logic_vector(to_unsigned(8,8) ,
72252	 => std_logic_vector(to_unsigned(11,8) ,
72253	 => std_logic_vector(to_unsigned(9,8) ,
72254	 => std_logic_vector(to_unsigned(9,8) ,
72255	 => std_logic_vector(to_unsigned(7,8) ,
72256	 => std_logic_vector(to_unsigned(8,8) ,
72257	 => std_logic_vector(to_unsigned(10,8) ,
72258	 => std_logic_vector(to_unsigned(9,8) ,
72259	 => std_logic_vector(to_unsigned(8,8) ,
72260	 => std_logic_vector(to_unsigned(6,8) ,
72261	 => std_logic_vector(to_unsigned(8,8) ,
72262	 => std_logic_vector(to_unsigned(8,8) ,
72263	 => std_logic_vector(to_unsigned(8,8) ,
72264	 => std_logic_vector(to_unsigned(10,8) ,
72265	 => std_logic_vector(to_unsigned(13,8) ,
72266	 => std_logic_vector(to_unsigned(13,8) ,
72267	 => std_logic_vector(to_unsigned(13,8) ,
72268	 => std_logic_vector(to_unsigned(15,8) ,
72269	 => std_logic_vector(to_unsigned(25,8) ,
72270	 => std_logic_vector(to_unsigned(17,8) ,
72271	 => std_logic_vector(to_unsigned(7,8) ,
72272	 => std_logic_vector(to_unsigned(19,8) ,
72273	 => std_logic_vector(to_unsigned(24,8) ,
72274	 => std_logic_vector(to_unsigned(15,8) ,
72275	 => std_logic_vector(to_unsigned(35,8) ,
72276	 => std_logic_vector(to_unsigned(17,8) ,
72277	 => std_logic_vector(to_unsigned(2,8) ,
72278	 => std_logic_vector(to_unsigned(0,8) ,
72279	 => std_logic_vector(to_unsigned(7,8) ,
72280	 => std_logic_vector(to_unsigned(39,8) ,
72281	 => std_logic_vector(to_unsigned(37,8) ,
72282	 => std_logic_vector(to_unsigned(24,8) ,
72283	 => std_logic_vector(to_unsigned(8,8) ,
72284	 => std_logic_vector(to_unsigned(23,8) ,
72285	 => std_logic_vector(to_unsigned(20,8) ,
72286	 => std_logic_vector(to_unsigned(18,8) ,
72287	 => std_logic_vector(to_unsigned(19,8) ,
72288	 => std_logic_vector(to_unsigned(4,8) ,
72289	 => std_logic_vector(to_unsigned(0,8) ,
72290	 => std_logic_vector(to_unsigned(0,8) ,
72291	 => std_logic_vector(to_unsigned(0,8) ,
72292	 => std_logic_vector(to_unsigned(1,8) ,
72293	 => std_logic_vector(to_unsigned(1,8) ,
72294	 => std_logic_vector(to_unsigned(1,8) ,
72295	 => std_logic_vector(to_unsigned(1,8) ,
72296	 => std_logic_vector(to_unsigned(1,8) ,
72297	 => std_logic_vector(to_unsigned(5,8) ,
72298	 => std_logic_vector(to_unsigned(5,8) ,
72299	 => std_logic_vector(to_unsigned(1,8) ,
72300	 => std_logic_vector(to_unsigned(0,8) ,
72301	 => std_logic_vector(to_unsigned(0,8) ,
72302	 => std_logic_vector(to_unsigned(1,8) ,
72303	 => std_logic_vector(to_unsigned(2,8) ,
72304	 => std_logic_vector(to_unsigned(1,8) ,
72305	 => std_logic_vector(to_unsigned(3,8) ,
72306	 => std_logic_vector(to_unsigned(31,8) ,
72307	 => std_logic_vector(to_unsigned(37,8) ,
72308	 => std_logic_vector(to_unsigned(25,8) ,
72309	 => std_logic_vector(to_unsigned(17,8) ,
72310	 => std_logic_vector(to_unsigned(92,8) ,
72311	 => std_logic_vector(to_unsigned(146,8) ,
72312	 => std_logic_vector(to_unsigned(70,8) ,
72313	 => std_logic_vector(to_unsigned(50,8) ,
72314	 => std_logic_vector(to_unsigned(57,8) ,
72315	 => std_logic_vector(to_unsigned(30,8) ,
72316	 => std_logic_vector(to_unsigned(51,8) ,
72317	 => std_logic_vector(to_unsigned(77,8) ,
72318	 => std_logic_vector(to_unsigned(72,8) ,
72319	 => std_logic_vector(to_unsigned(79,8) ,
72320	 => std_logic_vector(to_unsigned(85,8) ,
72321	 => std_logic_vector(to_unsigned(136,8) ,
72322	 => std_logic_vector(to_unsigned(133,8) ,
72323	 => std_logic_vector(to_unsigned(142,8) ,
72324	 => std_logic_vector(to_unsigned(134,8) ,
72325	 => std_logic_vector(to_unsigned(119,8) ,
72326	 => std_logic_vector(to_unsigned(103,8) ,
72327	 => std_logic_vector(to_unsigned(93,8) ,
72328	 => std_logic_vector(to_unsigned(103,8) ,
72329	 => std_logic_vector(to_unsigned(79,8) ,
72330	 => std_logic_vector(to_unsigned(68,8) ,
72331	 => std_logic_vector(to_unsigned(79,8) ,
72332	 => std_logic_vector(to_unsigned(91,8) ,
72333	 => std_logic_vector(to_unsigned(91,8) ,
72334	 => std_logic_vector(to_unsigned(79,8) ,
72335	 => std_logic_vector(to_unsigned(81,8) ,
72336	 => std_logic_vector(to_unsigned(80,8) ,
72337	 => std_logic_vector(to_unsigned(79,8) ,
72338	 => std_logic_vector(to_unsigned(80,8) ,
72339	 => std_logic_vector(to_unsigned(70,8) ,
72340	 => std_logic_vector(to_unsigned(63,8) ,
72341	 => std_logic_vector(to_unsigned(61,8) ,
72342	 => std_logic_vector(to_unsigned(55,8) ,
72343	 => std_logic_vector(to_unsigned(57,8) ,
72344	 => std_logic_vector(to_unsigned(55,8) ,
72345	 => std_logic_vector(to_unsigned(48,8) ,
72346	 => std_logic_vector(to_unsigned(40,8) ,
72347	 => std_logic_vector(to_unsigned(37,8) ,
72348	 => std_logic_vector(to_unsigned(40,8) ,
72349	 => std_logic_vector(to_unsigned(45,8) ,
72350	 => std_logic_vector(to_unsigned(66,8) ,
72351	 => std_logic_vector(to_unsigned(54,8) ,
72352	 => std_logic_vector(to_unsigned(25,8) ,
72353	 => std_logic_vector(to_unsigned(32,8) ,
72354	 => std_logic_vector(to_unsigned(10,8) ,
72355	 => std_logic_vector(to_unsigned(10,8) ,
72356	 => std_logic_vector(to_unsigned(13,8) ,
72357	 => std_logic_vector(to_unsigned(24,8) ,
72358	 => std_logic_vector(to_unsigned(45,8) ,
72359	 => std_logic_vector(to_unsigned(43,8) ,
72360	 => std_logic_vector(to_unsigned(25,8) ,
72361	 => std_logic_vector(to_unsigned(30,8) ,
72362	 => std_logic_vector(to_unsigned(32,8) ,
72363	 => std_logic_vector(to_unsigned(31,8) ,
72364	 => std_logic_vector(to_unsigned(32,8) ,
72365	 => std_logic_vector(to_unsigned(26,8) ,
72366	 => std_logic_vector(to_unsigned(41,8) ,
72367	 => std_logic_vector(to_unsigned(44,8) ,
72368	 => std_logic_vector(to_unsigned(34,8) ,
72369	 => std_logic_vector(to_unsigned(22,8) ,
72370	 => std_logic_vector(to_unsigned(33,8) ,
72371	 => std_logic_vector(to_unsigned(46,8) ,
72372	 => std_logic_vector(to_unsigned(37,8) ,
72373	 => std_logic_vector(to_unsigned(38,8) ,
72374	 => std_logic_vector(to_unsigned(37,8) ,
72375	 => std_logic_vector(to_unsigned(35,8) ,
72376	 => std_logic_vector(to_unsigned(41,8) ,
72377	 => std_logic_vector(to_unsigned(44,8) ,
72378	 => std_logic_vector(to_unsigned(41,8) ,
72379	 => std_logic_vector(to_unsigned(43,8) ,
72380	 => std_logic_vector(to_unsigned(49,8) ,
72381	 => std_logic_vector(to_unsigned(51,8) ,
72382	 => std_logic_vector(to_unsigned(44,8) ,
72383	 => std_logic_vector(to_unsigned(47,8) ,
72384	 => std_logic_vector(to_unsigned(67,8) ,
72385	 => std_logic_vector(to_unsigned(79,8) ,
72386	 => std_logic_vector(to_unsigned(68,8) ,
72387	 => std_logic_vector(to_unsigned(51,8) ,
72388	 => std_logic_vector(to_unsigned(47,8) ,
72389	 => std_logic_vector(to_unsigned(44,8) ,
72390	 => std_logic_vector(to_unsigned(47,8) ,
72391	 => std_logic_vector(to_unsigned(44,8) ,
72392	 => std_logic_vector(to_unsigned(40,8) ,
72393	 => std_logic_vector(to_unsigned(51,8) ,
72394	 => std_logic_vector(to_unsigned(70,8) ,
72395	 => std_logic_vector(to_unsigned(66,8) ,
72396	 => std_logic_vector(to_unsigned(68,8) ,
72397	 => std_logic_vector(to_unsigned(61,8) ,
72398	 => std_logic_vector(to_unsigned(69,8) ,
72399	 => std_logic_vector(to_unsigned(78,8) ,
72400	 => std_logic_vector(to_unsigned(81,8) ,
72401	 => std_logic_vector(to_unsigned(81,8) ,
72402	 => std_logic_vector(to_unsigned(61,8) ,
72403	 => std_logic_vector(to_unsigned(57,8) ,
72404	 => std_logic_vector(to_unsigned(76,8) ,
72405	 => std_logic_vector(to_unsigned(69,8) ,
72406	 => std_logic_vector(to_unsigned(65,8) ,
72407	 => std_logic_vector(to_unsigned(92,8) ,
72408	 => std_logic_vector(to_unsigned(78,8) ,
72409	 => std_logic_vector(to_unsigned(57,8) ,
72410	 => std_logic_vector(to_unsigned(41,8) ,
72411	 => std_logic_vector(to_unsigned(43,8) ,
72412	 => std_logic_vector(to_unsigned(51,8) ,
72413	 => std_logic_vector(to_unsigned(45,8) ,
72414	 => std_logic_vector(to_unsigned(40,8) ,
72415	 => std_logic_vector(to_unsigned(41,8) ,
72416	 => std_logic_vector(to_unsigned(45,8) ,
72417	 => std_logic_vector(to_unsigned(35,8) ,
72418	 => std_logic_vector(to_unsigned(24,8) ,
72419	 => std_logic_vector(to_unsigned(35,8) ,
72420	 => std_logic_vector(to_unsigned(39,8) ,
72421	 => std_logic_vector(to_unsigned(34,8) ,
72422	 => std_logic_vector(to_unsigned(30,8) ,
72423	 => std_logic_vector(to_unsigned(45,8) ,
72424	 => std_logic_vector(to_unsigned(93,8) ,
72425	 => std_logic_vector(to_unsigned(81,8) ,
72426	 => std_logic_vector(to_unsigned(80,8) ,
72427	 => std_logic_vector(to_unsigned(108,8) ,
72428	 => std_logic_vector(to_unsigned(134,8) ,
72429	 => std_logic_vector(to_unsigned(147,8) ,
72430	 => std_logic_vector(to_unsigned(163,8) ,
72431	 => std_logic_vector(to_unsigned(146,8) ,
72432	 => std_logic_vector(to_unsigned(82,8) ,
72433	 => std_logic_vector(to_unsigned(68,8) ,
72434	 => std_logic_vector(to_unsigned(69,8) ,
72435	 => std_logic_vector(to_unsigned(48,8) ,
72436	 => std_logic_vector(to_unsigned(61,8) ,
72437	 => std_logic_vector(to_unsigned(108,8) ,
72438	 => std_logic_vector(to_unsigned(108,8) ,
72439	 => std_logic_vector(to_unsigned(104,8) ,
72440	 => std_logic_vector(to_unsigned(101,8) ,
72441	 => std_logic_vector(to_unsigned(104,8) ,
72442	 => std_logic_vector(to_unsigned(109,8) ,
72443	 => std_logic_vector(to_unsigned(108,8) ,
72444	 => std_logic_vector(to_unsigned(107,8) ,
72445	 => std_logic_vector(to_unsigned(101,8) ,
72446	 => std_logic_vector(to_unsigned(96,8) ,
72447	 => std_logic_vector(to_unsigned(92,8) ,
72448	 => std_logic_vector(to_unsigned(66,8) ,
72449	 => std_logic_vector(to_unsigned(43,8) ,
72450	 => std_logic_vector(to_unsigned(24,8) ,
72451	 => std_logic_vector(to_unsigned(10,8) ,
72452	 => std_logic_vector(to_unsigned(29,8) ,
72453	 => std_logic_vector(to_unsigned(84,8) ,
72454	 => std_logic_vector(to_unsigned(101,8) ,
72455	 => std_logic_vector(to_unsigned(99,8) ,
72456	 => std_logic_vector(to_unsigned(87,8) ,
72457	 => std_logic_vector(to_unsigned(45,8) ,
72458	 => std_logic_vector(to_unsigned(27,8) ,
72459	 => std_logic_vector(to_unsigned(32,8) ,
72460	 => std_logic_vector(to_unsigned(32,8) ,
72461	 => std_logic_vector(to_unsigned(38,8) ,
72462	 => std_logic_vector(to_unsigned(55,8) ,
72463	 => std_logic_vector(to_unsigned(49,8) ,
72464	 => std_logic_vector(to_unsigned(60,8) ,
72465	 => std_logic_vector(to_unsigned(57,8) ,
72466	 => std_logic_vector(to_unsigned(51,8) ,
72467	 => std_logic_vector(to_unsigned(52,8) ,
72468	 => std_logic_vector(to_unsigned(47,8) ,
72469	 => std_logic_vector(to_unsigned(57,8) ,
72470	 => std_logic_vector(to_unsigned(80,8) ,
72471	 => std_logic_vector(to_unsigned(58,8) ,
72472	 => std_logic_vector(to_unsigned(40,8) ,
72473	 => std_logic_vector(to_unsigned(32,8) ,
72474	 => std_logic_vector(to_unsigned(19,8) ,
72475	 => std_logic_vector(to_unsigned(36,8) ,
72476	 => std_logic_vector(to_unsigned(88,8) ,
72477	 => std_logic_vector(to_unsigned(63,8) ,
72478	 => std_logic_vector(to_unsigned(52,8) ,
72479	 => std_logic_vector(to_unsigned(74,8) ,
72480	 => std_logic_vector(to_unsigned(73,8) ,
72481	 => std_logic_vector(to_unsigned(74,8) ,
72482	 => std_logic_vector(to_unsigned(55,8) ,
72483	 => std_logic_vector(to_unsigned(29,8) ,
72484	 => std_logic_vector(to_unsigned(25,8) ,
72485	 => std_logic_vector(to_unsigned(44,8) ,
72486	 => std_logic_vector(to_unsigned(34,8) ,
72487	 => std_logic_vector(to_unsigned(6,8) ,
72488	 => std_logic_vector(to_unsigned(5,8) ,
72489	 => std_logic_vector(to_unsigned(12,8) ,
72490	 => std_logic_vector(to_unsigned(10,8) ,
72491	 => std_logic_vector(to_unsigned(23,8) ,
72492	 => std_logic_vector(to_unsigned(43,8) ,
72493	 => std_logic_vector(to_unsigned(12,8) ,
72494	 => std_logic_vector(to_unsigned(17,8) ,
72495	 => std_logic_vector(to_unsigned(17,8) ,
72496	 => std_logic_vector(to_unsigned(14,8) ,
72497	 => std_logic_vector(to_unsigned(35,8) ,
72498	 => std_logic_vector(to_unsigned(32,8) ,
72499	 => std_logic_vector(to_unsigned(40,8) ,
72500	 => std_logic_vector(to_unsigned(60,8) ,
72501	 => std_logic_vector(to_unsigned(24,8) ,
72502	 => std_logic_vector(to_unsigned(9,8) ,
72503	 => std_logic_vector(to_unsigned(11,8) ,
72504	 => std_logic_vector(to_unsigned(10,8) ,
72505	 => std_logic_vector(to_unsigned(12,8) ,
72506	 => std_logic_vector(to_unsigned(19,8) ,
72507	 => std_logic_vector(to_unsigned(45,8) ,
72508	 => std_logic_vector(to_unsigned(78,8) ,
72509	 => std_logic_vector(to_unsigned(59,8) ,
72510	 => std_logic_vector(to_unsigned(27,8) ,
72511	 => std_logic_vector(to_unsigned(23,8) ,
72512	 => std_logic_vector(to_unsigned(35,8) ,
72513	 => std_logic_vector(to_unsigned(39,8) ,
72514	 => std_logic_vector(to_unsigned(29,8) ,
72515	 => std_logic_vector(to_unsigned(21,8) ,
72516	 => std_logic_vector(to_unsigned(23,8) ,
72517	 => std_logic_vector(to_unsigned(35,8) ,
72518	 => std_logic_vector(to_unsigned(45,8) ,
72519	 => std_logic_vector(to_unsigned(41,8) ,
72520	 => std_logic_vector(to_unsigned(27,8) ,
72521	 => std_logic_vector(to_unsigned(22,8) ,
72522	 => std_logic_vector(to_unsigned(9,8) ,
72523	 => std_logic_vector(to_unsigned(8,8) ,
72524	 => std_logic_vector(to_unsigned(17,8) ,
72525	 => std_logic_vector(to_unsigned(18,8) ,
72526	 => std_logic_vector(to_unsigned(10,8) ,
72527	 => std_logic_vector(to_unsigned(9,8) ,
72528	 => std_logic_vector(to_unsigned(18,8) ,
72529	 => std_logic_vector(to_unsigned(15,8) ,
72530	 => std_logic_vector(to_unsigned(17,8) ,
72531	 => std_logic_vector(to_unsigned(17,8) ,
72532	 => std_logic_vector(to_unsigned(19,8) ,
72533	 => std_logic_vector(to_unsigned(22,8) ,
72534	 => std_logic_vector(to_unsigned(28,8) ,
72535	 => std_logic_vector(to_unsigned(31,8) ,
72536	 => std_logic_vector(to_unsigned(25,8) ,
72537	 => std_logic_vector(to_unsigned(18,8) ,
72538	 => std_logic_vector(to_unsigned(19,8) ,
72539	 => std_logic_vector(to_unsigned(23,8) ,
72540	 => std_logic_vector(to_unsigned(17,8) ,
72541	 => std_logic_vector(to_unsigned(12,8) ,
72542	 => std_logic_vector(to_unsigned(16,8) ,
72543	 => std_logic_vector(to_unsigned(25,8) ,
72544	 => std_logic_vector(to_unsigned(38,8) ,
72545	 => std_logic_vector(to_unsigned(31,8) ,
72546	 => std_logic_vector(to_unsigned(25,8) ,
72547	 => std_logic_vector(to_unsigned(24,8) ,
72548	 => std_logic_vector(to_unsigned(13,8) ,
72549	 => std_logic_vector(to_unsigned(3,8) ,
72550	 => std_logic_vector(to_unsigned(14,8) ,
72551	 => std_logic_vector(to_unsigned(30,8) ,
72552	 => std_logic_vector(to_unsigned(23,8) ,
72553	 => std_logic_vector(to_unsigned(10,8) ,
72554	 => std_logic_vector(to_unsigned(23,8) ,
72555	 => std_logic_vector(to_unsigned(41,8) ,
72556	 => std_logic_vector(to_unsigned(27,8) ,
72557	 => std_logic_vector(to_unsigned(30,8) ,
72558	 => std_logic_vector(to_unsigned(51,8) ,
72559	 => std_logic_vector(to_unsigned(45,8) ,
72560	 => std_logic_vector(to_unsigned(29,8) ,
72561	 => std_logic_vector(to_unsigned(33,8) ,
72562	 => std_logic_vector(to_unsigned(35,8) ,
72563	 => std_logic_vector(to_unsigned(67,8) ,
72564	 => std_logic_vector(to_unsigned(104,8) ,
72565	 => std_logic_vector(to_unsigned(86,8) ,
72566	 => std_logic_vector(to_unsigned(39,8) ,
72567	 => std_logic_vector(to_unsigned(76,8) ,
72568	 => std_logic_vector(to_unsigned(121,8) ,
72569	 => std_logic_vector(to_unsigned(97,8) ,
72570	 => std_logic_vector(to_unsigned(13,8) ,
72571	 => std_logic_vector(to_unsigned(6,8) ,
72572	 => std_logic_vector(to_unsigned(8,8) ,
72573	 => std_logic_vector(to_unsigned(6,8) ,
72574	 => std_logic_vector(to_unsigned(9,8) ,
72575	 => std_logic_vector(to_unsigned(8,8) ,
72576	 => std_logic_vector(to_unsigned(8,8) ,
72577	 => std_logic_vector(to_unsigned(10,8) ,
72578	 => std_logic_vector(to_unsigned(10,8) ,
72579	 => std_logic_vector(to_unsigned(9,8) ,
72580	 => std_logic_vector(to_unsigned(8,8) ,
72581	 => std_logic_vector(to_unsigned(9,8) ,
72582	 => std_logic_vector(to_unsigned(8,8) ,
72583	 => std_logic_vector(to_unsigned(6,8) ,
72584	 => std_logic_vector(to_unsigned(8,8) ,
72585	 => std_logic_vector(to_unsigned(7,8) ,
72586	 => std_logic_vector(to_unsigned(7,8) ,
72587	 => std_logic_vector(to_unsigned(8,8) ,
72588	 => std_logic_vector(to_unsigned(12,8) ,
72589	 => std_logic_vector(to_unsigned(25,8) ,
72590	 => std_logic_vector(to_unsigned(19,8) ,
72591	 => std_logic_vector(to_unsigned(6,8) ,
72592	 => std_logic_vector(to_unsigned(8,8) ,
72593	 => std_logic_vector(to_unsigned(23,8) ,
72594	 => std_logic_vector(to_unsigned(46,8) ,
72595	 => std_logic_vector(to_unsigned(45,8) ,
72596	 => std_logic_vector(to_unsigned(21,8) ,
72597	 => std_logic_vector(to_unsigned(7,8) ,
72598	 => std_logic_vector(to_unsigned(0,8) ,
72599	 => std_logic_vector(to_unsigned(1,8) ,
72600	 => std_logic_vector(to_unsigned(30,8) ,
72601	 => std_logic_vector(to_unsigned(55,8) ,
72602	 => std_logic_vector(to_unsigned(10,8) ,
72603	 => std_logic_vector(to_unsigned(4,8) ,
72604	 => std_logic_vector(to_unsigned(35,8) ,
72605	 => std_logic_vector(to_unsigned(34,8) ,
72606	 => std_logic_vector(to_unsigned(30,8) ,
72607	 => std_logic_vector(to_unsigned(31,8) ,
72608	 => std_logic_vector(to_unsigned(19,8) ,
72609	 => std_logic_vector(to_unsigned(1,8) ,
72610	 => std_logic_vector(to_unsigned(0,8) ,
72611	 => std_logic_vector(to_unsigned(0,8) ,
72612	 => std_logic_vector(to_unsigned(0,8) ,
72613	 => std_logic_vector(to_unsigned(0,8) ,
72614	 => std_logic_vector(to_unsigned(1,8) ,
72615	 => std_logic_vector(to_unsigned(1,8) ,
72616	 => std_logic_vector(to_unsigned(0,8) ,
72617	 => std_logic_vector(to_unsigned(1,8) ,
72618	 => std_logic_vector(to_unsigned(3,8) ,
72619	 => std_logic_vector(to_unsigned(4,8) ,
72620	 => std_logic_vector(to_unsigned(1,8) ,
72621	 => std_logic_vector(to_unsigned(0,8) ,
72622	 => std_logic_vector(to_unsigned(1,8) ,
72623	 => std_logic_vector(to_unsigned(1,8) ,
72624	 => std_logic_vector(to_unsigned(0,8) ,
72625	 => std_logic_vector(to_unsigned(6,8) ,
72626	 => std_logic_vector(to_unsigned(34,8) ,
72627	 => std_logic_vector(to_unsigned(24,8) ,
72628	 => std_logic_vector(to_unsigned(25,8) ,
72629	 => std_logic_vector(to_unsigned(33,8) ,
72630	 => std_logic_vector(to_unsigned(58,8) ,
72631	 => std_logic_vector(to_unsigned(91,8) ,
72632	 => std_logic_vector(to_unsigned(59,8) ,
72633	 => std_logic_vector(to_unsigned(53,8) ,
72634	 => std_logic_vector(to_unsigned(67,8) ,
72635	 => std_logic_vector(to_unsigned(49,8) ,
72636	 => std_logic_vector(to_unsigned(49,8) ,
72637	 => std_logic_vector(to_unsigned(45,8) ,
72638	 => std_logic_vector(to_unsigned(45,8) ,
72639	 => std_logic_vector(to_unsigned(53,8) ,
72640	 => std_logic_vector(to_unsigned(71,8) ,
72641	 => std_logic_vector(to_unsigned(157,8) ,
72642	 => std_logic_vector(to_unsigned(131,8) ,
72643	 => std_logic_vector(to_unsigned(111,8) ,
72644	 => std_logic_vector(to_unsigned(112,8) ,
72645	 => std_logic_vector(to_unsigned(107,8) ,
72646	 => std_logic_vector(to_unsigned(109,8) ,
72647	 => std_logic_vector(to_unsigned(93,8) ,
72648	 => std_logic_vector(to_unsigned(79,8) ,
72649	 => std_logic_vector(to_unsigned(82,8) ,
72650	 => std_logic_vector(to_unsigned(88,8) ,
72651	 => std_logic_vector(to_unsigned(84,8) ,
72652	 => std_logic_vector(to_unsigned(91,8) ,
72653	 => std_logic_vector(to_unsigned(87,8) ,
72654	 => std_logic_vector(to_unsigned(81,8) ,
72655	 => std_logic_vector(to_unsigned(81,8) ,
72656	 => std_logic_vector(to_unsigned(74,8) ,
72657	 => std_logic_vector(to_unsigned(77,8) ,
72658	 => std_logic_vector(to_unsigned(79,8) ,
72659	 => std_logic_vector(to_unsigned(73,8) ,
72660	 => std_logic_vector(to_unsigned(67,8) ,
72661	 => std_logic_vector(to_unsigned(64,8) ,
72662	 => std_logic_vector(to_unsigned(59,8) ,
72663	 => std_logic_vector(to_unsigned(49,8) ,
72664	 => std_logic_vector(to_unsigned(45,8) ,
72665	 => std_logic_vector(to_unsigned(39,8) ,
72666	 => std_logic_vector(to_unsigned(40,8) ,
72667	 => std_logic_vector(to_unsigned(40,8) ,
72668	 => std_logic_vector(to_unsigned(43,8) ,
72669	 => std_logic_vector(to_unsigned(42,8) ,
72670	 => std_logic_vector(to_unsigned(76,8) ,
72671	 => std_logic_vector(to_unsigned(72,8) ,
72672	 => std_logic_vector(to_unsigned(28,8) ,
72673	 => std_logic_vector(to_unsigned(25,8) ,
72674	 => std_logic_vector(to_unsigned(18,8) ,
72675	 => std_logic_vector(to_unsigned(26,8) ,
72676	 => std_logic_vector(to_unsigned(33,8) ,
72677	 => std_logic_vector(to_unsigned(21,8) ,
72678	 => std_logic_vector(to_unsigned(20,8) ,
72679	 => std_logic_vector(to_unsigned(34,8) ,
72680	 => std_logic_vector(to_unsigned(25,8) ,
72681	 => std_logic_vector(to_unsigned(17,8) ,
72682	 => std_logic_vector(to_unsigned(16,8) ,
72683	 => std_logic_vector(to_unsigned(34,8) ,
72684	 => std_logic_vector(to_unsigned(30,8) ,
72685	 => std_logic_vector(to_unsigned(25,8) ,
72686	 => std_logic_vector(to_unsigned(34,8) ,
72687	 => std_logic_vector(to_unsigned(39,8) ,
72688	 => std_logic_vector(to_unsigned(42,8) ,
72689	 => std_logic_vector(to_unsigned(37,8) ,
72690	 => std_logic_vector(to_unsigned(31,8) ,
72691	 => std_logic_vector(to_unsigned(36,8) ,
72692	 => std_logic_vector(to_unsigned(33,8) ,
72693	 => std_logic_vector(to_unsigned(38,8) ,
72694	 => std_logic_vector(to_unsigned(42,8) ,
72695	 => std_logic_vector(to_unsigned(51,8) ,
72696	 => std_logic_vector(to_unsigned(56,8) ,
72697	 => std_logic_vector(to_unsigned(56,8) ,
72698	 => std_logic_vector(to_unsigned(47,8) ,
72699	 => std_logic_vector(to_unsigned(45,8) ,
72700	 => std_logic_vector(to_unsigned(44,8) ,
72701	 => std_logic_vector(to_unsigned(43,8) ,
72702	 => std_logic_vector(to_unsigned(48,8) ,
72703	 => std_logic_vector(to_unsigned(69,8) ,
72704	 => std_logic_vector(to_unsigned(91,8) ,
72705	 => std_logic_vector(to_unsigned(97,8) ,
72706	 => std_logic_vector(to_unsigned(87,8) ,
72707	 => std_logic_vector(to_unsigned(101,8) ,
72708	 => std_logic_vector(to_unsigned(73,8) ,
72709	 => std_logic_vector(to_unsigned(42,8) ,
72710	 => std_logic_vector(to_unsigned(49,8) ,
72711	 => std_logic_vector(to_unsigned(40,8) ,
72712	 => std_logic_vector(to_unsigned(36,8) ,
72713	 => std_logic_vector(to_unsigned(47,8) ,
72714	 => std_logic_vector(to_unsigned(66,8) ,
72715	 => std_logic_vector(to_unsigned(60,8) ,
72716	 => std_logic_vector(to_unsigned(52,8) ,
72717	 => std_logic_vector(to_unsigned(66,8) ,
72718	 => std_logic_vector(to_unsigned(67,8) ,
72719	 => std_logic_vector(to_unsigned(73,8) ,
72720	 => std_logic_vector(to_unsigned(68,8) ,
72721	 => std_logic_vector(to_unsigned(51,8) ,
72722	 => std_logic_vector(to_unsigned(60,8) ,
72723	 => std_logic_vector(to_unsigned(80,8) ,
72724	 => std_logic_vector(to_unsigned(88,8) ,
72725	 => std_logic_vector(to_unsigned(86,8) ,
72726	 => std_logic_vector(to_unsigned(74,8) ,
72727	 => std_logic_vector(to_unsigned(69,8) ,
72728	 => std_logic_vector(to_unsigned(51,8) ,
72729	 => std_logic_vector(to_unsigned(35,8) ,
72730	 => std_logic_vector(to_unsigned(45,8) ,
72731	 => std_logic_vector(to_unsigned(44,8) ,
72732	 => std_logic_vector(to_unsigned(35,8) ,
72733	 => std_logic_vector(to_unsigned(45,8) ,
72734	 => std_logic_vector(to_unsigned(52,8) ,
72735	 => std_logic_vector(to_unsigned(47,8) ,
72736	 => std_logic_vector(to_unsigned(33,8) ,
72737	 => std_logic_vector(to_unsigned(29,8) ,
72738	 => std_logic_vector(to_unsigned(34,8) ,
72739	 => std_logic_vector(to_unsigned(29,8) ,
72740	 => std_logic_vector(to_unsigned(23,8) ,
72741	 => std_logic_vector(to_unsigned(36,8) ,
72742	 => std_logic_vector(to_unsigned(38,8) ,
72743	 => std_logic_vector(to_unsigned(40,8) ,
72744	 => std_logic_vector(to_unsigned(108,8) ,
72745	 => std_logic_vector(to_unsigned(114,8) ,
72746	 => std_logic_vector(to_unsigned(100,8) ,
72747	 => std_logic_vector(to_unsigned(104,8) ,
72748	 => std_logic_vector(to_unsigned(100,8) ,
72749	 => std_logic_vector(to_unsigned(100,8) ,
72750	 => std_logic_vector(to_unsigned(96,8) ,
72751	 => std_logic_vector(to_unsigned(91,8) ,
72752	 => std_logic_vector(to_unsigned(84,8) ,
72753	 => std_logic_vector(to_unsigned(64,8) ,
72754	 => std_logic_vector(to_unsigned(64,8) ,
72755	 => std_logic_vector(to_unsigned(61,8) ,
72756	 => std_logic_vector(to_unsigned(72,8) ,
72757	 => std_logic_vector(to_unsigned(121,8) ,
72758	 => std_logic_vector(to_unsigned(124,8) ,
72759	 => std_logic_vector(to_unsigned(118,8) ,
72760	 => std_logic_vector(to_unsigned(109,8) ,
72761	 => std_logic_vector(to_unsigned(104,8) ,
72762	 => std_logic_vector(to_unsigned(105,8) ,
72763	 => std_logic_vector(to_unsigned(95,8) ,
72764	 => std_logic_vector(to_unsigned(90,8) ,
72765	 => std_logic_vector(to_unsigned(84,8) ,
72766	 => std_logic_vector(to_unsigned(87,8) ,
72767	 => std_logic_vector(to_unsigned(91,8) ,
72768	 => std_logic_vector(to_unsigned(69,8) ,
72769	 => std_logic_vector(to_unsigned(45,8) ,
72770	 => std_logic_vector(to_unsigned(45,8) ,
72771	 => std_logic_vector(to_unsigned(35,8) ,
72772	 => std_logic_vector(to_unsigned(37,8) ,
72773	 => std_logic_vector(to_unsigned(68,8) ,
72774	 => std_logic_vector(to_unsigned(80,8) ,
72775	 => std_logic_vector(to_unsigned(84,8) ,
72776	 => std_logic_vector(to_unsigned(78,8) ,
72777	 => std_logic_vector(to_unsigned(52,8) ,
72778	 => std_logic_vector(to_unsigned(46,8) ,
72779	 => std_logic_vector(to_unsigned(57,8) ,
72780	 => std_logic_vector(to_unsigned(53,8) ,
72781	 => std_logic_vector(to_unsigned(45,8) ,
72782	 => std_logic_vector(to_unsigned(45,8) ,
72783	 => std_logic_vector(to_unsigned(25,8) ,
72784	 => std_logic_vector(to_unsigned(32,8) ,
72785	 => std_logic_vector(to_unsigned(28,8) ,
72786	 => std_logic_vector(to_unsigned(25,8) ,
72787	 => std_logic_vector(to_unsigned(46,8) ,
72788	 => std_logic_vector(to_unsigned(31,8) ,
72789	 => std_logic_vector(to_unsigned(51,8) ,
72790	 => std_logic_vector(to_unsigned(100,8) ,
72791	 => std_logic_vector(to_unsigned(92,8) ,
72792	 => std_logic_vector(to_unsigned(80,8) ,
72793	 => std_logic_vector(to_unsigned(72,8) ,
72794	 => std_logic_vector(to_unsigned(80,8) ,
72795	 => std_logic_vector(to_unsigned(97,8) ,
72796	 => std_logic_vector(to_unsigned(92,8) ,
72797	 => std_logic_vector(to_unsigned(74,8) ,
72798	 => std_logic_vector(to_unsigned(73,8) ,
72799	 => std_logic_vector(to_unsigned(80,8) ,
72800	 => std_logic_vector(to_unsigned(78,8) ,
72801	 => std_logic_vector(to_unsigned(45,8) ,
72802	 => std_logic_vector(to_unsigned(25,8) ,
72803	 => std_logic_vector(to_unsigned(27,8) ,
72804	 => std_logic_vector(to_unsigned(28,8) ,
72805	 => std_logic_vector(to_unsigned(37,8) ,
72806	 => std_logic_vector(to_unsigned(31,8) ,
72807	 => std_logic_vector(to_unsigned(4,8) ,
72808	 => std_logic_vector(to_unsigned(4,8) ,
72809	 => std_logic_vector(to_unsigned(10,8) ,
72810	 => std_logic_vector(to_unsigned(18,8) ,
72811	 => std_logic_vector(to_unsigned(37,8) ,
72812	 => std_logic_vector(to_unsigned(18,8) ,
72813	 => std_logic_vector(to_unsigned(19,8) ,
72814	 => std_logic_vector(to_unsigned(16,8) ,
72815	 => std_logic_vector(to_unsigned(14,8) ,
72816	 => std_logic_vector(to_unsigned(37,8) ,
72817	 => std_logic_vector(to_unsigned(37,8) ,
72818	 => std_logic_vector(to_unsigned(45,8) ,
72819	 => std_logic_vector(to_unsigned(72,8) ,
72820	 => std_logic_vector(to_unsigned(64,8) ,
72821	 => std_logic_vector(to_unsigned(20,8) ,
72822	 => std_logic_vector(to_unsigned(8,8) ,
72823	 => std_logic_vector(to_unsigned(14,8) ,
72824	 => std_logic_vector(to_unsigned(10,8) ,
72825	 => std_logic_vector(to_unsigned(10,8) ,
72826	 => std_logic_vector(to_unsigned(22,8) ,
72827	 => std_logic_vector(to_unsigned(41,8) ,
72828	 => std_logic_vector(to_unsigned(43,8) ,
72829	 => std_logic_vector(to_unsigned(40,8) ,
72830	 => std_logic_vector(to_unsigned(25,8) ,
72831	 => std_logic_vector(to_unsigned(25,8) ,
72832	 => std_logic_vector(to_unsigned(35,8) ,
72833	 => std_logic_vector(to_unsigned(45,8) ,
72834	 => std_logic_vector(to_unsigned(41,8) ,
72835	 => std_logic_vector(to_unsigned(25,8) ,
72836	 => std_logic_vector(to_unsigned(23,8) ,
72837	 => std_logic_vector(to_unsigned(22,8) ,
72838	 => std_logic_vector(to_unsigned(27,8) ,
72839	 => std_logic_vector(to_unsigned(29,8) ,
72840	 => std_logic_vector(to_unsigned(29,8) ,
72841	 => std_logic_vector(to_unsigned(17,8) ,
72842	 => std_logic_vector(to_unsigned(10,8) ,
72843	 => std_logic_vector(to_unsigned(12,8) ,
72844	 => std_logic_vector(to_unsigned(13,8) ,
72845	 => std_logic_vector(to_unsigned(13,8) ,
72846	 => std_logic_vector(to_unsigned(8,8) ,
72847	 => std_logic_vector(to_unsigned(8,8) ,
72848	 => std_logic_vector(to_unsigned(23,8) ,
72849	 => std_logic_vector(to_unsigned(14,8) ,
72850	 => std_logic_vector(to_unsigned(5,8) ,
72851	 => std_logic_vector(to_unsigned(8,8) ,
72852	 => std_logic_vector(to_unsigned(20,8) ,
72853	 => std_logic_vector(to_unsigned(20,8) ,
72854	 => std_logic_vector(to_unsigned(23,8) ,
72855	 => std_logic_vector(to_unsigned(30,8) ,
72856	 => std_logic_vector(to_unsigned(29,8) ,
72857	 => std_logic_vector(to_unsigned(18,8) ,
72858	 => std_logic_vector(to_unsigned(17,8) ,
72859	 => std_logic_vector(to_unsigned(24,8) ,
72860	 => std_logic_vector(to_unsigned(37,8) ,
72861	 => std_logic_vector(to_unsigned(32,8) ,
72862	 => std_logic_vector(to_unsigned(20,8) ,
72863	 => std_logic_vector(to_unsigned(22,8) ,
72864	 => std_logic_vector(to_unsigned(25,8) ,
72865	 => std_logic_vector(to_unsigned(27,8) ,
72866	 => std_logic_vector(to_unsigned(25,8) ,
72867	 => std_logic_vector(to_unsigned(22,8) ,
72868	 => std_logic_vector(to_unsigned(12,8) ,
72869	 => std_logic_vector(to_unsigned(3,8) ,
72870	 => std_logic_vector(to_unsigned(14,8) ,
72871	 => std_logic_vector(to_unsigned(24,8) ,
72872	 => std_logic_vector(to_unsigned(15,8) ,
72873	 => std_logic_vector(to_unsigned(11,8) ,
72874	 => std_logic_vector(to_unsigned(24,8) ,
72875	 => std_logic_vector(to_unsigned(36,8) ,
72876	 => std_logic_vector(to_unsigned(5,8) ,
72877	 => std_logic_vector(to_unsigned(7,8) ,
72878	 => std_logic_vector(to_unsigned(45,8) ,
72879	 => std_logic_vector(to_unsigned(45,8) ,
72880	 => std_logic_vector(to_unsigned(11,8) ,
72881	 => std_logic_vector(to_unsigned(5,8) ,
72882	 => std_logic_vector(to_unsigned(25,8) ,
72883	 => std_logic_vector(to_unsigned(62,8) ,
72884	 => std_logic_vector(to_unsigned(101,8) ,
72885	 => std_logic_vector(to_unsigned(96,8) ,
72886	 => std_logic_vector(to_unsigned(39,8) ,
72887	 => std_logic_vector(to_unsigned(77,8) ,
72888	 => std_logic_vector(to_unsigned(122,8) ,
72889	 => std_logic_vector(to_unsigned(90,8) ,
72890	 => std_logic_vector(to_unsigned(12,8) ,
72891	 => std_logic_vector(to_unsigned(6,8) ,
72892	 => std_logic_vector(to_unsigned(6,8) ,
72893	 => std_logic_vector(to_unsigned(6,8) ,
72894	 => std_logic_vector(to_unsigned(9,8) ,
72895	 => std_logic_vector(to_unsigned(8,8) ,
72896	 => std_logic_vector(to_unsigned(8,8) ,
72897	 => std_logic_vector(to_unsigned(7,8) ,
72898	 => std_logic_vector(to_unsigned(9,8) ,
72899	 => std_logic_vector(to_unsigned(8,8) ,
72900	 => std_logic_vector(to_unsigned(8,8) ,
72901	 => std_logic_vector(to_unsigned(10,8) ,
72902	 => std_logic_vector(to_unsigned(9,8) ,
72903	 => std_logic_vector(to_unsigned(8,8) ,
72904	 => std_logic_vector(to_unsigned(9,8) ,
72905	 => std_logic_vector(to_unsigned(9,8) ,
72906	 => std_logic_vector(to_unsigned(9,8) ,
72907	 => std_logic_vector(to_unsigned(7,8) ,
72908	 => std_logic_vector(to_unsigned(10,8) ,
72909	 => std_logic_vector(to_unsigned(28,8) ,
72910	 => std_logic_vector(to_unsigned(23,8) ,
72911	 => std_logic_vector(to_unsigned(8,8) ,
72912	 => std_logic_vector(to_unsigned(8,8) ,
72913	 => std_logic_vector(to_unsigned(13,8) ,
72914	 => std_logic_vector(to_unsigned(26,8) ,
72915	 => std_logic_vector(to_unsigned(22,8) ,
72916	 => std_logic_vector(to_unsigned(14,8) ,
72917	 => std_logic_vector(to_unsigned(11,8) ,
72918	 => std_logic_vector(to_unsigned(1,8) ,
72919	 => std_logic_vector(to_unsigned(0,8) ,
72920	 => std_logic_vector(to_unsigned(10,8) ,
72921	 => std_logic_vector(to_unsigned(48,8) ,
72922	 => std_logic_vector(to_unsigned(6,8) ,
72923	 => std_logic_vector(to_unsigned(6,8) ,
72924	 => std_logic_vector(to_unsigned(41,8) ,
72925	 => std_logic_vector(to_unsigned(35,8) ,
72926	 => std_logic_vector(to_unsigned(35,8) ,
72927	 => std_logic_vector(to_unsigned(35,8) ,
72928	 => std_logic_vector(to_unsigned(41,8) ,
72929	 => std_logic_vector(to_unsigned(17,8) ,
72930	 => std_logic_vector(to_unsigned(1,8) ,
72931	 => std_logic_vector(to_unsigned(0,8) ,
72932	 => std_logic_vector(to_unsigned(0,8) ,
72933	 => std_logic_vector(to_unsigned(1,8) ,
72934	 => std_logic_vector(to_unsigned(4,8) ,
72935	 => std_logic_vector(to_unsigned(4,8) ,
72936	 => std_logic_vector(to_unsigned(4,8) ,
72937	 => std_logic_vector(to_unsigned(3,8) ,
72938	 => std_logic_vector(to_unsigned(1,8) ,
72939	 => std_logic_vector(to_unsigned(2,8) ,
72940	 => std_logic_vector(to_unsigned(1,8) ,
72941	 => std_logic_vector(to_unsigned(0,8) ,
72942	 => std_logic_vector(to_unsigned(0,8) ,
72943	 => std_logic_vector(to_unsigned(0,8) ,
72944	 => std_logic_vector(to_unsigned(0,8) ,
72945	 => std_logic_vector(to_unsigned(18,8) ,
72946	 => std_logic_vector(to_unsigned(47,8) ,
72947	 => std_logic_vector(to_unsigned(30,8) ,
72948	 => std_logic_vector(to_unsigned(25,8) ,
72949	 => std_logic_vector(to_unsigned(34,8) ,
72950	 => std_logic_vector(to_unsigned(38,8) ,
72951	 => std_logic_vector(to_unsigned(46,8) ,
72952	 => std_logic_vector(to_unsigned(57,8) ,
72953	 => std_logic_vector(to_unsigned(61,8) ,
72954	 => std_logic_vector(to_unsigned(62,8) ,
72955	 => std_logic_vector(to_unsigned(39,8) ,
72956	 => std_logic_vector(to_unsigned(21,8) ,
72957	 => std_logic_vector(to_unsigned(25,8) ,
72958	 => std_logic_vector(to_unsigned(31,8) ,
72959	 => std_logic_vector(to_unsigned(29,8) ,
72960	 => std_logic_vector(to_unsigned(30,8) ,
72961	 => std_logic_vector(to_unsigned(138,8) ,
72962	 => std_logic_vector(to_unsigned(116,8) ,
72963	 => std_logic_vector(to_unsigned(99,8) ,
72964	 => std_logic_vector(to_unsigned(109,8) ,
72965	 => std_logic_vector(to_unsigned(108,8) ,
72966	 => std_logic_vector(to_unsigned(103,8) ,
72967	 => std_logic_vector(to_unsigned(91,8) ,
72968	 => std_logic_vector(to_unsigned(86,8) ,
72969	 => std_logic_vector(to_unsigned(92,8) ,
72970	 => std_logic_vector(to_unsigned(87,8) ,
72971	 => std_logic_vector(to_unsigned(90,8) ,
72972	 => std_logic_vector(to_unsigned(86,8) ,
72973	 => std_logic_vector(to_unsigned(84,8) ,
72974	 => std_logic_vector(to_unsigned(84,8) ,
72975	 => std_logic_vector(to_unsigned(84,8) ,
72976	 => std_logic_vector(to_unsigned(82,8) ,
72977	 => std_logic_vector(to_unsigned(79,8) ,
72978	 => std_logic_vector(to_unsigned(76,8) ,
72979	 => std_logic_vector(to_unsigned(72,8) ,
72980	 => std_logic_vector(to_unsigned(66,8) ,
72981	 => std_logic_vector(to_unsigned(57,8) ,
72982	 => std_logic_vector(to_unsigned(59,8) ,
72983	 => std_logic_vector(to_unsigned(51,8) ,
72984	 => std_logic_vector(to_unsigned(45,8) ,
72985	 => std_logic_vector(to_unsigned(25,8) ,
72986	 => std_logic_vector(to_unsigned(27,8) ,
72987	 => std_logic_vector(to_unsigned(40,8) ,
72988	 => std_logic_vector(to_unsigned(41,8) ,
72989	 => std_logic_vector(to_unsigned(42,8) ,
72990	 => std_logic_vector(to_unsigned(67,8) ,
72991	 => std_logic_vector(to_unsigned(59,8) ,
72992	 => std_logic_vector(to_unsigned(33,8) ,
72993	 => std_logic_vector(to_unsigned(45,8) ,
72994	 => std_logic_vector(to_unsigned(50,8) ,
72995	 => std_logic_vector(to_unsigned(56,8) ,
72996	 => std_logic_vector(to_unsigned(67,8) ,
72997	 => std_logic_vector(to_unsigned(45,8) ,
72998	 => std_logic_vector(to_unsigned(38,8) ,
72999	 => std_logic_vector(to_unsigned(29,8) ,
73000	 => std_logic_vector(to_unsigned(28,8) ,
73001	 => std_logic_vector(to_unsigned(20,8) ,
73002	 => std_logic_vector(to_unsigned(10,8) ,
73003	 => std_logic_vector(to_unsigned(22,8) ,
73004	 => std_logic_vector(to_unsigned(25,8) ,
73005	 => std_logic_vector(to_unsigned(32,8) ,
73006	 => std_logic_vector(to_unsigned(30,8) ,
73007	 => std_logic_vector(to_unsigned(29,8) ,
73008	 => std_logic_vector(to_unsigned(29,8) ,
73009	 => std_logic_vector(to_unsigned(36,8) ,
73010	 => std_logic_vector(to_unsigned(35,8) ,
73011	 => std_logic_vector(to_unsigned(40,8) ,
73012	 => std_logic_vector(to_unsigned(41,8) ,
73013	 => std_logic_vector(to_unsigned(37,8) ,
73014	 => std_logic_vector(to_unsigned(41,8) ,
73015	 => std_logic_vector(to_unsigned(61,8) ,
73016	 => std_logic_vector(to_unsigned(85,8) ,
73017	 => std_logic_vector(to_unsigned(96,8) ,
73018	 => std_logic_vector(to_unsigned(86,8) ,
73019	 => std_logic_vector(to_unsigned(77,8) ,
73020	 => std_logic_vector(to_unsigned(68,8) ,
73021	 => std_logic_vector(to_unsigned(70,8) ,
73022	 => std_logic_vector(to_unsigned(91,8) ,
73023	 => std_logic_vector(to_unsigned(103,8) ,
73024	 => std_logic_vector(to_unsigned(97,8) ,
73025	 => std_logic_vector(to_unsigned(96,8) ,
73026	 => std_logic_vector(to_unsigned(105,8) ,
73027	 => std_logic_vector(to_unsigned(131,8) ,
73028	 => std_logic_vector(to_unsigned(78,8) ,
73029	 => std_logic_vector(to_unsigned(39,8) ,
73030	 => std_logic_vector(to_unsigned(44,8) ,
73031	 => std_logic_vector(to_unsigned(40,8) ,
73032	 => std_logic_vector(to_unsigned(33,8) ,
73033	 => std_logic_vector(to_unsigned(45,8) ,
73034	 => std_logic_vector(to_unsigned(64,8) ,
73035	 => std_logic_vector(to_unsigned(55,8) ,
73036	 => std_logic_vector(to_unsigned(58,8) ,
73037	 => std_logic_vector(to_unsigned(65,8) ,
73038	 => std_logic_vector(to_unsigned(69,8) ,
73039	 => std_logic_vector(to_unsigned(52,8) ,
73040	 => std_logic_vector(to_unsigned(37,8) ,
73041	 => std_logic_vector(to_unsigned(52,8) ,
73042	 => std_logic_vector(to_unsigned(86,8) ,
73043	 => std_logic_vector(to_unsigned(93,8) ,
73044	 => std_logic_vector(to_unsigned(90,8) ,
73045	 => std_logic_vector(to_unsigned(101,8) ,
73046	 => std_logic_vector(to_unsigned(72,8) ,
73047	 => std_logic_vector(to_unsigned(41,8) ,
73048	 => std_logic_vector(to_unsigned(51,8) ,
73049	 => std_logic_vector(to_unsigned(49,8) ,
73050	 => std_logic_vector(to_unsigned(54,8) ,
73051	 => std_logic_vector(to_unsigned(39,8) ,
73052	 => std_logic_vector(to_unsigned(45,8) ,
73053	 => std_logic_vector(to_unsigned(90,8) ,
73054	 => std_logic_vector(to_unsigned(70,8) ,
73055	 => std_logic_vector(to_unsigned(39,8) ,
73056	 => std_logic_vector(to_unsigned(32,8) ,
73057	 => std_logic_vector(to_unsigned(30,8) ,
73058	 => std_logic_vector(to_unsigned(30,8) ,
73059	 => std_logic_vector(to_unsigned(30,8) ,
73060	 => std_logic_vector(to_unsigned(29,8) ,
73061	 => std_logic_vector(to_unsigned(41,8) ,
73062	 => std_logic_vector(to_unsigned(34,8) ,
73063	 => std_logic_vector(to_unsigned(43,8) ,
73064	 => std_logic_vector(to_unsigned(95,8) ,
73065	 => std_logic_vector(to_unsigned(65,8) ,
73066	 => std_logic_vector(to_unsigned(109,8) ,
73067	 => std_logic_vector(to_unsigned(133,8) ,
73068	 => std_logic_vector(to_unsigned(92,8) ,
73069	 => std_logic_vector(to_unsigned(122,8) ,
73070	 => std_logic_vector(to_unsigned(118,8) ,
73071	 => std_logic_vector(to_unsigned(90,8) ,
73072	 => std_logic_vector(to_unsigned(95,8) ,
73073	 => std_logic_vector(to_unsigned(74,8) ,
73074	 => std_logic_vector(to_unsigned(79,8) ,
73075	 => std_logic_vector(to_unsigned(77,8) ,
73076	 => std_logic_vector(to_unsigned(91,8) ,
73077	 => std_logic_vector(to_unsigned(118,8) ,
73078	 => std_logic_vector(to_unsigned(116,8) ,
73079	 => std_logic_vector(to_unsigned(122,8) ,
73080	 => std_logic_vector(to_unsigned(119,8) ,
73081	 => std_logic_vector(to_unsigned(114,8) ,
73082	 => std_logic_vector(to_unsigned(109,8) ,
73083	 => std_logic_vector(to_unsigned(99,8) ,
73084	 => std_logic_vector(to_unsigned(90,8) ,
73085	 => std_logic_vector(to_unsigned(82,8) ,
73086	 => std_logic_vector(to_unsigned(90,8) ,
73087	 => std_logic_vector(to_unsigned(90,8) ,
73088	 => std_logic_vector(to_unsigned(88,8) ,
73089	 => std_logic_vector(to_unsigned(86,8) ,
73090	 => std_logic_vector(to_unsigned(93,8) ,
73091	 => std_logic_vector(to_unsigned(105,8) ,
73092	 => std_logic_vector(to_unsigned(107,8) ,
73093	 => std_logic_vector(to_unsigned(95,8) ,
73094	 => std_logic_vector(to_unsigned(101,8) ,
73095	 => std_logic_vector(to_unsigned(97,8) ,
73096	 => std_logic_vector(to_unsigned(79,8) ,
73097	 => std_logic_vector(to_unsigned(53,8) ,
73098	 => std_logic_vector(to_unsigned(41,8) ,
73099	 => std_logic_vector(to_unsigned(49,8) ,
73100	 => std_logic_vector(to_unsigned(51,8) ,
73101	 => std_logic_vector(to_unsigned(56,8) ,
73102	 => std_logic_vector(to_unsigned(55,8) ,
73103	 => std_logic_vector(to_unsigned(55,8) ,
73104	 => std_logic_vector(to_unsigned(55,8) ,
73105	 => std_logic_vector(to_unsigned(45,8) ,
73106	 => std_logic_vector(to_unsigned(28,8) ,
73107	 => std_logic_vector(to_unsigned(35,8) ,
73108	 => std_logic_vector(to_unsigned(15,8) ,
73109	 => std_logic_vector(to_unsigned(25,8) ,
73110	 => std_logic_vector(to_unsigned(97,8) ,
73111	 => std_logic_vector(to_unsigned(114,8) ,
73112	 => std_logic_vector(to_unsigned(112,8) ,
73113	 => std_logic_vector(to_unsigned(107,8) ,
73114	 => std_logic_vector(to_unsigned(100,8) ,
73115	 => std_logic_vector(to_unsigned(93,8) ,
73116	 => std_logic_vector(to_unsigned(88,8) ,
73117	 => std_logic_vector(to_unsigned(85,8) ,
73118	 => std_logic_vector(to_unsigned(72,8) ,
73119	 => std_logic_vector(to_unsigned(62,8) ,
73120	 => std_logic_vector(to_unsigned(55,8) ,
73121	 => std_logic_vector(to_unsigned(22,8) ,
73122	 => std_logic_vector(to_unsigned(36,8) ,
73123	 => std_logic_vector(to_unsigned(32,8) ,
73124	 => std_logic_vector(to_unsigned(20,8) ,
73125	 => std_logic_vector(to_unsigned(31,8) ,
73126	 => std_logic_vector(to_unsigned(32,8) ,
73127	 => std_logic_vector(to_unsigned(6,8) ,
73128	 => std_logic_vector(to_unsigned(5,8) ,
73129	 => std_logic_vector(to_unsigned(10,8) ,
73130	 => std_logic_vector(to_unsigned(17,8) ,
73131	 => std_logic_vector(to_unsigned(22,8) ,
73132	 => std_logic_vector(to_unsigned(18,8) ,
73133	 => std_logic_vector(to_unsigned(20,8) ,
73134	 => std_logic_vector(to_unsigned(17,8) ,
73135	 => std_logic_vector(to_unsigned(28,8) ,
73136	 => std_logic_vector(to_unsigned(27,8) ,
73137	 => std_logic_vector(to_unsigned(35,8) ,
73138	 => std_logic_vector(to_unsigned(62,8) ,
73139	 => std_logic_vector(to_unsigned(45,8) ,
73140	 => std_logic_vector(to_unsigned(36,8) ,
73141	 => std_logic_vector(to_unsigned(24,8) ,
73142	 => std_logic_vector(to_unsigned(12,8) ,
73143	 => std_logic_vector(to_unsigned(14,8) ,
73144	 => std_logic_vector(to_unsigned(12,8) ,
73145	 => std_logic_vector(to_unsigned(10,8) ,
73146	 => std_logic_vector(to_unsigned(23,8) ,
73147	 => std_logic_vector(to_unsigned(44,8) ,
73148	 => std_logic_vector(to_unsigned(51,8) ,
73149	 => std_logic_vector(to_unsigned(41,8) ,
73150	 => std_logic_vector(to_unsigned(27,8) ,
73151	 => std_logic_vector(to_unsigned(32,8) ,
73152	 => std_logic_vector(to_unsigned(32,8) ,
73153	 => std_logic_vector(to_unsigned(27,8) ,
73154	 => std_logic_vector(to_unsigned(29,8) ,
73155	 => std_logic_vector(to_unsigned(24,8) ,
73156	 => std_logic_vector(to_unsigned(22,8) ,
73157	 => std_logic_vector(to_unsigned(30,8) ,
73158	 => std_logic_vector(to_unsigned(45,8) ,
73159	 => std_logic_vector(to_unsigned(45,8) ,
73160	 => std_logic_vector(to_unsigned(32,8) ,
73161	 => std_logic_vector(to_unsigned(21,8) ,
73162	 => std_logic_vector(to_unsigned(12,8) ,
73163	 => std_logic_vector(to_unsigned(8,8) ,
73164	 => std_logic_vector(to_unsigned(18,8) ,
73165	 => std_logic_vector(to_unsigned(19,8) ,
73166	 => std_logic_vector(to_unsigned(9,8) ,
73167	 => std_logic_vector(to_unsigned(9,8) ,
73168	 => std_logic_vector(to_unsigned(25,8) ,
73169	 => std_logic_vector(to_unsigned(31,8) ,
73170	 => std_logic_vector(to_unsigned(25,8) ,
73171	 => std_logic_vector(to_unsigned(20,8) ,
73172	 => std_logic_vector(to_unsigned(19,8) ,
73173	 => std_logic_vector(to_unsigned(21,8) ,
73174	 => std_logic_vector(to_unsigned(37,8) ,
73175	 => std_logic_vector(to_unsigned(62,8) ,
73176	 => std_logic_vector(to_unsigned(47,8) ,
73177	 => std_logic_vector(to_unsigned(20,8) ,
73178	 => std_logic_vector(to_unsigned(16,8) ,
73179	 => std_logic_vector(to_unsigned(24,8) ,
73180	 => std_logic_vector(to_unsigned(37,8) ,
73181	 => std_logic_vector(to_unsigned(38,8) ,
73182	 => std_logic_vector(to_unsigned(23,8) ,
73183	 => std_logic_vector(to_unsigned(22,8) ,
73184	 => std_logic_vector(to_unsigned(28,8) ,
73185	 => std_logic_vector(to_unsigned(25,8) ,
73186	 => std_logic_vector(to_unsigned(30,8) ,
73187	 => std_logic_vector(to_unsigned(37,8) ,
73188	 => std_logic_vector(to_unsigned(14,8) ,
73189	 => std_logic_vector(to_unsigned(3,8) ,
73190	 => std_logic_vector(to_unsigned(15,8) ,
73191	 => std_logic_vector(to_unsigned(35,8) ,
73192	 => std_logic_vector(to_unsigned(28,8) ,
73193	 => std_logic_vector(to_unsigned(24,8) ,
73194	 => std_logic_vector(to_unsigned(34,8) ,
73195	 => std_logic_vector(to_unsigned(35,8) ,
73196	 => std_logic_vector(to_unsigned(11,8) ,
73197	 => std_logic_vector(to_unsigned(9,8) ,
73198	 => std_logic_vector(to_unsigned(41,8) ,
73199	 => std_logic_vector(to_unsigned(45,8) ,
73200	 => std_logic_vector(to_unsigned(17,8) ,
73201	 => std_logic_vector(to_unsigned(5,8) ,
73202	 => std_logic_vector(to_unsigned(30,8) ,
73203	 => std_logic_vector(to_unsigned(51,8) ,
73204	 => std_logic_vector(to_unsigned(63,8) ,
73205	 => std_logic_vector(to_unsigned(71,8) ,
73206	 => std_logic_vector(to_unsigned(37,8) ,
73207	 => std_logic_vector(to_unsigned(81,8) ,
73208	 => std_logic_vector(to_unsigned(128,8) ,
73209	 => std_logic_vector(to_unsigned(61,8) ,
73210	 => std_logic_vector(to_unsigned(8,8) ,
73211	 => std_logic_vector(to_unsigned(8,8) ,
73212	 => std_logic_vector(to_unsigned(8,8) ,
73213	 => std_logic_vector(to_unsigned(8,8) ,
73214	 => std_logic_vector(to_unsigned(9,8) ,
73215	 => std_logic_vector(to_unsigned(8,8) ,
73216	 => std_logic_vector(to_unsigned(9,8) ,
73217	 => std_logic_vector(to_unsigned(10,8) ,
73218	 => std_logic_vector(to_unsigned(12,8) ,
73219	 => std_logic_vector(to_unsigned(9,8) ,
73220	 => std_logic_vector(to_unsigned(6,8) ,
73221	 => std_logic_vector(to_unsigned(7,8) ,
73222	 => std_logic_vector(to_unsigned(6,8) ,
73223	 => std_logic_vector(to_unsigned(7,8) ,
73224	 => std_logic_vector(to_unsigned(10,8) ,
73225	 => std_logic_vector(to_unsigned(12,8) ,
73226	 => std_logic_vector(to_unsigned(11,8) ,
73227	 => std_logic_vector(to_unsigned(12,8) ,
73228	 => std_logic_vector(to_unsigned(15,8) ,
73229	 => std_logic_vector(to_unsigned(24,8) ,
73230	 => std_logic_vector(to_unsigned(20,8) ,
73231	 => std_logic_vector(to_unsigned(9,8) ,
73232	 => std_logic_vector(to_unsigned(9,8) ,
73233	 => std_logic_vector(to_unsigned(9,8) ,
73234	 => std_logic_vector(to_unsigned(23,8) ,
73235	 => std_logic_vector(to_unsigned(23,8) ,
73236	 => std_logic_vector(to_unsigned(14,8) ,
73237	 => std_logic_vector(to_unsigned(22,8) ,
73238	 => std_logic_vector(to_unsigned(4,8) ,
73239	 => std_logic_vector(to_unsigned(0,8) ,
73240	 => std_logic_vector(to_unsigned(3,8) ,
73241	 => std_logic_vector(to_unsigned(37,8) ,
73242	 => std_logic_vector(to_unsigned(10,8) ,
73243	 => std_logic_vector(to_unsigned(17,8) ,
73244	 => std_logic_vector(to_unsigned(40,8) ,
73245	 => std_logic_vector(to_unsigned(32,8) ,
73246	 => std_logic_vector(to_unsigned(29,8) ,
73247	 => std_logic_vector(to_unsigned(30,8) ,
73248	 => std_logic_vector(to_unsigned(33,8) ,
73249	 => std_logic_vector(to_unsigned(46,8) ,
73250	 => std_logic_vector(to_unsigned(8,8) ,
73251	 => std_logic_vector(to_unsigned(0,8) ,
73252	 => std_logic_vector(to_unsigned(0,8) ,
73253	 => std_logic_vector(to_unsigned(1,8) ,
73254	 => std_logic_vector(to_unsigned(1,8) ,
73255	 => std_logic_vector(to_unsigned(2,8) ,
73256	 => std_logic_vector(to_unsigned(3,8) ,
73257	 => std_logic_vector(to_unsigned(5,8) ,
73258	 => std_logic_vector(to_unsigned(3,8) ,
73259	 => std_logic_vector(to_unsigned(1,8) ,
73260	 => std_logic_vector(to_unsigned(2,8) ,
73261	 => std_logic_vector(to_unsigned(0,8) ,
73262	 => std_logic_vector(to_unsigned(1,8) ,
73263	 => std_logic_vector(to_unsigned(0,8) ,
73264	 => std_logic_vector(to_unsigned(2,8) ,
73265	 => std_logic_vector(to_unsigned(27,8) ,
73266	 => std_logic_vector(to_unsigned(34,8) ,
73267	 => std_logic_vector(to_unsigned(30,8) ,
73268	 => std_logic_vector(to_unsigned(28,8) ,
73269	 => std_logic_vector(to_unsigned(33,8) ,
73270	 => std_logic_vector(to_unsigned(57,8) ,
73271	 => std_logic_vector(to_unsigned(64,8) ,
73272	 => std_logic_vector(to_unsigned(69,8) ,
73273	 => std_logic_vector(to_unsigned(68,8) ,
73274	 => std_logic_vector(to_unsigned(37,8) ,
73275	 => std_logic_vector(to_unsigned(35,8) ,
73276	 => std_logic_vector(to_unsigned(45,8) ,
73277	 => std_logic_vector(to_unsigned(39,8) ,
73278	 => std_logic_vector(to_unsigned(38,8) ,
73279	 => std_logic_vector(to_unsigned(35,8) ,
73280	 => std_logic_vector(to_unsigned(22,8) ,
73281	 => std_logic_vector(to_unsigned(108,8) ,
73282	 => std_logic_vector(to_unsigned(112,8) ,
73283	 => std_logic_vector(to_unsigned(116,8) ,
73284	 => std_logic_vector(to_unsigned(100,8) ,
73285	 => std_logic_vector(to_unsigned(99,8) ,
73286	 => std_logic_vector(to_unsigned(101,8) ,
73287	 => std_logic_vector(to_unsigned(96,8) ,
73288	 => std_logic_vector(to_unsigned(96,8) ,
73289	 => std_logic_vector(to_unsigned(101,8) ,
73290	 => std_logic_vector(to_unsigned(96,8) ,
73291	 => std_logic_vector(to_unsigned(107,8) ,
73292	 => std_logic_vector(to_unsigned(85,8) ,
73293	 => std_logic_vector(to_unsigned(80,8) ,
73294	 => std_logic_vector(to_unsigned(85,8) ,
73295	 => std_logic_vector(to_unsigned(85,8) ,
73296	 => std_logic_vector(to_unsigned(84,8) ,
73297	 => std_logic_vector(to_unsigned(81,8) ,
73298	 => std_logic_vector(to_unsigned(76,8) ,
73299	 => std_logic_vector(to_unsigned(73,8) ,
73300	 => std_logic_vector(to_unsigned(64,8) ,
73301	 => std_logic_vector(to_unsigned(57,8) ,
73302	 => std_logic_vector(to_unsigned(50,8) ,
73303	 => std_logic_vector(to_unsigned(45,8) ,
73304	 => std_logic_vector(to_unsigned(45,8) ,
73305	 => std_logic_vector(to_unsigned(44,8) ,
73306	 => std_logic_vector(to_unsigned(34,8) ,
73307	 => std_logic_vector(to_unsigned(33,8) ,
73308	 => std_logic_vector(to_unsigned(38,8) ,
73309	 => std_logic_vector(to_unsigned(41,8) ,
73310	 => std_logic_vector(to_unsigned(41,8) ,
73311	 => std_logic_vector(to_unsigned(45,8) ,
73312	 => std_logic_vector(to_unsigned(46,8) ,
73313	 => std_logic_vector(to_unsigned(61,8) ,
73314	 => std_logic_vector(to_unsigned(65,8) ,
73315	 => std_logic_vector(to_unsigned(60,8) ,
73316	 => std_logic_vector(to_unsigned(69,8) ,
73317	 => std_logic_vector(to_unsigned(69,8) ,
73318	 => std_logic_vector(to_unsigned(60,8) ,
73319	 => std_logic_vector(to_unsigned(37,8) ,
73320	 => std_logic_vector(to_unsigned(32,8) ,
73321	 => std_logic_vector(to_unsigned(30,8) ,
73322	 => std_logic_vector(to_unsigned(24,8) ,
73323	 => std_logic_vector(to_unsigned(29,8) ,
73324	 => std_logic_vector(to_unsigned(31,8) ,
73325	 => std_logic_vector(to_unsigned(33,8) ,
73326	 => std_logic_vector(to_unsigned(32,8) ,
73327	 => std_logic_vector(to_unsigned(29,8) ,
73328	 => std_logic_vector(to_unsigned(32,8) ,
73329	 => std_logic_vector(to_unsigned(37,8) ,
73330	 => std_logic_vector(to_unsigned(36,8) ,
73331	 => std_logic_vector(to_unsigned(41,8) ,
73332	 => std_logic_vector(to_unsigned(41,8) ,
73333	 => std_logic_vector(to_unsigned(45,8) ,
73334	 => std_logic_vector(to_unsigned(51,8) ,
73335	 => std_logic_vector(to_unsigned(86,8) ,
73336	 => std_logic_vector(to_unsigned(109,8) ,
73337	 => std_logic_vector(to_unsigned(96,8) ,
73338	 => std_logic_vector(to_unsigned(91,8) ,
73339	 => std_logic_vector(to_unsigned(91,8) ,
73340	 => std_logic_vector(to_unsigned(90,8) ,
73341	 => std_logic_vector(to_unsigned(100,8) ,
73342	 => std_logic_vector(to_unsigned(103,8) ,
73343	 => std_logic_vector(to_unsigned(97,8) ,
73344	 => std_logic_vector(to_unsigned(107,8) ,
73345	 => std_logic_vector(to_unsigned(116,8) ,
73346	 => std_logic_vector(to_unsigned(133,8) ,
73347	 => std_logic_vector(to_unsigned(131,8) ,
73348	 => std_logic_vector(to_unsigned(85,8) ,
73349	 => std_logic_vector(to_unsigned(39,8) ,
73350	 => std_logic_vector(to_unsigned(37,8) ,
73351	 => std_logic_vector(to_unsigned(42,8) ,
73352	 => std_logic_vector(to_unsigned(40,8) ,
73353	 => std_logic_vector(to_unsigned(43,8) ,
73354	 => std_logic_vector(to_unsigned(56,8) ,
73355	 => std_logic_vector(to_unsigned(57,8) ,
73356	 => std_logic_vector(to_unsigned(63,8) ,
73357	 => std_logic_vector(to_unsigned(68,8) ,
73358	 => std_logic_vector(to_unsigned(68,8) ,
73359	 => std_logic_vector(to_unsigned(59,8) ,
73360	 => std_logic_vector(to_unsigned(54,8) ,
73361	 => std_logic_vector(to_unsigned(66,8) ,
73362	 => std_logic_vector(to_unsigned(63,8) ,
73363	 => std_logic_vector(to_unsigned(68,8) ,
73364	 => std_logic_vector(to_unsigned(78,8) ,
73365	 => std_logic_vector(to_unsigned(62,8) ,
73366	 => std_logic_vector(to_unsigned(45,8) ,
73367	 => std_logic_vector(to_unsigned(45,8) ,
73368	 => std_logic_vector(to_unsigned(61,8) ,
73369	 => std_logic_vector(to_unsigned(53,8) ,
73370	 => std_logic_vector(to_unsigned(45,8) ,
73371	 => std_logic_vector(to_unsigned(53,8) ,
73372	 => std_logic_vector(to_unsigned(54,8) ,
73373	 => std_logic_vector(to_unsigned(51,8) ,
73374	 => std_logic_vector(to_unsigned(43,8) ,
73375	 => std_logic_vector(to_unsigned(35,8) ,
73376	 => std_logic_vector(to_unsigned(41,8) ,
73377	 => std_logic_vector(to_unsigned(38,8) ,
73378	 => std_logic_vector(to_unsigned(24,8) ,
73379	 => std_logic_vector(to_unsigned(35,8) ,
73380	 => std_logic_vector(to_unsigned(37,8) ,
73381	 => std_logic_vector(to_unsigned(35,8) ,
73382	 => std_logic_vector(to_unsigned(52,8) ,
73383	 => std_logic_vector(to_unsigned(82,8) ,
73384	 => std_logic_vector(to_unsigned(109,8) ,
73385	 => std_logic_vector(to_unsigned(43,8) ,
73386	 => std_logic_vector(to_unsigned(82,8) ,
73387	 => std_logic_vector(to_unsigned(134,8) ,
73388	 => std_logic_vector(to_unsigned(37,8) ,
73389	 => std_logic_vector(to_unsigned(74,8) ,
73390	 => std_logic_vector(to_unsigned(125,8) ,
73391	 => std_logic_vector(to_unsigned(58,8) ,
73392	 => std_logic_vector(to_unsigned(99,8) ,
73393	 => std_logic_vector(to_unsigned(119,8) ,
73394	 => std_logic_vector(to_unsigned(95,8) ,
73395	 => std_logic_vector(to_unsigned(100,8) ,
73396	 => std_logic_vector(to_unsigned(93,8) ,
73397	 => std_logic_vector(to_unsigned(86,8) ,
73398	 => std_logic_vector(to_unsigned(104,8) ,
73399	 => std_logic_vector(to_unsigned(121,8) ,
73400	 => std_logic_vector(to_unsigned(119,8) ,
73401	 => std_logic_vector(to_unsigned(112,8) ,
73402	 => std_logic_vector(to_unsigned(109,8) ,
73403	 => std_logic_vector(to_unsigned(105,8) ,
73404	 => std_logic_vector(to_unsigned(96,8) ,
73405	 => std_logic_vector(to_unsigned(90,8) ,
73406	 => std_logic_vector(to_unsigned(100,8) ,
73407	 => std_logic_vector(to_unsigned(96,8) ,
73408	 => std_logic_vector(to_unsigned(86,8) ,
73409	 => std_logic_vector(to_unsigned(85,8) ,
73410	 => std_logic_vector(to_unsigned(87,8) ,
73411	 => std_logic_vector(to_unsigned(88,8) ,
73412	 => std_logic_vector(to_unsigned(80,8) ,
73413	 => std_logic_vector(to_unsigned(79,8) ,
73414	 => std_logic_vector(to_unsigned(90,8) ,
73415	 => std_logic_vector(to_unsigned(92,8) ,
73416	 => std_logic_vector(to_unsigned(92,8) ,
73417	 => std_logic_vector(to_unsigned(90,8) ,
73418	 => std_logic_vector(to_unsigned(73,8) ,
73419	 => std_logic_vector(to_unsigned(67,8) ,
73420	 => std_logic_vector(to_unsigned(60,8) ,
73421	 => std_logic_vector(to_unsigned(46,8) ,
73422	 => std_logic_vector(to_unsigned(38,8) ,
73423	 => std_logic_vector(to_unsigned(47,8) ,
73424	 => std_logic_vector(to_unsigned(49,8) ,
73425	 => std_logic_vector(to_unsigned(46,8) ,
73426	 => std_logic_vector(to_unsigned(43,8) ,
73427	 => std_logic_vector(to_unsigned(44,8) ,
73428	 => std_logic_vector(to_unsigned(39,8) ,
73429	 => std_logic_vector(to_unsigned(28,8) ,
73430	 => std_logic_vector(to_unsigned(88,8) ,
73431	 => std_logic_vector(to_unsigned(115,8) ,
73432	 => std_logic_vector(to_unsigned(103,8) ,
73433	 => std_logic_vector(to_unsigned(101,8) ,
73434	 => std_logic_vector(to_unsigned(92,8) ,
73435	 => std_logic_vector(to_unsigned(87,8) ,
73436	 => std_logic_vector(to_unsigned(88,8) ,
73437	 => std_logic_vector(to_unsigned(79,8) ,
73438	 => std_logic_vector(to_unsigned(53,8) ,
73439	 => std_logic_vector(to_unsigned(18,8) ,
73440	 => std_logic_vector(to_unsigned(45,8) ,
73441	 => std_logic_vector(to_unsigned(27,8) ,
73442	 => std_logic_vector(to_unsigned(33,8) ,
73443	 => std_logic_vector(to_unsigned(32,8) ,
73444	 => std_logic_vector(to_unsigned(20,8) ,
73445	 => std_logic_vector(to_unsigned(37,8) ,
73446	 => std_logic_vector(to_unsigned(52,8) ,
73447	 => std_logic_vector(to_unsigned(8,8) ,
73448	 => std_logic_vector(to_unsigned(4,8) ,
73449	 => std_logic_vector(to_unsigned(12,8) ,
73450	 => std_logic_vector(to_unsigned(10,8) ,
73451	 => std_logic_vector(to_unsigned(17,8) ,
73452	 => std_logic_vector(to_unsigned(20,8) ,
73453	 => std_logic_vector(to_unsigned(12,8) ,
73454	 => std_logic_vector(to_unsigned(26,8) ,
73455	 => std_logic_vector(to_unsigned(17,8) ,
73456	 => std_logic_vector(to_unsigned(29,8) ,
73457	 => std_logic_vector(to_unsigned(66,8) ,
73458	 => std_logic_vector(to_unsigned(52,8) ,
73459	 => std_logic_vector(to_unsigned(17,8) ,
73460	 => std_logic_vector(to_unsigned(43,8) ,
73461	 => std_logic_vector(to_unsigned(52,8) ,
73462	 => std_logic_vector(to_unsigned(23,8) ,
73463	 => std_logic_vector(to_unsigned(29,8) ,
73464	 => std_logic_vector(to_unsigned(27,8) ,
73465	 => std_logic_vector(to_unsigned(12,8) ,
73466	 => std_logic_vector(to_unsigned(17,8) ,
73467	 => std_logic_vector(to_unsigned(46,8) ,
73468	 => std_logic_vector(to_unsigned(85,8) ,
73469	 => std_logic_vector(to_unsigned(61,8) ,
73470	 => std_logic_vector(to_unsigned(29,8) ,
73471	 => std_logic_vector(to_unsigned(25,8) ,
73472	 => std_logic_vector(to_unsigned(40,8) ,
73473	 => std_logic_vector(to_unsigned(47,8) ,
73474	 => std_logic_vector(to_unsigned(32,8) ,
73475	 => std_logic_vector(to_unsigned(22,8) ,
73476	 => std_logic_vector(to_unsigned(22,8) ,
73477	 => std_logic_vector(to_unsigned(38,8) ,
73478	 => std_logic_vector(to_unsigned(52,8) ,
73479	 => std_logic_vector(to_unsigned(49,8) ,
73480	 => std_logic_vector(to_unsigned(27,8) ,
73481	 => std_logic_vector(to_unsigned(19,8) ,
73482	 => std_logic_vector(to_unsigned(9,8) ,
73483	 => std_logic_vector(to_unsigned(8,8) ,
73484	 => std_logic_vector(to_unsigned(16,8) ,
73485	 => std_logic_vector(to_unsigned(14,8) ,
73486	 => std_logic_vector(to_unsigned(10,8) ,
73487	 => std_logic_vector(to_unsigned(10,8) ,
73488	 => std_logic_vector(to_unsigned(15,8) ,
73489	 => std_logic_vector(to_unsigned(27,8) ,
73490	 => std_logic_vector(to_unsigned(37,8) ,
73491	 => std_logic_vector(to_unsigned(22,8) ,
73492	 => std_logic_vector(to_unsigned(13,8) ,
73493	 => std_logic_vector(to_unsigned(17,8) ,
73494	 => std_logic_vector(to_unsigned(32,8) ,
73495	 => std_logic_vector(to_unsigned(50,8) ,
73496	 => std_logic_vector(to_unsigned(50,8) ,
73497	 => std_logic_vector(to_unsigned(21,8) ,
73498	 => std_logic_vector(to_unsigned(18,8) ,
73499	 => std_logic_vector(to_unsigned(32,8) ,
73500	 => std_logic_vector(to_unsigned(64,8) ,
73501	 => std_logic_vector(to_unsigned(61,8) ,
73502	 => std_logic_vector(to_unsigned(24,8) ,
73503	 => std_logic_vector(to_unsigned(19,8) ,
73504	 => std_logic_vector(to_unsigned(35,8) ,
73505	 => std_logic_vector(to_unsigned(28,8) ,
73506	 => std_logic_vector(to_unsigned(27,8) ,
73507	 => std_logic_vector(to_unsigned(27,8) ,
73508	 => std_logic_vector(to_unsigned(14,8) ,
73509	 => std_logic_vector(to_unsigned(3,8) ,
73510	 => std_logic_vector(to_unsigned(15,8) ,
73511	 => std_logic_vector(to_unsigned(24,8) ,
73512	 => std_logic_vector(to_unsigned(19,8) ,
73513	 => std_logic_vector(to_unsigned(17,8) ,
73514	 => std_logic_vector(to_unsigned(28,8) ,
73515	 => std_logic_vector(to_unsigned(40,8) ,
73516	 => std_logic_vector(to_unsigned(32,8) ,
73517	 => std_logic_vector(to_unsigned(30,8) ,
73518	 => std_logic_vector(to_unsigned(39,8) ,
73519	 => std_logic_vector(to_unsigned(37,8) ,
73520	 => std_logic_vector(to_unsigned(32,8) ,
73521	 => std_logic_vector(to_unsigned(27,8) ,
73522	 => std_logic_vector(to_unsigned(30,8) ,
73523	 => std_logic_vector(to_unsigned(25,8) ,
73524	 => std_logic_vector(to_unsigned(15,8) ,
73525	 => std_logic_vector(to_unsigned(16,8) ,
73526	 => std_logic_vector(to_unsigned(18,8) ,
73527	 => std_logic_vector(to_unsigned(30,8) ,
73528	 => std_logic_vector(to_unsigned(65,8) ,
73529	 => std_logic_vector(to_unsigned(27,8) ,
73530	 => std_logic_vector(to_unsigned(5,8) ,
73531	 => std_logic_vector(to_unsigned(10,8) ,
73532	 => std_logic_vector(to_unsigned(10,8) ,
73533	 => std_logic_vector(to_unsigned(8,8) ,
73534	 => std_logic_vector(to_unsigned(9,8) ,
73535	 => std_logic_vector(to_unsigned(11,8) ,
73536	 => std_logic_vector(to_unsigned(13,8) ,
73537	 => std_logic_vector(to_unsigned(11,8) ,
73538	 => std_logic_vector(to_unsigned(10,8) ,
73539	 => std_logic_vector(to_unsigned(12,8) ,
73540	 => std_logic_vector(to_unsigned(8,8) ,
73541	 => std_logic_vector(to_unsigned(5,8) ,
73542	 => std_logic_vector(to_unsigned(5,8) ,
73543	 => std_logic_vector(to_unsigned(5,8) ,
73544	 => std_logic_vector(to_unsigned(6,8) ,
73545	 => std_logic_vector(to_unsigned(11,8) ,
73546	 => std_logic_vector(to_unsigned(11,8) ,
73547	 => std_logic_vector(to_unsigned(18,8) ,
73548	 => std_logic_vector(to_unsigned(16,8) ,
73549	 => std_logic_vector(to_unsigned(11,8) ,
73550	 => std_logic_vector(to_unsigned(12,8) ,
73551	 => std_logic_vector(to_unsigned(11,8) ,
73552	 => std_logic_vector(to_unsigned(15,8) ,
73553	 => std_logic_vector(to_unsigned(9,8) ,
73554	 => std_logic_vector(to_unsigned(10,8) ,
73555	 => std_logic_vector(to_unsigned(11,8) ,
73556	 => std_logic_vector(to_unsigned(11,8) ,
73557	 => std_logic_vector(to_unsigned(32,8) ,
73558	 => std_logic_vector(to_unsigned(14,8) ,
73559	 => std_logic_vector(to_unsigned(0,8) ,
73560	 => std_logic_vector(to_unsigned(1,8) ,
73561	 => std_logic_vector(to_unsigned(17,8) ,
73562	 => std_logic_vector(to_unsigned(11,8) ,
73563	 => std_logic_vector(to_unsigned(20,8) ,
73564	 => std_logic_vector(to_unsigned(35,8) ,
73565	 => std_logic_vector(to_unsigned(29,8) ,
73566	 => std_logic_vector(to_unsigned(27,8) ,
73567	 => std_logic_vector(to_unsigned(28,8) ,
73568	 => std_logic_vector(to_unsigned(27,8) ,
73569	 => std_logic_vector(to_unsigned(40,8) ,
73570	 => std_logic_vector(to_unsigned(22,8) ,
73571	 => std_logic_vector(to_unsigned(5,8) ,
73572	 => std_logic_vector(to_unsigned(1,8) ,
73573	 => std_logic_vector(to_unsigned(0,8) ,
73574	 => std_logic_vector(to_unsigned(0,8) ,
73575	 => std_logic_vector(to_unsigned(0,8) ,
73576	 => std_logic_vector(to_unsigned(1,8) ,
73577	 => std_logic_vector(to_unsigned(2,8) ,
73578	 => std_logic_vector(to_unsigned(4,8) ,
73579	 => std_logic_vector(to_unsigned(1,8) ,
73580	 => std_logic_vector(to_unsigned(1,8) ,
73581	 => std_logic_vector(to_unsigned(1,8) ,
73582	 => std_logic_vector(to_unsigned(1,8) ,
73583	 => std_logic_vector(to_unsigned(0,8) ,
73584	 => std_logic_vector(to_unsigned(10,8) ,
73585	 => std_logic_vector(to_unsigned(45,8) ,
73586	 => std_logic_vector(to_unsigned(24,8) ,
73587	 => std_logic_vector(to_unsigned(24,8) ,
73588	 => std_logic_vector(to_unsigned(21,8) ,
73589	 => std_logic_vector(to_unsigned(17,8) ,
73590	 => std_logic_vector(to_unsigned(29,8) ,
73591	 => std_logic_vector(to_unsigned(33,8) ,
73592	 => std_logic_vector(to_unsigned(35,8) ,
73593	 => std_logic_vector(to_unsigned(47,8) ,
73594	 => std_logic_vector(to_unsigned(62,8) ,
73595	 => std_logic_vector(to_unsigned(79,8) ,
73596	 => std_logic_vector(to_unsigned(82,8) ,
73597	 => std_logic_vector(to_unsigned(70,8) ,
73598	 => std_logic_vector(to_unsigned(64,8) ,
73599	 => std_logic_vector(to_unsigned(69,8) ,
73600	 => std_logic_vector(to_unsigned(73,8) ,
73601	 => std_logic_vector(to_unsigned(107,8) ,
73602	 => std_logic_vector(to_unsigned(109,8) ,
73603	 => std_logic_vector(to_unsigned(114,8) ,
73604	 => std_logic_vector(to_unsigned(92,8) ,
73605	 => std_logic_vector(to_unsigned(112,8) ,
73606	 => std_logic_vector(to_unsigned(122,8) ,
73607	 => std_logic_vector(to_unsigned(111,8) ,
73608	 => std_logic_vector(to_unsigned(108,8) ,
73609	 => std_logic_vector(to_unsigned(122,8) ,
73610	 => std_logic_vector(to_unsigned(119,8) ,
73611	 => std_logic_vector(to_unsigned(118,8) ,
73612	 => std_logic_vector(to_unsigned(93,8) ,
73613	 => std_logic_vector(to_unsigned(80,8) ,
73614	 => std_logic_vector(to_unsigned(80,8) ,
73615	 => std_logic_vector(to_unsigned(82,8) ,
73616	 => std_logic_vector(to_unsigned(80,8) ,
73617	 => std_logic_vector(to_unsigned(81,8) ,
73618	 => std_logic_vector(to_unsigned(77,8) ,
73619	 => std_logic_vector(to_unsigned(74,8) ,
73620	 => std_logic_vector(to_unsigned(66,8) ,
73621	 => std_logic_vector(to_unsigned(58,8) ,
73622	 => std_logic_vector(to_unsigned(54,8) ,
73623	 => std_logic_vector(to_unsigned(46,8) ,
73624	 => std_logic_vector(to_unsigned(48,8) ,
73625	 => std_logic_vector(to_unsigned(59,8) ,
73626	 => std_logic_vector(to_unsigned(41,8) ,
73627	 => std_logic_vector(to_unsigned(41,8) ,
73628	 => std_logic_vector(to_unsigned(37,8) ,
73629	 => std_logic_vector(to_unsigned(37,8) ,
73630	 => std_logic_vector(to_unsigned(41,8) ,
73631	 => std_logic_vector(to_unsigned(51,8) ,
73632	 => std_logic_vector(to_unsigned(52,8) ,
73633	 => std_logic_vector(to_unsigned(56,8) ,
73634	 => std_logic_vector(to_unsigned(63,8) ,
73635	 => std_logic_vector(to_unsigned(70,8) ,
73636	 => std_logic_vector(to_unsigned(71,8) ,
73637	 => std_logic_vector(to_unsigned(56,8) ,
73638	 => std_logic_vector(to_unsigned(43,8) ,
73639	 => std_logic_vector(to_unsigned(55,8) ,
73640	 => std_logic_vector(to_unsigned(59,8) ,
73641	 => std_logic_vector(to_unsigned(57,8) ,
73642	 => std_logic_vector(to_unsigned(57,8) ,
73643	 => std_logic_vector(to_unsigned(45,8) ,
73644	 => std_logic_vector(to_unsigned(31,8) ,
73645	 => std_logic_vector(to_unsigned(29,8) ,
73646	 => std_logic_vector(to_unsigned(32,8) ,
73647	 => std_logic_vector(to_unsigned(35,8) ,
73648	 => std_logic_vector(to_unsigned(30,8) ,
73649	 => std_logic_vector(to_unsigned(16,8) ,
73650	 => std_logic_vector(to_unsigned(25,8) ,
73651	 => std_logic_vector(to_unsigned(46,8) ,
73652	 => std_logic_vector(to_unsigned(41,8) ,
73653	 => std_logic_vector(to_unsigned(54,8) ,
73654	 => std_logic_vector(to_unsigned(79,8) ,
73655	 => std_logic_vector(to_unsigned(104,8) ,
73656	 => std_logic_vector(to_unsigned(104,8) ,
73657	 => std_logic_vector(to_unsigned(101,8) ,
73658	 => std_logic_vector(to_unsigned(93,8) ,
73659	 => std_logic_vector(to_unsigned(81,8) ,
73660	 => std_logic_vector(to_unsigned(84,8) ,
73661	 => std_logic_vector(to_unsigned(90,8) ,
73662	 => std_logic_vector(to_unsigned(65,8) ,
73663	 => std_logic_vector(to_unsigned(67,8) ,
73664	 => std_logic_vector(to_unsigned(108,8) ,
73665	 => std_logic_vector(to_unsigned(144,8) ,
73666	 => std_logic_vector(to_unsigned(138,8) ,
73667	 => std_logic_vector(to_unsigned(142,8) ,
73668	 => std_logic_vector(to_unsigned(95,8) ,
73669	 => std_logic_vector(to_unsigned(32,8) ,
73670	 => std_logic_vector(to_unsigned(29,8) ,
73671	 => std_logic_vector(to_unsigned(38,8) ,
73672	 => std_logic_vector(to_unsigned(39,8) ,
73673	 => std_logic_vector(to_unsigned(41,8) ,
73674	 => std_logic_vector(to_unsigned(44,8) ,
73675	 => std_logic_vector(to_unsigned(43,8) ,
73676	 => std_logic_vector(to_unsigned(41,8) ,
73677	 => std_logic_vector(to_unsigned(51,8) ,
73678	 => std_logic_vector(to_unsigned(57,8) ,
73679	 => std_logic_vector(to_unsigned(81,8) ,
73680	 => std_logic_vector(to_unsigned(96,8) ,
73681	 => std_logic_vector(to_unsigned(91,8) ,
73682	 => std_logic_vector(to_unsigned(71,8) ,
73683	 => std_logic_vector(to_unsigned(76,8) ,
73684	 => std_logic_vector(to_unsigned(62,8) ,
73685	 => std_logic_vector(to_unsigned(51,8) ,
73686	 => std_logic_vector(to_unsigned(41,8) ,
73687	 => std_logic_vector(to_unsigned(45,8) ,
73688	 => std_logic_vector(to_unsigned(46,8) ,
73689	 => std_logic_vector(to_unsigned(44,8) ,
73690	 => std_logic_vector(to_unsigned(42,8) ,
73691	 => std_logic_vector(to_unsigned(45,8) ,
73692	 => std_logic_vector(to_unsigned(45,8) ,
73693	 => std_logic_vector(to_unsigned(45,8) ,
73694	 => std_logic_vector(to_unsigned(47,8) ,
73695	 => std_logic_vector(to_unsigned(49,8) ,
73696	 => std_logic_vector(to_unsigned(45,8) ,
73697	 => std_logic_vector(to_unsigned(40,8) ,
73698	 => std_logic_vector(to_unsigned(43,8) ,
73699	 => std_logic_vector(to_unsigned(41,8) ,
73700	 => std_logic_vector(to_unsigned(32,8) ,
73701	 => std_logic_vector(to_unsigned(51,8) ,
73702	 => std_logic_vector(to_unsigned(84,8) ,
73703	 => std_logic_vector(to_unsigned(86,8) ,
73704	 => std_logic_vector(to_unsigned(107,8) ,
73705	 => std_logic_vector(to_unsigned(88,8) ,
73706	 => std_logic_vector(to_unsigned(111,8) ,
73707	 => std_logic_vector(to_unsigned(133,8) ,
73708	 => std_logic_vector(to_unsigned(52,8) ,
73709	 => std_logic_vector(to_unsigned(78,8) ,
73710	 => std_logic_vector(to_unsigned(111,8) ,
73711	 => std_logic_vector(to_unsigned(19,8) ,
73712	 => std_logic_vector(to_unsigned(58,8) ,
73713	 => std_logic_vector(to_unsigned(127,8) ,
73714	 => std_logic_vector(to_unsigned(51,8) ,
73715	 => std_logic_vector(to_unsigned(58,8) ,
73716	 => std_logic_vector(to_unsigned(81,8) ,
73717	 => std_logic_vector(to_unsigned(71,8) ,
73718	 => std_logic_vector(to_unsigned(101,8) ,
73719	 => std_logic_vector(to_unsigned(107,8) ,
73720	 => std_logic_vector(to_unsigned(108,8) ,
73721	 => std_logic_vector(to_unsigned(105,8) ,
73722	 => std_logic_vector(to_unsigned(105,8) ,
73723	 => std_logic_vector(to_unsigned(108,8) ,
73724	 => std_logic_vector(to_unsigned(101,8) ,
73725	 => std_logic_vector(to_unsigned(100,8) ,
73726	 => std_logic_vector(to_unsigned(105,8) ,
73727	 => std_logic_vector(to_unsigned(97,8) ,
73728	 => std_logic_vector(to_unsigned(84,8) ,
73729	 => std_logic_vector(to_unsigned(72,8) ,
73730	 => std_logic_vector(to_unsigned(81,8) ,
73731	 => std_logic_vector(to_unsigned(72,8) ,
73732	 => std_logic_vector(to_unsigned(58,8) ,
73733	 => std_logic_vector(to_unsigned(56,8) ,
73734	 => std_logic_vector(to_unsigned(65,8) ,
73735	 => std_logic_vector(to_unsigned(56,8) ,
73736	 => std_logic_vector(to_unsigned(59,8) ,
73737	 => std_logic_vector(to_unsigned(87,8) ,
73738	 => std_logic_vector(to_unsigned(87,8) ,
73739	 => std_logic_vector(to_unsigned(85,8) ,
73740	 => std_logic_vector(to_unsigned(87,8) ,
73741	 => std_logic_vector(to_unsigned(74,8) ,
73742	 => std_logic_vector(to_unsigned(68,8) ,
73743	 => std_logic_vector(to_unsigned(63,8) ,
73744	 => std_logic_vector(to_unsigned(52,8) ,
73745	 => std_logic_vector(to_unsigned(46,8) ,
73746	 => std_logic_vector(to_unsigned(45,8) ,
73747	 => std_logic_vector(to_unsigned(41,8) ,
73748	 => std_logic_vector(to_unsigned(37,8) ,
73749	 => std_logic_vector(to_unsigned(40,8) ,
73750	 => std_logic_vector(to_unsigned(95,8) ,
73751	 => std_logic_vector(to_unsigned(107,8) ,
73752	 => std_logic_vector(to_unsigned(101,8) ,
73753	 => std_logic_vector(to_unsigned(103,8) ,
73754	 => std_logic_vector(to_unsigned(100,8) ,
73755	 => std_logic_vector(to_unsigned(93,8) ,
73756	 => std_logic_vector(to_unsigned(72,8) ,
73757	 => std_logic_vector(to_unsigned(69,8) ,
73758	 => std_logic_vector(to_unsigned(53,8) ,
73759	 => std_logic_vector(to_unsigned(20,8) ,
73760	 => std_logic_vector(to_unsigned(50,8) ,
73761	 => std_logic_vector(to_unsigned(53,8) ,
73762	 => std_logic_vector(to_unsigned(24,8) ,
73763	 => std_logic_vector(to_unsigned(23,8) ,
73764	 => std_logic_vector(to_unsigned(41,8) ,
73765	 => std_logic_vector(to_unsigned(56,8) ,
73766	 => std_logic_vector(to_unsigned(51,8) ,
73767	 => std_logic_vector(to_unsigned(6,8) ,
73768	 => std_logic_vector(to_unsigned(4,8) ,
73769	 => std_logic_vector(to_unsigned(11,8) ,
73770	 => std_logic_vector(to_unsigned(12,8) ,
73771	 => std_logic_vector(to_unsigned(13,8) ,
73772	 => std_logic_vector(to_unsigned(12,8) ,
73773	 => std_logic_vector(to_unsigned(24,8) ,
73774	 => std_logic_vector(to_unsigned(19,8) ,
73775	 => std_logic_vector(to_unsigned(20,8) ,
73776	 => std_logic_vector(to_unsigned(69,8) ,
73777	 => std_logic_vector(to_unsigned(63,8) ,
73778	 => std_logic_vector(to_unsigned(31,8) ,
73779	 => std_logic_vector(to_unsigned(41,8) ,
73780	 => std_logic_vector(to_unsigned(67,8) ,
73781	 => std_logic_vector(to_unsigned(27,8) ,
73782	 => std_logic_vector(to_unsigned(25,8) ,
73783	 => std_logic_vector(to_unsigned(37,8) ,
73784	 => std_logic_vector(to_unsigned(45,8) ,
73785	 => std_logic_vector(to_unsigned(20,8) ,
73786	 => std_logic_vector(to_unsigned(18,8) ,
73787	 => std_logic_vector(to_unsigned(42,8) ,
73788	 => std_logic_vector(to_unsigned(76,8) ,
73789	 => std_logic_vector(to_unsigned(64,8) ,
73790	 => std_logic_vector(to_unsigned(27,8) ,
73791	 => std_logic_vector(to_unsigned(24,8) ,
73792	 => std_logic_vector(to_unsigned(46,8) ,
73793	 => std_logic_vector(to_unsigned(68,8) ,
73794	 => std_logic_vector(to_unsigned(45,8) ,
73795	 => std_logic_vector(to_unsigned(21,8) ,
73796	 => std_logic_vector(to_unsigned(24,8) ,
73797	 => std_logic_vector(to_unsigned(27,8) ,
73798	 => std_logic_vector(to_unsigned(37,8) ,
73799	 => std_logic_vector(to_unsigned(35,8) ,
73800	 => std_logic_vector(to_unsigned(26,8) ,
73801	 => std_logic_vector(to_unsigned(15,8) ,
73802	 => std_logic_vector(to_unsigned(11,8) ,
73803	 => std_logic_vector(to_unsigned(9,8) ,
73804	 => std_logic_vector(to_unsigned(9,8) ,
73805	 => std_logic_vector(to_unsigned(13,8) ,
73806	 => std_logic_vector(to_unsigned(9,8) ,
73807	 => std_logic_vector(to_unsigned(9,8) ,
73808	 => std_logic_vector(to_unsigned(13,8) ,
73809	 => std_logic_vector(to_unsigned(41,8) ,
73810	 => std_logic_vector(to_unsigned(68,8) ,
73811	 => std_logic_vector(to_unsigned(39,8) ,
73812	 => std_logic_vector(to_unsigned(14,8) ,
73813	 => std_logic_vector(to_unsigned(16,8) ,
73814	 => std_logic_vector(to_unsigned(17,8) ,
73815	 => std_logic_vector(to_unsigned(20,8) ,
73816	 => std_logic_vector(to_unsigned(25,8) ,
73817	 => std_logic_vector(to_unsigned(18,8) ,
73818	 => std_logic_vector(to_unsigned(19,8) ,
73819	 => std_logic_vector(to_unsigned(20,8) ,
73820	 => std_logic_vector(to_unsigned(37,8) ,
73821	 => std_logic_vector(to_unsigned(45,8) ,
73822	 => std_logic_vector(to_unsigned(23,8) ,
73823	 => std_logic_vector(to_unsigned(23,8) ,
73824	 => std_logic_vector(to_unsigned(30,8) ,
73825	 => std_logic_vector(to_unsigned(28,8) ,
73826	 => std_logic_vector(to_unsigned(27,8) ,
73827	 => std_logic_vector(to_unsigned(23,8) ,
73828	 => std_logic_vector(to_unsigned(14,8) ,
73829	 => std_logic_vector(to_unsigned(3,8) ,
73830	 => std_logic_vector(to_unsigned(13,8) ,
73831	 => std_logic_vector(to_unsigned(12,8) ,
73832	 => std_logic_vector(to_unsigned(7,8) ,
73833	 => std_logic_vector(to_unsigned(8,8) ,
73834	 => std_logic_vector(to_unsigned(20,8) ,
73835	 => std_logic_vector(to_unsigned(34,8) ,
73836	 => std_logic_vector(to_unsigned(15,8) ,
73837	 => std_logic_vector(to_unsigned(23,8) ,
73838	 => std_logic_vector(to_unsigned(37,8) ,
73839	 => std_logic_vector(to_unsigned(31,8) ,
73840	 => std_logic_vector(to_unsigned(23,8) ,
73841	 => std_logic_vector(to_unsigned(17,8) ,
73842	 => std_logic_vector(to_unsigned(22,8) ,
73843	 => std_logic_vector(to_unsigned(15,8) ,
73844	 => std_logic_vector(to_unsigned(16,8) ,
73845	 => std_logic_vector(to_unsigned(21,8) ,
73846	 => std_logic_vector(to_unsigned(13,8) ,
73847	 => std_logic_vector(to_unsigned(14,8) ,
73848	 => std_logic_vector(to_unsigned(44,8) ,
73849	 => std_logic_vector(to_unsigned(14,8) ,
73850	 => std_logic_vector(to_unsigned(8,8) ,
73851	 => std_logic_vector(to_unsigned(10,8) ,
73852	 => std_logic_vector(to_unsigned(6,8) ,
73853	 => std_logic_vector(to_unsigned(11,8) ,
73854	 => std_logic_vector(to_unsigned(20,8) ,
73855	 => std_logic_vector(to_unsigned(19,8) ,
73856	 => std_logic_vector(to_unsigned(19,8) ,
73857	 => std_logic_vector(to_unsigned(13,8) ,
73858	 => std_logic_vector(to_unsigned(7,8) ,
73859	 => std_logic_vector(to_unsigned(9,8) ,
73860	 => std_logic_vector(to_unsigned(8,8) ,
73861	 => std_logic_vector(to_unsigned(8,8) ,
73862	 => std_logic_vector(to_unsigned(14,8) ,
73863	 => std_logic_vector(to_unsigned(10,8) ,
73864	 => std_logic_vector(to_unsigned(10,8) ,
73865	 => std_logic_vector(to_unsigned(8,8) ,
73866	 => std_logic_vector(to_unsigned(8,8) ,
73867	 => std_logic_vector(to_unsigned(17,8) ,
73868	 => std_logic_vector(to_unsigned(18,8) ,
73869	 => std_logic_vector(to_unsigned(6,8) ,
73870	 => std_logic_vector(to_unsigned(5,8) ,
73871	 => std_logic_vector(to_unsigned(16,8) ,
73872	 => std_logic_vector(to_unsigned(32,8) ,
73873	 => std_logic_vector(to_unsigned(12,8) ,
73874	 => std_logic_vector(to_unsigned(6,8) ,
73875	 => std_logic_vector(to_unsigned(10,8) ,
73876	 => std_logic_vector(to_unsigned(13,8) ,
73877	 => std_logic_vector(to_unsigned(29,8) ,
73878	 => std_logic_vector(to_unsigned(23,8) ,
73879	 => std_logic_vector(to_unsigned(2,8) ,
73880	 => std_logic_vector(to_unsigned(0,8) ,
73881	 => std_logic_vector(to_unsigned(3,8) ,
73882	 => std_logic_vector(to_unsigned(8,8) ,
73883	 => std_logic_vector(to_unsigned(29,8) ,
73884	 => std_logic_vector(to_unsigned(38,8) ,
73885	 => std_logic_vector(to_unsigned(33,8) ,
73886	 => std_logic_vector(to_unsigned(35,8) ,
73887	 => std_logic_vector(to_unsigned(33,8) ,
73888	 => std_logic_vector(to_unsigned(37,8) ,
73889	 => std_logic_vector(to_unsigned(39,8) ,
73890	 => std_logic_vector(to_unsigned(28,8) ,
73891	 => std_logic_vector(to_unsigned(25,8) ,
73892	 => std_logic_vector(to_unsigned(7,8) ,
73893	 => std_logic_vector(to_unsigned(0,8) ,
73894	 => std_logic_vector(to_unsigned(0,8) ,
73895	 => std_logic_vector(to_unsigned(0,8) ,
73896	 => std_logic_vector(to_unsigned(0,8) ,
73897	 => std_logic_vector(to_unsigned(0,8) ,
73898	 => std_logic_vector(to_unsigned(1,8) ,
73899	 => std_logic_vector(to_unsigned(0,8) ,
73900	 => std_logic_vector(to_unsigned(0,8) ,
73901	 => std_logic_vector(to_unsigned(0,8) ,
73902	 => std_logic_vector(to_unsigned(0,8) ,
73903	 => std_logic_vector(to_unsigned(1,8) ,
73904	 => std_logic_vector(to_unsigned(30,8) ,
73905	 => std_logic_vector(to_unsigned(47,8) ,
73906	 => std_logic_vector(to_unsigned(22,8) ,
73907	 => std_logic_vector(to_unsigned(36,8) ,
73908	 => std_logic_vector(to_unsigned(22,8) ,
73909	 => std_logic_vector(to_unsigned(10,8) ,
73910	 => std_logic_vector(to_unsigned(8,8) ,
73911	 => std_logic_vector(to_unsigned(11,8) ,
73912	 => std_logic_vector(to_unsigned(13,8) ,
73913	 => std_logic_vector(to_unsigned(12,8) ,
73914	 => std_logic_vector(to_unsigned(26,8) ,
73915	 => std_logic_vector(to_unsigned(87,8) ,
73916	 => std_logic_vector(to_unsigned(84,8) ,
73917	 => std_logic_vector(to_unsigned(79,8) ,
73918	 => std_logic_vector(to_unsigned(84,8) ,
73919	 => std_logic_vector(to_unsigned(84,8) ,
73920	 => std_logic_vector(to_unsigned(99,8) ,
73921	 => std_logic_vector(to_unsigned(104,8) ,
73922	 => std_logic_vector(to_unsigned(104,8) ,
73923	 => std_logic_vector(to_unsigned(112,8) ,
73924	 => std_logic_vector(to_unsigned(99,8) ,
73925	 => std_logic_vector(to_unsigned(121,8) ,
73926	 => std_logic_vector(to_unsigned(138,8) ,
73927	 => std_logic_vector(to_unsigned(133,8) ,
73928	 => std_logic_vector(to_unsigned(125,8) ,
73929	 => std_logic_vector(to_unsigned(128,8) ,
73930	 => std_logic_vector(to_unsigned(128,8) ,
73931	 => std_logic_vector(to_unsigned(121,8) ,
73932	 => std_logic_vector(to_unsigned(96,8) ,
73933	 => std_logic_vector(to_unsigned(85,8) ,
73934	 => std_logic_vector(to_unsigned(79,8) ,
73935	 => std_logic_vector(to_unsigned(77,8) ,
73936	 => std_logic_vector(to_unsigned(79,8) ,
73937	 => std_logic_vector(to_unsigned(86,8) ,
73938	 => std_logic_vector(to_unsigned(79,8) ,
73939	 => std_logic_vector(to_unsigned(71,8) ,
73940	 => std_logic_vector(to_unsigned(62,8) ,
73941	 => std_logic_vector(to_unsigned(58,8) ,
73942	 => std_logic_vector(to_unsigned(56,8) ,
73943	 => std_logic_vector(to_unsigned(41,8) ,
73944	 => std_logic_vector(to_unsigned(64,8) ,
73945	 => std_logic_vector(to_unsigned(55,8) ,
73946	 => std_logic_vector(to_unsigned(33,8) ,
73947	 => std_logic_vector(to_unsigned(41,8) ,
73948	 => std_logic_vector(to_unsigned(37,8) ,
73949	 => std_logic_vector(to_unsigned(35,8) ,
73950	 => std_logic_vector(to_unsigned(42,8) ,
73951	 => std_logic_vector(to_unsigned(56,8) ,
73952	 => std_logic_vector(to_unsigned(55,8) ,
73953	 => std_logic_vector(to_unsigned(59,8) ,
73954	 => std_logic_vector(to_unsigned(73,8) ,
73955	 => std_logic_vector(to_unsigned(72,8) ,
73956	 => std_logic_vector(to_unsigned(48,8) ,
73957	 => std_logic_vector(to_unsigned(31,8) ,
73958	 => std_logic_vector(to_unsigned(36,8) ,
73959	 => std_logic_vector(to_unsigned(58,8) ,
73960	 => std_logic_vector(to_unsigned(51,8) ,
73961	 => std_logic_vector(to_unsigned(41,8) ,
73962	 => std_logic_vector(to_unsigned(51,8) ,
73963	 => std_logic_vector(to_unsigned(66,8) ,
73964	 => std_logic_vector(to_unsigned(52,8) ,
73965	 => std_logic_vector(to_unsigned(43,8) ,
73966	 => std_logic_vector(to_unsigned(43,8) ,
73967	 => std_logic_vector(to_unsigned(56,8) ,
73968	 => std_logic_vector(to_unsigned(25,8) ,
73969	 => std_logic_vector(to_unsigned(16,8) ,
73970	 => std_logic_vector(to_unsigned(32,8) ,
73971	 => std_logic_vector(to_unsigned(52,8) ,
73972	 => std_logic_vector(to_unsigned(60,8) ,
73973	 => std_logic_vector(to_unsigned(79,8) ,
73974	 => std_logic_vector(to_unsigned(104,8) ,
73975	 => std_logic_vector(to_unsigned(100,8) ,
73976	 => std_logic_vector(to_unsigned(95,8) ,
73977	 => std_logic_vector(to_unsigned(107,8) ,
73978	 => std_logic_vector(to_unsigned(104,8) ,
73979	 => std_logic_vector(to_unsigned(82,8) ,
73980	 => std_logic_vector(to_unsigned(90,8) ,
73981	 => std_logic_vector(to_unsigned(100,8) ,
73982	 => std_logic_vector(to_unsigned(47,8) ,
73983	 => std_logic_vector(to_unsigned(58,8) ,
73984	 => std_logic_vector(to_unsigned(101,8) ,
73985	 => std_logic_vector(to_unsigned(139,8) ,
73986	 => std_logic_vector(to_unsigned(142,8) ,
73987	 => std_logic_vector(to_unsigned(100,8) ,
73988	 => std_logic_vector(to_unsigned(46,8) ,
73989	 => std_logic_vector(to_unsigned(27,8) ,
73990	 => std_logic_vector(to_unsigned(25,8) ,
73991	 => std_logic_vector(to_unsigned(26,8) ,
73992	 => std_logic_vector(to_unsigned(35,8) ,
73993	 => std_logic_vector(to_unsigned(37,8) ,
73994	 => std_logic_vector(to_unsigned(37,8) ,
73995	 => std_logic_vector(to_unsigned(30,8) ,
73996	 => std_logic_vector(to_unsigned(32,8) ,
73997	 => std_logic_vector(to_unsigned(35,8) ,
73998	 => std_logic_vector(to_unsigned(35,8) ,
73999	 => std_logic_vector(to_unsigned(73,8) ,
74000	 => std_logic_vector(to_unsigned(114,8) ,
74001	 => std_logic_vector(to_unsigned(125,8) ,
74002	 => std_logic_vector(to_unsigned(109,8) ,
74003	 => std_logic_vector(to_unsigned(118,8) ,
74004	 => std_logic_vector(to_unsigned(87,8) ,
74005	 => std_logic_vector(to_unsigned(121,8) ,
74006	 => std_logic_vector(to_unsigned(88,8) ,
74007	 => std_logic_vector(to_unsigned(85,8) ,
74008	 => std_logic_vector(to_unsigned(66,8) ,
74009	 => std_logic_vector(to_unsigned(56,8) ,
74010	 => std_logic_vector(to_unsigned(50,8) ,
74011	 => std_logic_vector(to_unsigned(42,8) ,
74012	 => std_logic_vector(to_unsigned(41,8) ,
74013	 => std_logic_vector(to_unsigned(42,8) ,
74014	 => std_logic_vector(to_unsigned(38,8) ,
74015	 => std_logic_vector(to_unsigned(37,8) ,
74016	 => std_logic_vector(to_unsigned(35,8) ,
74017	 => std_logic_vector(to_unsigned(39,8) ,
74018	 => std_logic_vector(to_unsigned(54,8) ,
74019	 => std_logic_vector(to_unsigned(55,8) ,
74020	 => std_logic_vector(to_unsigned(72,8) ,
74021	 => std_logic_vector(to_unsigned(90,8) ,
74022	 => std_logic_vector(to_unsigned(73,8) ,
74023	 => std_logic_vector(to_unsigned(63,8) ,
74024	 => std_logic_vector(to_unsigned(96,8) ,
74025	 => std_logic_vector(to_unsigned(111,8) ,
74026	 => std_logic_vector(to_unsigned(121,8) ,
74027	 => std_logic_vector(to_unsigned(131,8) ,
74028	 => std_logic_vector(to_unsigned(124,8) ,
74029	 => std_logic_vector(to_unsigned(141,8) ,
74030	 => std_logic_vector(to_unsigned(125,8) ,
74031	 => std_logic_vector(to_unsigned(61,8) ,
74032	 => std_logic_vector(to_unsigned(84,8) ,
74033	 => std_logic_vector(to_unsigned(122,8) ,
74034	 => std_logic_vector(to_unsigned(51,8) ,
74035	 => std_logic_vector(to_unsigned(35,8) ,
74036	 => std_logic_vector(to_unsigned(65,8) ,
74037	 => std_logic_vector(to_unsigned(69,8) ,
74038	 => std_logic_vector(to_unsigned(104,8) ,
74039	 => std_logic_vector(to_unsigned(108,8) ,
74040	 => std_logic_vector(to_unsigned(109,8) ,
74041	 => std_logic_vector(to_unsigned(105,8) ,
74042	 => std_logic_vector(to_unsigned(104,8) ,
74043	 => std_logic_vector(to_unsigned(101,8) ,
74044	 => std_logic_vector(to_unsigned(101,8) ,
74045	 => std_logic_vector(to_unsigned(104,8) ,
74046	 => std_logic_vector(to_unsigned(107,8) ,
74047	 => std_logic_vector(to_unsigned(107,8) ,
74048	 => std_logic_vector(to_unsigned(66,8) ,
74049	 => std_logic_vector(to_unsigned(28,8) ,
74050	 => std_logic_vector(to_unsigned(47,8) ,
74051	 => std_logic_vector(to_unsigned(51,8) ,
74052	 => std_logic_vector(to_unsigned(52,8) ,
74053	 => std_logic_vector(to_unsigned(54,8) ,
74054	 => std_logic_vector(to_unsigned(62,8) ,
74055	 => std_logic_vector(to_unsigned(53,8) ,
74056	 => std_logic_vector(to_unsigned(46,8) ,
74057	 => std_logic_vector(to_unsigned(76,8) ,
74058	 => std_logic_vector(to_unsigned(84,8) ,
74059	 => std_logic_vector(to_unsigned(77,8) ,
74060	 => std_logic_vector(to_unsigned(79,8) ,
74061	 => std_logic_vector(to_unsigned(85,8) ,
74062	 => std_logic_vector(to_unsigned(86,8) ,
74063	 => std_logic_vector(to_unsigned(80,8) ,
74064	 => std_logic_vector(to_unsigned(79,8) ,
74065	 => std_logic_vector(to_unsigned(78,8) ,
74066	 => std_logic_vector(to_unsigned(73,8) ,
74067	 => std_logic_vector(to_unsigned(63,8) ,
74068	 => std_logic_vector(to_unsigned(48,8) ,
74069	 => std_logic_vector(to_unsigned(40,8) ,
74070	 => std_logic_vector(to_unsigned(91,8) ,
74071	 => std_logic_vector(to_unsigned(100,8) ,
74072	 => std_logic_vector(to_unsigned(95,8) ,
74073	 => std_logic_vector(to_unsigned(91,8) ,
74074	 => std_logic_vector(to_unsigned(92,8) ,
74075	 => std_logic_vector(to_unsigned(88,8) ,
74076	 => std_logic_vector(to_unsigned(73,8) ,
74077	 => std_logic_vector(to_unsigned(71,8) ,
74078	 => std_logic_vector(to_unsigned(70,8) ,
74079	 => std_logic_vector(to_unsigned(67,8) ,
74080	 => std_logic_vector(to_unsigned(63,8) ,
74081	 => std_logic_vector(to_unsigned(37,8) ,
74082	 => std_logic_vector(to_unsigned(25,8) ,
74083	 => std_logic_vector(to_unsigned(31,8) ,
74084	 => std_logic_vector(to_unsigned(72,8) ,
74085	 => std_logic_vector(to_unsigned(67,8) ,
74086	 => std_logic_vector(to_unsigned(29,8) ,
74087	 => std_logic_vector(to_unsigned(5,8) ,
74088	 => std_logic_vector(to_unsigned(4,8) ,
74089	 => std_logic_vector(to_unsigned(10,8) ,
74090	 => std_logic_vector(to_unsigned(13,8) ,
74091	 => std_logic_vector(to_unsigned(14,8) ,
74092	 => std_logic_vector(to_unsigned(23,8) ,
74093	 => std_logic_vector(to_unsigned(21,8) ,
74094	 => std_logic_vector(to_unsigned(17,8) ,
74095	 => std_logic_vector(to_unsigned(59,8) ,
74096	 => std_logic_vector(to_unsigned(74,8) ,
74097	 => std_logic_vector(to_unsigned(49,8) ,
74098	 => std_logic_vector(to_unsigned(12,8) ,
74099	 => std_logic_vector(to_unsigned(14,8) ,
74100	 => std_logic_vector(to_unsigned(18,8) ,
74101	 => std_logic_vector(to_unsigned(16,8) ,
74102	 => std_logic_vector(to_unsigned(32,8) ,
74103	 => std_logic_vector(to_unsigned(33,8) ,
74104	 => std_logic_vector(to_unsigned(37,8) ,
74105	 => std_logic_vector(to_unsigned(19,8) ,
74106	 => std_logic_vector(to_unsigned(20,8) ,
74107	 => std_logic_vector(to_unsigned(32,8) ,
74108	 => std_logic_vector(to_unsigned(28,8) ,
74109	 => std_logic_vector(to_unsigned(30,8) ,
74110	 => std_logic_vector(to_unsigned(24,8) ,
74111	 => std_logic_vector(to_unsigned(27,8) ,
74112	 => std_logic_vector(to_unsigned(38,8) ,
74113	 => std_logic_vector(to_unsigned(51,8) ,
74114	 => std_logic_vector(to_unsigned(43,8) ,
74115	 => std_logic_vector(to_unsigned(23,8) ,
74116	 => std_logic_vector(to_unsigned(24,8) ,
74117	 => std_logic_vector(to_unsigned(25,8) ,
74118	 => std_logic_vector(to_unsigned(30,8) ,
74119	 => std_logic_vector(to_unsigned(32,8) ,
74120	 => std_logic_vector(to_unsigned(27,8) ,
74121	 => std_logic_vector(to_unsigned(17,8) ,
74122	 => std_logic_vector(to_unsigned(11,8) ,
74123	 => std_logic_vector(to_unsigned(7,8) ,
74124	 => std_logic_vector(to_unsigned(9,8) ,
74125	 => std_logic_vector(to_unsigned(14,8) ,
74126	 => std_logic_vector(to_unsigned(10,8) ,
74127	 => std_logic_vector(to_unsigned(8,8) ,
74128	 => std_logic_vector(to_unsigned(14,8) ,
74129	 => std_logic_vector(to_unsigned(37,8) ,
74130	 => std_logic_vector(to_unsigned(72,8) ,
74131	 => std_logic_vector(to_unsigned(54,8) ,
74132	 => std_logic_vector(to_unsigned(16,8) ,
74133	 => std_logic_vector(to_unsigned(17,8) ,
74134	 => std_logic_vector(to_unsigned(9,8) ,
74135	 => std_logic_vector(to_unsigned(5,8) ,
74136	 => std_logic_vector(to_unsigned(8,8) ,
74137	 => std_logic_vector(to_unsigned(16,8) ,
74138	 => std_logic_vector(to_unsigned(19,8) ,
74139	 => std_logic_vector(to_unsigned(18,8) ,
74140	 => std_logic_vector(to_unsigned(29,8) ,
74141	 => std_logic_vector(to_unsigned(30,8) ,
74142	 => std_logic_vector(to_unsigned(18,8) ,
74143	 => std_logic_vector(to_unsigned(24,8) ,
74144	 => std_logic_vector(to_unsigned(29,8) ,
74145	 => std_logic_vector(to_unsigned(26,8) ,
74146	 => std_logic_vector(to_unsigned(34,8) ,
74147	 => std_logic_vector(to_unsigned(30,8) ,
74148	 => std_logic_vector(to_unsigned(9,8) ,
74149	 => std_logic_vector(to_unsigned(2,8) ,
74150	 => std_logic_vector(to_unsigned(14,8) ,
74151	 => std_logic_vector(to_unsigned(18,8) ,
74152	 => std_logic_vector(to_unsigned(11,8) ,
74153	 => std_logic_vector(to_unsigned(16,8) ,
74154	 => std_logic_vector(to_unsigned(31,8) ,
74155	 => std_logic_vector(to_unsigned(30,8) ,
74156	 => std_logic_vector(to_unsigned(7,8) ,
74157	 => std_logic_vector(to_unsigned(10,8) ,
74158	 => std_logic_vector(to_unsigned(37,8) ,
74159	 => std_logic_vector(to_unsigned(29,8) ,
74160	 => std_logic_vector(to_unsigned(9,8) ,
74161	 => std_logic_vector(to_unsigned(7,8) ,
74162	 => std_logic_vector(to_unsigned(25,8) ,
74163	 => std_logic_vector(to_unsigned(20,8) ,
74164	 => std_logic_vector(to_unsigned(25,8) ,
74165	 => std_logic_vector(to_unsigned(23,8) ,
74166	 => std_logic_vector(to_unsigned(9,8) ,
74167	 => std_logic_vector(to_unsigned(38,8) ,
74168	 => std_logic_vector(to_unsigned(50,8) ,
74169	 => std_logic_vector(to_unsigned(9,8) ,
74170	 => std_logic_vector(to_unsigned(12,8) ,
74171	 => std_logic_vector(to_unsigned(12,8) ,
74172	 => std_logic_vector(to_unsigned(8,8) ,
74173	 => std_logic_vector(to_unsigned(15,8) ,
74174	 => std_logic_vector(to_unsigned(26,8) ,
74175	 => std_logic_vector(to_unsigned(23,8) ,
74176	 => std_logic_vector(to_unsigned(24,8) ,
74177	 => std_logic_vector(to_unsigned(17,8) ,
74178	 => std_logic_vector(to_unsigned(7,8) ,
74179	 => std_logic_vector(to_unsigned(11,8) ,
74180	 => std_logic_vector(to_unsigned(13,8) ,
74181	 => std_logic_vector(to_unsigned(11,8) ,
74182	 => std_logic_vector(to_unsigned(9,8) ,
74183	 => std_logic_vector(to_unsigned(10,8) ,
74184	 => std_logic_vector(to_unsigned(12,8) ,
74185	 => std_logic_vector(to_unsigned(12,8) ,
74186	 => std_logic_vector(to_unsigned(12,8) ,
74187	 => std_logic_vector(to_unsigned(15,8) ,
74188	 => std_logic_vector(to_unsigned(16,8) ,
74189	 => std_logic_vector(to_unsigned(22,8) ,
74190	 => std_logic_vector(to_unsigned(15,8) ,
74191	 => std_logic_vector(to_unsigned(15,8) ,
74192	 => std_logic_vector(to_unsigned(20,8) ,
74193	 => std_logic_vector(to_unsigned(12,8) ,
74194	 => std_logic_vector(to_unsigned(20,8) ,
74195	 => std_logic_vector(to_unsigned(24,8) ,
74196	 => std_logic_vector(to_unsigned(25,8) ,
74197	 => std_logic_vector(to_unsigned(23,8) ,
74198	 => std_logic_vector(to_unsigned(29,8) ,
74199	 => std_logic_vector(to_unsigned(7,8) ,
74200	 => std_logic_vector(to_unsigned(0,8) ,
74201	 => std_logic_vector(to_unsigned(1,8) ,
74202	 => std_logic_vector(to_unsigned(5,8) ,
74203	 => std_logic_vector(to_unsigned(29,8) ,
74204	 => std_logic_vector(to_unsigned(32,8) ,
74205	 => std_logic_vector(to_unsigned(29,8) ,
74206	 => std_logic_vector(to_unsigned(23,8) ,
74207	 => std_logic_vector(to_unsigned(27,8) ,
74208	 => std_logic_vector(to_unsigned(38,8) ,
74209	 => std_logic_vector(to_unsigned(38,8) ,
74210	 => std_logic_vector(to_unsigned(19,8) ,
74211	 => std_logic_vector(to_unsigned(19,8) ,
74212	 => std_logic_vector(to_unsigned(23,8) ,
74213	 => std_logic_vector(to_unsigned(6,8) ,
74214	 => std_logic_vector(to_unsigned(0,8) ,
74215	 => std_logic_vector(to_unsigned(0,8) ,
74216	 => std_logic_vector(to_unsigned(0,8) ,
74217	 => std_logic_vector(to_unsigned(0,8) ,
74218	 => std_logic_vector(to_unsigned(0,8) ,
74219	 => std_logic_vector(to_unsigned(0,8) ,
74220	 => std_logic_vector(to_unsigned(0,8) ,
74221	 => std_logic_vector(to_unsigned(1,8) ,
74222	 => std_logic_vector(to_unsigned(8,8) ,
74223	 => std_logic_vector(to_unsigned(23,8) ,
74224	 => std_logic_vector(to_unsigned(45,8) ,
74225	 => std_logic_vector(to_unsigned(37,8) ,
74226	 => std_logic_vector(to_unsigned(33,8) ,
74227	 => std_logic_vector(to_unsigned(28,8) ,
74228	 => std_logic_vector(to_unsigned(24,8) ,
74229	 => std_logic_vector(to_unsigned(12,8) ,
74230	 => std_logic_vector(to_unsigned(8,8) ,
74231	 => std_logic_vector(to_unsigned(10,8) ,
74232	 => std_logic_vector(to_unsigned(14,8) ,
74233	 => std_logic_vector(to_unsigned(23,8) ,
74234	 => std_logic_vector(to_unsigned(26,8) ,
74235	 => std_logic_vector(to_unsigned(56,8) ,
74236	 => std_logic_vector(to_unsigned(66,8) ,
74237	 => std_logic_vector(to_unsigned(74,8) ,
74238	 => std_logic_vector(to_unsigned(80,8) ,
74239	 => std_logic_vector(to_unsigned(67,8) ,
74240	 => std_logic_vector(to_unsigned(58,8) ,
74241	 => std_logic_vector(to_unsigned(124,8) ,
74242	 => std_logic_vector(to_unsigned(111,8) ,
74243	 => std_logic_vector(to_unsigned(108,8) ,
74244	 => std_logic_vector(to_unsigned(99,8) ,
74245	 => std_logic_vector(to_unsigned(111,8) ,
74246	 => std_logic_vector(to_unsigned(133,8) ,
74247	 => std_logic_vector(to_unsigned(131,8) ,
74248	 => std_logic_vector(to_unsigned(128,8) ,
74249	 => std_logic_vector(to_unsigned(133,8) ,
74250	 => std_logic_vector(to_unsigned(112,8) ,
74251	 => std_logic_vector(to_unsigned(91,8) ,
74252	 => std_logic_vector(to_unsigned(81,8) ,
74253	 => std_logic_vector(to_unsigned(86,8) ,
74254	 => std_logic_vector(to_unsigned(84,8) ,
74255	 => std_logic_vector(to_unsigned(82,8) ,
74256	 => std_logic_vector(to_unsigned(85,8) ,
74257	 => std_logic_vector(to_unsigned(81,8) ,
74258	 => std_logic_vector(to_unsigned(61,8) ,
74259	 => std_logic_vector(to_unsigned(57,8) ,
74260	 => std_logic_vector(to_unsigned(63,8) ,
74261	 => std_logic_vector(to_unsigned(54,8) ,
74262	 => std_logic_vector(to_unsigned(60,8) ,
74263	 => std_logic_vector(to_unsigned(35,8) ,
74264	 => std_logic_vector(to_unsigned(60,8) ,
74265	 => std_logic_vector(to_unsigned(57,8) ,
74266	 => std_logic_vector(to_unsigned(30,8) ,
74267	 => std_logic_vector(to_unsigned(38,8) ,
74268	 => std_logic_vector(to_unsigned(49,8) ,
74269	 => std_logic_vector(to_unsigned(37,8) ,
74270	 => std_logic_vector(to_unsigned(45,8) ,
74271	 => std_logic_vector(to_unsigned(62,8) ,
74272	 => std_logic_vector(to_unsigned(51,8) ,
74273	 => std_logic_vector(to_unsigned(62,8) ,
74274	 => std_logic_vector(to_unsigned(62,8) ,
74275	 => std_logic_vector(to_unsigned(40,8) ,
74276	 => std_logic_vector(to_unsigned(35,8) ,
74277	 => std_logic_vector(to_unsigned(37,8) ,
74278	 => std_logic_vector(to_unsigned(30,8) ,
74279	 => std_logic_vector(to_unsigned(33,8) ,
74280	 => std_logic_vector(to_unsigned(20,8) ,
74281	 => std_logic_vector(to_unsigned(11,8) ,
74282	 => std_logic_vector(to_unsigned(29,8) ,
74283	 => std_logic_vector(to_unsigned(67,8) ,
74284	 => std_logic_vector(to_unsigned(70,8) ,
74285	 => std_logic_vector(to_unsigned(72,8) ,
74286	 => std_logic_vector(to_unsigned(69,8) ,
74287	 => std_logic_vector(to_unsigned(63,8) ,
74288	 => std_logic_vector(to_unsigned(48,8) ,
74289	 => std_logic_vector(to_unsigned(47,8) ,
74290	 => std_logic_vector(to_unsigned(53,8) ,
74291	 => std_logic_vector(to_unsigned(67,8) ,
74292	 => std_logic_vector(to_unsigned(86,8) ,
74293	 => std_logic_vector(to_unsigned(101,8) ,
74294	 => std_logic_vector(to_unsigned(100,8) ,
74295	 => std_logic_vector(to_unsigned(99,8) ,
74296	 => std_logic_vector(to_unsigned(100,8) ,
74297	 => std_logic_vector(to_unsigned(104,8) ,
74298	 => std_logic_vector(to_unsigned(103,8) ,
74299	 => std_logic_vector(to_unsigned(96,8) ,
74300	 => std_logic_vector(to_unsigned(93,8) ,
74301	 => std_logic_vector(to_unsigned(112,8) ,
74302	 => std_logic_vector(to_unsigned(71,8) ,
74303	 => std_logic_vector(to_unsigned(61,8) ,
74304	 => std_logic_vector(to_unsigned(104,8) ,
74305	 => std_logic_vector(to_unsigned(141,8) ,
74306	 => std_logic_vector(to_unsigned(95,8) ,
74307	 => std_logic_vector(to_unsigned(51,8) ,
74308	 => std_logic_vector(to_unsigned(36,8) ,
74309	 => std_logic_vector(to_unsigned(35,8) ,
74310	 => std_logic_vector(to_unsigned(36,8) ,
74311	 => std_logic_vector(to_unsigned(33,8) ,
74312	 => std_logic_vector(to_unsigned(37,8) ,
74313	 => std_logic_vector(to_unsigned(35,8) ,
74314	 => std_logic_vector(to_unsigned(39,8) ,
74315	 => std_logic_vector(to_unsigned(32,8) ,
74316	 => std_logic_vector(to_unsigned(33,8) ,
74317	 => std_logic_vector(to_unsigned(35,8) ,
74318	 => std_logic_vector(to_unsigned(31,8) ,
74319	 => std_logic_vector(to_unsigned(61,8) ,
74320	 => std_logic_vector(to_unsigned(86,8) ,
74321	 => std_logic_vector(to_unsigned(105,8) ,
74322	 => std_logic_vector(to_unsigned(95,8) ,
74323	 => std_logic_vector(to_unsigned(114,8) ,
74324	 => std_logic_vector(to_unsigned(92,8) ,
74325	 => std_logic_vector(to_unsigned(128,8) ,
74326	 => std_logic_vector(to_unsigned(96,8) ,
74327	 => std_logic_vector(to_unsigned(119,8) ,
74328	 => std_logic_vector(to_unsigned(95,8) ,
74329	 => std_logic_vector(to_unsigned(109,8) ,
74330	 => std_logic_vector(to_unsigned(85,8) ,
74331	 => std_logic_vector(to_unsigned(95,8) ,
74332	 => std_logic_vector(to_unsigned(68,8) ,
74333	 => std_logic_vector(to_unsigned(51,8) ,
74334	 => std_logic_vector(to_unsigned(50,8) ,
74335	 => std_logic_vector(to_unsigned(38,8) ,
74336	 => std_logic_vector(to_unsigned(37,8) ,
74337	 => std_logic_vector(to_unsigned(35,8) ,
74338	 => std_logic_vector(to_unsigned(32,8) ,
74339	 => std_logic_vector(to_unsigned(58,8) ,
74340	 => std_logic_vector(to_unsigned(90,8) ,
74341	 => std_logic_vector(to_unsigned(88,8) ,
74342	 => std_logic_vector(to_unsigned(72,8) ,
74343	 => std_logic_vector(to_unsigned(65,8) ,
74344	 => std_logic_vector(to_unsigned(97,8) ,
74345	 => std_logic_vector(to_unsigned(72,8) ,
74346	 => std_logic_vector(to_unsigned(95,8) ,
74347	 => std_logic_vector(to_unsigned(133,8) ,
74348	 => std_logic_vector(to_unsigned(87,8) ,
74349	 => std_logic_vector(to_unsigned(109,8) ,
74350	 => std_logic_vector(to_unsigned(130,8) ,
74351	 => std_logic_vector(to_unsigned(104,8) ,
74352	 => std_logic_vector(to_unsigned(114,8) ,
74353	 => std_logic_vector(to_unsigned(108,8) ,
74354	 => std_logic_vector(to_unsigned(91,8) ,
74355	 => std_logic_vector(to_unsigned(77,8) ,
74356	 => std_logic_vector(to_unsigned(60,8) ,
74357	 => std_logic_vector(to_unsigned(65,8) ,
74358	 => std_logic_vector(to_unsigned(97,8) ,
74359	 => std_logic_vector(to_unsigned(100,8) ,
74360	 => std_logic_vector(to_unsigned(105,8) ,
74361	 => std_logic_vector(to_unsigned(111,8) ,
74362	 => std_logic_vector(to_unsigned(105,8) ,
74363	 => std_logic_vector(to_unsigned(99,8) ,
74364	 => std_logic_vector(to_unsigned(99,8) ,
74365	 => std_logic_vector(to_unsigned(96,8) ,
74366	 => std_logic_vector(to_unsigned(99,8) ,
74367	 => std_logic_vector(to_unsigned(104,8) ,
74368	 => std_logic_vector(to_unsigned(70,8) ,
74369	 => std_logic_vector(to_unsigned(35,8) ,
74370	 => std_logic_vector(to_unsigned(24,8) ,
74371	 => std_logic_vector(to_unsigned(9,8) ,
74372	 => std_logic_vector(to_unsigned(10,8) ,
74373	 => std_logic_vector(to_unsigned(19,8) ,
74374	 => std_logic_vector(to_unsigned(29,8) ,
74375	 => std_logic_vector(to_unsigned(44,8) ,
74376	 => std_logic_vector(to_unsigned(38,8) ,
74377	 => std_logic_vector(to_unsigned(51,8) ,
74378	 => std_logic_vector(to_unsigned(82,8) ,
74379	 => std_logic_vector(to_unsigned(77,8) ,
74380	 => std_logic_vector(to_unsigned(66,8) ,
74381	 => std_logic_vector(to_unsigned(80,8) ,
74382	 => std_logic_vector(to_unsigned(74,8) ,
74383	 => std_logic_vector(to_unsigned(68,8) ,
74384	 => std_logic_vector(to_unsigned(80,8) ,
74385	 => std_logic_vector(to_unsigned(80,8) ,
74386	 => std_logic_vector(to_unsigned(69,8) ,
74387	 => std_logic_vector(to_unsigned(77,8) ,
74388	 => std_logic_vector(to_unsigned(84,8) ,
74389	 => std_logic_vector(to_unsigned(66,8) ,
74390	 => std_logic_vector(to_unsigned(92,8) ,
74391	 => std_logic_vector(to_unsigned(84,8) ,
74392	 => std_logic_vector(to_unsigned(35,8) ,
74393	 => std_logic_vector(to_unsigned(77,8) ,
74394	 => std_logic_vector(to_unsigned(93,8) ,
74395	 => std_logic_vector(to_unsigned(85,8) ,
74396	 => std_logic_vector(to_unsigned(80,8) ,
74397	 => std_logic_vector(to_unsigned(72,8) ,
74398	 => std_logic_vector(to_unsigned(62,8) ,
74399	 => std_logic_vector(to_unsigned(44,8) ,
74400	 => std_logic_vector(to_unsigned(48,8) ,
74401	 => std_logic_vector(to_unsigned(14,8) ,
74402	 => std_logic_vector(to_unsigned(28,8) ,
74403	 => std_logic_vector(to_unsigned(63,8) ,
74404	 => std_logic_vector(to_unsigned(76,8) ,
74405	 => std_logic_vector(to_unsigned(73,8) ,
74406	 => std_logic_vector(to_unsigned(32,8) ,
74407	 => std_logic_vector(to_unsigned(7,8) ,
74408	 => std_logic_vector(to_unsigned(5,8) ,
74409	 => std_logic_vector(to_unsigned(12,8) ,
74410	 => std_logic_vector(to_unsigned(11,8) ,
74411	 => std_logic_vector(to_unsigned(27,8) ,
74412	 => std_logic_vector(to_unsigned(41,8) ,
74413	 => std_logic_vector(to_unsigned(15,8) ,
74414	 => std_logic_vector(to_unsigned(50,8) ,
74415	 => std_logic_vector(to_unsigned(64,8) ,
74416	 => std_logic_vector(to_unsigned(66,8) ,
74417	 => std_logic_vector(to_unsigned(18,8) ,
74418	 => std_logic_vector(to_unsigned(2,8) ,
74419	 => std_logic_vector(to_unsigned(5,8) ,
74420	 => std_logic_vector(to_unsigned(8,8) ,
74421	 => std_logic_vector(to_unsigned(22,8) ,
74422	 => std_logic_vector(to_unsigned(32,8) ,
74423	 => std_logic_vector(to_unsigned(15,8) ,
74424	 => std_logic_vector(to_unsigned(16,8) ,
74425	 => std_logic_vector(to_unsigned(7,8) ,
74426	 => std_logic_vector(to_unsigned(19,8) ,
74427	 => std_logic_vector(to_unsigned(22,8) ,
74428	 => std_logic_vector(to_unsigned(7,8) ,
74429	 => std_logic_vector(to_unsigned(8,8) ,
74430	 => std_logic_vector(to_unsigned(20,8) ,
74431	 => std_logic_vector(to_unsigned(28,8) ,
74432	 => std_logic_vector(to_unsigned(27,8) ,
74433	 => std_logic_vector(to_unsigned(29,8) ,
74434	 => std_logic_vector(to_unsigned(32,8) ,
74435	 => std_logic_vector(to_unsigned(26,8) ,
74436	 => std_logic_vector(to_unsigned(23,8) ,
74437	 => std_logic_vector(to_unsigned(24,8) ,
74438	 => std_logic_vector(to_unsigned(24,8) ,
74439	 => std_logic_vector(to_unsigned(20,8) ,
74440	 => std_logic_vector(to_unsigned(23,8) ,
74441	 => std_logic_vector(to_unsigned(22,8) ,
74442	 => std_logic_vector(to_unsigned(10,8) ,
74443	 => std_logic_vector(to_unsigned(7,8) ,
74444	 => std_logic_vector(to_unsigned(13,8) ,
74445	 => std_logic_vector(to_unsigned(13,8) ,
74446	 => std_logic_vector(to_unsigned(9,8) ,
74447	 => std_logic_vector(to_unsigned(8,8) ,
74448	 => std_logic_vector(to_unsigned(17,8) ,
74449	 => std_logic_vector(to_unsigned(25,8) ,
74450	 => std_logic_vector(to_unsigned(30,8) ,
74451	 => std_logic_vector(to_unsigned(25,8) ,
74452	 => std_logic_vector(to_unsigned(17,8) ,
74453	 => std_logic_vector(to_unsigned(18,8) ,
74454	 => std_logic_vector(to_unsigned(16,8) ,
74455	 => std_logic_vector(to_unsigned(15,8) ,
74456	 => std_logic_vector(to_unsigned(13,8) ,
74457	 => std_logic_vector(to_unsigned(16,8) ,
74458	 => std_logic_vector(to_unsigned(18,8) ,
74459	 => std_logic_vector(to_unsigned(21,8) ,
74460	 => std_logic_vector(to_unsigned(34,8) ,
74461	 => std_logic_vector(to_unsigned(35,8) ,
74462	 => std_logic_vector(to_unsigned(20,8) ,
74463	 => std_logic_vector(to_unsigned(23,8) ,
74464	 => std_logic_vector(to_unsigned(33,8) ,
74465	 => std_logic_vector(to_unsigned(28,8) ,
74466	 => std_logic_vector(to_unsigned(27,8) ,
74467	 => std_logic_vector(to_unsigned(24,8) ,
74468	 => std_logic_vector(to_unsigned(9,8) ,
74469	 => std_logic_vector(to_unsigned(3,8) ,
74470	 => std_logic_vector(to_unsigned(16,8) ,
74471	 => std_logic_vector(to_unsigned(31,8) ,
74472	 => std_logic_vector(to_unsigned(20,8) ,
74473	 => std_logic_vector(to_unsigned(16,8) ,
74474	 => std_logic_vector(to_unsigned(32,8) ,
74475	 => std_logic_vector(to_unsigned(34,8) ,
74476	 => std_logic_vector(to_unsigned(22,8) ,
74477	 => std_logic_vector(to_unsigned(20,8) ,
74478	 => std_logic_vector(to_unsigned(30,8) ,
74479	 => std_logic_vector(to_unsigned(21,8) ,
74480	 => std_logic_vector(to_unsigned(20,8) ,
74481	 => std_logic_vector(to_unsigned(21,8) ,
74482	 => std_logic_vector(to_unsigned(30,8) ,
74483	 => std_logic_vector(to_unsigned(23,8) ,
74484	 => std_logic_vector(to_unsigned(19,8) ,
74485	 => std_logic_vector(to_unsigned(12,8) ,
74486	 => std_logic_vector(to_unsigned(18,8) ,
74487	 => std_logic_vector(to_unsigned(54,8) ,
74488	 => std_logic_vector(to_unsigned(10,8) ,
74489	 => std_logic_vector(to_unsigned(5,8) ,
74490	 => std_logic_vector(to_unsigned(12,8) ,
74491	 => std_logic_vector(to_unsigned(12,8) ,
74492	 => std_logic_vector(to_unsigned(11,8) ,
74493	 => std_logic_vector(to_unsigned(12,8) ,
74494	 => std_logic_vector(to_unsigned(18,8) ,
74495	 => std_logic_vector(to_unsigned(25,8) ,
74496	 => std_logic_vector(to_unsigned(24,8) ,
74497	 => std_logic_vector(to_unsigned(13,8) ,
74498	 => std_logic_vector(to_unsigned(11,8) ,
74499	 => std_logic_vector(to_unsigned(12,8) ,
74500	 => std_logic_vector(to_unsigned(11,8) ,
74501	 => std_logic_vector(to_unsigned(7,8) ,
74502	 => std_logic_vector(to_unsigned(4,8) ,
74503	 => std_logic_vector(to_unsigned(6,8) ,
74504	 => std_logic_vector(to_unsigned(13,8) ,
74505	 => std_logic_vector(to_unsigned(24,8) ,
74506	 => std_logic_vector(to_unsigned(25,8) ,
74507	 => std_logic_vector(to_unsigned(17,8) ,
74508	 => std_logic_vector(to_unsigned(12,8) ,
74509	 => std_logic_vector(to_unsigned(22,8) ,
74510	 => std_logic_vector(to_unsigned(32,8) ,
74511	 => std_logic_vector(to_unsigned(18,8) ,
74512	 => std_logic_vector(to_unsigned(13,8) ,
74513	 => std_logic_vector(to_unsigned(10,8) ,
74514	 => std_logic_vector(to_unsigned(10,8) ,
74515	 => std_logic_vector(to_unsigned(8,8) ,
74516	 => std_logic_vector(to_unsigned(8,8) ,
74517	 => std_logic_vector(to_unsigned(16,8) ,
74518	 => std_logic_vector(to_unsigned(27,8) ,
74519	 => std_logic_vector(to_unsigned(12,8) ,
74520	 => std_logic_vector(to_unsigned(0,8) ,
74521	 => std_logic_vector(to_unsigned(0,8) ,
74522	 => std_logic_vector(to_unsigned(3,8) ,
74523	 => std_logic_vector(to_unsigned(19,8) ,
74524	 => std_logic_vector(to_unsigned(30,8) ,
74525	 => std_logic_vector(to_unsigned(26,8) ,
74526	 => std_logic_vector(to_unsigned(19,8) ,
74527	 => std_logic_vector(to_unsigned(22,8) ,
74528	 => std_logic_vector(to_unsigned(35,8) ,
74529	 => std_logic_vector(to_unsigned(35,8) ,
74530	 => std_logic_vector(to_unsigned(13,8) ,
74531	 => std_logic_vector(to_unsigned(18,8) ,
74532	 => std_logic_vector(to_unsigned(28,8) ,
74533	 => std_logic_vector(to_unsigned(22,8) ,
74534	 => std_logic_vector(to_unsigned(8,8) ,
74535	 => std_logic_vector(to_unsigned(2,8) ,
74536	 => std_logic_vector(to_unsigned(0,8) ,
74537	 => std_logic_vector(to_unsigned(0,8) ,
74538	 => std_logic_vector(to_unsigned(1,8) ,
74539	 => std_logic_vector(to_unsigned(1,8) ,
74540	 => std_logic_vector(to_unsigned(1,8) ,
74541	 => std_logic_vector(to_unsigned(5,8) ,
74542	 => std_logic_vector(to_unsigned(18,8) ,
74543	 => std_logic_vector(to_unsigned(24,8) ,
74544	 => std_logic_vector(to_unsigned(41,8) ,
74545	 => std_logic_vector(to_unsigned(47,8) ,
74546	 => std_logic_vector(to_unsigned(53,8) ,
74547	 => std_logic_vector(to_unsigned(51,8) ,
74548	 => std_logic_vector(to_unsigned(41,8) ,
74549	 => std_logic_vector(to_unsigned(14,8) ,
74550	 => std_logic_vector(to_unsigned(13,8) ,
74551	 => std_logic_vector(to_unsigned(11,8) ,
74552	 => std_logic_vector(to_unsigned(13,8) ,
74553	 => std_logic_vector(to_unsigned(11,8) ,
74554	 => std_logic_vector(to_unsigned(22,8) ,
74555	 => std_logic_vector(to_unsigned(48,8) ,
74556	 => std_logic_vector(to_unsigned(48,8) ,
74557	 => std_logic_vector(to_unsigned(51,8) ,
74558	 => std_logic_vector(to_unsigned(54,8) ,
74559	 => std_logic_vector(to_unsigned(66,8) ,
74560	 => std_logic_vector(to_unsigned(80,8) ,
74561	 => std_logic_vector(to_unsigned(128,8) ,
74562	 => std_logic_vector(to_unsigned(121,8) ,
74563	 => std_logic_vector(to_unsigned(118,8) ,
74564	 => std_logic_vector(to_unsigned(112,8) ,
74565	 => std_logic_vector(to_unsigned(108,8) ,
74566	 => std_logic_vector(to_unsigned(111,8) ,
74567	 => std_logic_vector(to_unsigned(115,8) ,
74568	 => std_logic_vector(to_unsigned(114,8) ,
74569	 => std_logic_vector(to_unsigned(108,8) ,
74570	 => std_logic_vector(to_unsigned(92,8) ,
74571	 => std_logic_vector(to_unsigned(88,8) ,
74572	 => std_logic_vector(to_unsigned(87,8) ,
74573	 => std_logic_vector(to_unsigned(90,8) ,
74574	 => std_logic_vector(to_unsigned(90,8) ,
74575	 => std_logic_vector(to_unsigned(80,8) ,
74576	 => std_logic_vector(to_unsigned(72,8) ,
74577	 => std_logic_vector(to_unsigned(69,8) ,
74578	 => std_logic_vector(to_unsigned(59,8) ,
74579	 => std_logic_vector(to_unsigned(58,8) ,
74580	 => std_logic_vector(to_unsigned(65,8) ,
74581	 => std_logic_vector(to_unsigned(51,8) ,
74582	 => std_logic_vector(to_unsigned(44,8) ,
74583	 => std_logic_vector(to_unsigned(34,8) ,
74584	 => std_logic_vector(to_unsigned(42,8) ,
74585	 => std_logic_vector(to_unsigned(41,8) ,
74586	 => std_logic_vector(to_unsigned(36,8) ,
74587	 => std_logic_vector(to_unsigned(49,8) ,
74588	 => std_logic_vector(to_unsigned(50,8) ,
74589	 => std_logic_vector(to_unsigned(51,8) ,
74590	 => std_logic_vector(to_unsigned(54,8) ,
74591	 => std_logic_vector(to_unsigned(53,8) ,
74592	 => std_logic_vector(to_unsigned(58,8) ,
74593	 => std_logic_vector(to_unsigned(49,8) ,
74594	 => std_logic_vector(to_unsigned(35,8) ,
74595	 => std_logic_vector(to_unsigned(34,8) ,
74596	 => std_logic_vector(to_unsigned(37,8) ,
74597	 => std_logic_vector(to_unsigned(48,8) ,
74598	 => std_logic_vector(to_unsigned(45,8) ,
74599	 => std_logic_vector(to_unsigned(43,8) ,
74600	 => std_logic_vector(to_unsigned(36,8) ,
74601	 => std_logic_vector(to_unsigned(25,8) ,
74602	 => std_logic_vector(to_unsigned(24,8) ,
74603	 => std_logic_vector(to_unsigned(33,8) ,
74604	 => std_logic_vector(to_unsigned(45,8) ,
74605	 => std_logic_vector(to_unsigned(69,8) ,
74606	 => std_logic_vector(to_unsigned(73,8) ,
74607	 => std_logic_vector(to_unsigned(73,8) ,
74608	 => std_logic_vector(to_unsigned(70,8) ,
74609	 => std_logic_vector(to_unsigned(65,8) ,
74610	 => std_logic_vector(to_unsigned(91,8) ,
74611	 => std_logic_vector(to_unsigned(99,8) ,
74612	 => std_logic_vector(to_unsigned(91,8) ,
74613	 => std_logic_vector(to_unsigned(97,8) ,
74614	 => std_logic_vector(to_unsigned(100,8) ,
74615	 => std_logic_vector(to_unsigned(105,8) ,
74616	 => std_logic_vector(to_unsigned(104,8) ,
74617	 => std_logic_vector(to_unsigned(104,8) ,
74618	 => std_logic_vector(to_unsigned(105,8) ,
74619	 => std_logic_vector(to_unsigned(104,8) ,
74620	 => std_logic_vector(to_unsigned(91,8) ,
74621	 => std_logic_vector(to_unsigned(95,8) ,
74622	 => std_logic_vector(to_unsigned(84,8) ,
74623	 => std_logic_vector(to_unsigned(71,8) ,
74624	 => std_logic_vector(to_unsigned(85,8) ,
74625	 => std_logic_vector(to_unsigned(82,8) ,
74626	 => std_logic_vector(to_unsigned(59,8) ,
74627	 => std_logic_vector(to_unsigned(58,8) ,
74628	 => std_logic_vector(to_unsigned(45,8) ,
74629	 => std_logic_vector(to_unsigned(32,8) ,
74630	 => std_logic_vector(to_unsigned(37,8) ,
74631	 => std_logic_vector(to_unsigned(37,8) ,
74632	 => std_logic_vector(to_unsigned(34,8) ,
74633	 => std_logic_vector(to_unsigned(35,8) ,
74634	 => std_logic_vector(to_unsigned(39,8) ,
74635	 => std_logic_vector(to_unsigned(45,8) ,
74636	 => std_logic_vector(to_unsigned(41,8) ,
74637	 => std_logic_vector(to_unsigned(34,8) ,
74638	 => std_logic_vector(to_unsigned(29,8) ,
74639	 => std_logic_vector(to_unsigned(55,8) ,
74640	 => std_logic_vector(to_unsigned(62,8) ,
74641	 => std_logic_vector(to_unsigned(67,8) ,
74642	 => std_logic_vector(to_unsigned(50,8) ,
74643	 => std_logic_vector(to_unsigned(74,8) ,
74644	 => std_logic_vector(to_unsigned(73,8) ,
74645	 => std_logic_vector(to_unsigned(116,8) ,
74646	 => std_logic_vector(to_unsigned(85,8) ,
74647	 => std_logic_vector(to_unsigned(104,8) ,
74648	 => std_logic_vector(to_unsigned(80,8) ,
74649	 => std_logic_vector(to_unsigned(107,8) ,
74650	 => std_logic_vector(to_unsigned(82,8) ,
74651	 => std_logic_vector(to_unsigned(121,8) ,
74652	 => std_logic_vector(to_unsigned(61,8) ,
74653	 => std_logic_vector(to_unsigned(86,8) ,
74654	 => std_logic_vector(to_unsigned(70,8) ,
74655	 => std_logic_vector(to_unsigned(79,8) ,
74656	 => std_logic_vector(to_unsigned(84,8) ,
74657	 => std_logic_vector(to_unsigned(57,8) ,
74658	 => std_logic_vector(to_unsigned(51,8) ,
74659	 => std_logic_vector(to_unsigned(43,8) ,
74660	 => std_logic_vector(to_unsigned(38,8) ,
74661	 => std_logic_vector(to_unsigned(48,8) ,
74662	 => std_logic_vector(to_unsigned(55,8) ,
74663	 => std_logic_vector(to_unsigned(57,8) ,
74664	 => std_logic_vector(to_unsigned(97,8) ,
74665	 => std_logic_vector(to_unsigned(63,8) ,
74666	 => std_logic_vector(to_unsigned(74,8) ,
74667	 => std_logic_vector(to_unsigned(136,8) ,
74668	 => std_logic_vector(to_unsigned(41,8) ,
74669	 => std_logic_vector(to_unsigned(50,8) ,
74670	 => std_logic_vector(to_unsigned(124,8) ,
74671	 => std_logic_vector(to_unsigned(40,8) ,
74672	 => std_logic_vector(to_unsigned(63,8) ,
74673	 => std_logic_vector(to_unsigned(116,8) ,
74674	 => std_logic_vector(to_unsigned(86,8) ,
74675	 => std_logic_vector(to_unsigned(78,8) ,
74676	 => std_logic_vector(to_unsigned(57,8) ,
74677	 => std_logic_vector(to_unsigned(62,8) ,
74678	 => std_logic_vector(to_unsigned(91,8) ,
74679	 => std_logic_vector(to_unsigned(92,8) ,
74680	 => std_logic_vector(to_unsigned(100,8) ,
74681	 => std_logic_vector(to_unsigned(111,8) ,
74682	 => std_logic_vector(to_unsigned(104,8) ,
74683	 => std_logic_vector(to_unsigned(100,8) ,
74684	 => std_logic_vector(to_unsigned(103,8) ,
74685	 => std_logic_vector(to_unsigned(101,8) ,
74686	 => std_logic_vector(to_unsigned(99,8) ,
74687	 => std_logic_vector(to_unsigned(97,8) ,
74688	 => std_logic_vector(to_unsigned(86,8) ,
74689	 => std_logic_vector(to_unsigned(55,8) ,
74690	 => std_logic_vector(to_unsigned(17,8) ,
74691	 => std_logic_vector(to_unsigned(6,8) ,
74692	 => std_logic_vector(to_unsigned(5,8) ,
74693	 => std_logic_vector(to_unsigned(5,8) ,
74694	 => std_logic_vector(to_unsigned(8,8) ,
74695	 => std_logic_vector(to_unsigned(8,8) ,
74696	 => std_logic_vector(to_unsigned(8,8) ,
74697	 => std_logic_vector(to_unsigned(45,8) ,
74698	 => std_logic_vector(to_unsigned(41,8) ,
74699	 => std_logic_vector(to_unsigned(57,8) ,
74700	 => std_logic_vector(to_unsigned(46,8) ,
74701	 => std_logic_vector(to_unsigned(61,8) ,
74702	 => std_logic_vector(to_unsigned(80,8) ,
74703	 => std_logic_vector(to_unsigned(76,8) ,
74704	 => std_logic_vector(to_unsigned(79,8) ,
74705	 => std_logic_vector(to_unsigned(73,8) ,
74706	 => std_logic_vector(to_unsigned(73,8) ,
74707	 => std_logic_vector(to_unsigned(78,8) ,
74708	 => std_logic_vector(to_unsigned(84,8) ,
74709	 => std_logic_vector(to_unsigned(80,8) ,
74710	 => std_logic_vector(to_unsigned(88,8) ,
74711	 => std_logic_vector(to_unsigned(81,8) ,
74712	 => std_logic_vector(to_unsigned(17,8) ,
74713	 => std_logic_vector(to_unsigned(68,8) ,
74714	 => std_logic_vector(to_unsigned(111,8) ,
74715	 => std_logic_vector(to_unsigned(84,8) ,
74716	 => std_logic_vector(to_unsigned(77,8) ,
74717	 => std_logic_vector(to_unsigned(74,8) ,
74718	 => std_logic_vector(to_unsigned(55,8) ,
74719	 => std_logic_vector(to_unsigned(26,8) ,
74720	 => std_logic_vector(to_unsigned(43,8) ,
74721	 => std_logic_vector(to_unsigned(45,8) ,
74722	 => std_logic_vector(to_unsigned(51,8) ,
74723	 => std_logic_vector(to_unsigned(72,8) ,
74724	 => std_logic_vector(to_unsigned(80,8) ,
74725	 => std_logic_vector(to_unsigned(80,8) ,
74726	 => std_logic_vector(to_unsigned(28,8) ,
74727	 => std_logic_vector(to_unsigned(6,8) ,
74728	 => std_logic_vector(to_unsigned(6,8) ,
74729	 => std_logic_vector(to_unsigned(12,8) ,
74730	 => std_logic_vector(to_unsigned(11,8) ,
74731	 => std_logic_vector(to_unsigned(19,8) ,
74732	 => std_logic_vector(to_unsigned(30,8) ,
74733	 => std_logic_vector(to_unsigned(52,8) ,
74734	 => std_logic_vector(to_unsigned(68,8) ,
74735	 => std_logic_vector(to_unsigned(51,8) ,
74736	 => std_logic_vector(to_unsigned(30,8) ,
74737	 => std_logic_vector(to_unsigned(4,8) ,
74738	 => std_logic_vector(to_unsigned(6,8) ,
74739	 => std_logic_vector(to_unsigned(17,8) ,
74740	 => std_logic_vector(to_unsigned(21,8) ,
74741	 => std_logic_vector(to_unsigned(19,8) ,
74742	 => std_logic_vector(to_unsigned(25,8) ,
74743	 => std_logic_vector(to_unsigned(14,8) ,
74744	 => std_logic_vector(to_unsigned(9,8) ,
74745	 => std_logic_vector(to_unsigned(6,8) ,
74746	 => std_logic_vector(to_unsigned(16,8) ,
74747	 => std_logic_vector(to_unsigned(33,8) ,
74748	 => std_logic_vector(to_unsigned(24,8) ,
74749	 => std_logic_vector(to_unsigned(17,8) ,
74750	 => std_logic_vector(to_unsigned(24,8) ,
74751	 => std_logic_vector(to_unsigned(29,8) ,
74752	 => std_logic_vector(to_unsigned(13,8) ,
74753	 => std_logic_vector(to_unsigned(8,8) ,
74754	 => std_logic_vector(to_unsigned(12,8) ,
74755	 => std_logic_vector(to_unsigned(22,8) ,
74756	 => std_logic_vector(to_unsigned(22,8) ,
74757	 => std_logic_vector(to_unsigned(21,8) ,
74758	 => std_logic_vector(to_unsigned(27,8) ,
74759	 => std_logic_vector(to_unsigned(29,8) ,
74760	 => std_logic_vector(to_unsigned(21,8) ,
74761	 => std_logic_vector(to_unsigned(16,8) ,
74762	 => std_logic_vector(to_unsigned(10,8) ,
74763	 => std_logic_vector(to_unsigned(9,8) ,
74764	 => std_logic_vector(to_unsigned(11,8) ,
74765	 => std_logic_vector(to_unsigned(12,8) ,
74766	 => std_logic_vector(to_unsigned(8,8) ,
74767	 => std_logic_vector(to_unsigned(9,8) ,
74768	 => std_logic_vector(to_unsigned(17,8) ,
74769	 => std_logic_vector(to_unsigned(42,8) ,
74770	 => std_logic_vector(to_unsigned(53,8) ,
74771	 => std_logic_vector(to_unsigned(34,8) ,
74772	 => std_logic_vector(to_unsigned(17,8) ,
74773	 => std_logic_vector(to_unsigned(17,8) ,
74774	 => std_logic_vector(to_unsigned(25,8) ,
74775	 => std_logic_vector(to_unsigned(33,8) ,
74776	 => std_logic_vector(to_unsigned(27,8) ,
74777	 => std_logic_vector(to_unsigned(18,8) ,
74778	 => std_logic_vector(to_unsigned(18,8) ,
74779	 => std_logic_vector(to_unsigned(18,8) ,
74780	 => std_logic_vector(to_unsigned(23,8) ,
74781	 => std_logic_vector(to_unsigned(29,8) ,
74782	 => std_logic_vector(to_unsigned(17,8) ,
74783	 => std_logic_vector(to_unsigned(20,8) ,
74784	 => std_logic_vector(to_unsigned(27,8) ,
74785	 => std_logic_vector(to_unsigned(27,8) ,
74786	 => std_logic_vector(to_unsigned(26,8) ,
74787	 => std_logic_vector(to_unsigned(20,8) ,
74788	 => std_logic_vector(to_unsigned(9,8) ,
74789	 => std_logic_vector(to_unsigned(2,8) ,
74790	 => std_logic_vector(to_unsigned(13,8) ,
74791	 => std_logic_vector(to_unsigned(13,8) ,
74792	 => std_logic_vector(to_unsigned(9,8) ,
74793	 => std_logic_vector(to_unsigned(9,8) ,
74794	 => std_logic_vector(to_unsigned(22,8) ,
74795	 => std_logic_vector(to_unsigned(30,8) ,
74796	 => std_logic_vector(to_unsigned(25,8) ,
74797	 => std_logic_vector(to_unsigned(23,8) ,
74798	 => std_logic_vector(to_unsigned(36,8) ,
74799	 => std_logic_vector(to_unsigned(38,8) ,
74800	 => std_logic_vector(to_unsigned(33,8) ,
74801	 => std_logic_vector(to_unsigned(27,8) ,
74802	 => std_logic_vector(to_unsigned(17,8) ,
74803	 => std_logic_vector(to_unsigned(13,8) ,
74804	 => std_logic_vector(to_unsigned(13,8) ,
74805	 => std_logic_vector(to_unsigned(12,8) ,
74806	 => std_logic_vector(to_unsigned(46,8) ,
74807	 => std_logic_vector(to_unsigned(37,8) ,
74808	 => std_logic_vector(to_unsigned(3,8) ,
74809	 => std_logic_vector(to_unsigned(4,8) ,
74810	 => std_logic_vector(to_unsigned(4,8) ,
74811	 => std_logic_vector(to_unsigned(5,8) ,
74812	 => std_logic_vector(to_unsigned(7,8) ,
74813	 => std_logic_vector(to_unsigned(8,8) ,
74814	 => std_logic_vector(to_unsigned(8,8) ,
74815	 => std_logic_vector(to_unsigned(18,8) ,
74816	 => std_logic_vector(to_unsigned(20,8) ,
74817	 => std_logic_vector(to_unsigned(8,8) ,
74818	 => std_logic_vector(to_unsigned(7,8) ,
74819	 => std_logic_vector(to_unsigned(9,8) ,
74820	 => std_logic_vector(to_unsigned(8,8) ,
74821	 => std_logic_vector(to_unsigned(5,8) ,
74822	 => std_logic_vector(to_unsigned(3,8) ,
74823	 => std_logic_vector(to_unsigned(10,8) ,
74824	 => std_logic_vector(to_unsigned(24,8) ,
74825	 => std_logic_vector(to_unsigned(29,8) ,
74826	 => std_logic_vector(to_unsigned(21,8) ,
74827	 => std_logic_vector(to_unsigned(11,8) ,
74828	 => std_logic_vector(to_unsigned(13,8) ,
74829	 => std_logic_vector(to_unsigned(16,8) ,
74830	 => std_logic_vector(to_unsigned(28,8) ,
74831	 => std_logic_vector(to_unsigned(20,8) ,
74832	 => std_logic_vector(to_unsigned(17,8) ,
74833	 => std_logic_vector(to_unsigned(22,8) ,
74834	 => std_logic_vector(to_unsigned(21,8) ,
74835	 => std_logic_vector(to_unsigned(17,8) ,
74836	 => std_logic_vector(to_unsigned(14,8) ,
74837	 => std_logic_vector(to_unsigned(15,8) ,
74838	 => std_logic_vector(to_unsigned(17,8) ,
74839	 => std_logic_vector(to_unsigned(13,8) ,
74840	 => std_logic_vector(to_unsigned(1,8) ,
74841	 => std_logic_vector(to_unsigned(0,8) ,
74842	 => std_logic_vector(to_unsigned(3,8) ,
74843	 => std_logic_vector(to_unsigned(17,8) ,
74844	 => std_logic_vector(to_unsigned(23,8) ,
74845	 => std_logic_vector(to_unsigned(18,8) ,
74846	 => std_logic_vector(to_unsigned(13,8) ,
74847	 => std_logic_vector(to_unsigned(17,8) ,
74848	 => std_logic_vector(to_unsigned(26,8) ,
74849	 => std_logic_vector(to_unsigned(51,8) ,
74850	 => std_logic_vector(to_unsigned(27,8) ,
74851	 => std_logic_vector(to_unsigned(7,8) ,
74852	 => std_logic_vector(to_unsigned(9,8) ,
74853	 => std_logic_vector(to_unsigned(9,8) ,
74854	 => std_logic_vector(to_unsigned(21,8) ,
74855	 => std_logic_vector(to_unsigned(14,8) ,
74856	 => std_logic_vector(to_unsigned(0,8) ,
74857	 => std_logic_vector(to_unsigned(0,8) ,
74858	 => std_logic_vector(to_unsigned(0,8) ,
74859	 => std_logic_vector(to_unsigned(2,8) ,
74860	 => std_logic_vector(to_unsigned(5,8) ,
74861	 => std_logic_vector(to_unsigned(3,8) ,
74862	 => std_logic_vector(to_unsigned(17,8) ,
74863	 => std_logic_vector(to_unsigned(13,8) ,
74864	 => std_logic_vector(to_unsigned(26,8) ,
74865	 => std_logic_vector(to_unsigned(20,8) ,
74866	 => std_logic_vector(to_unsigned(17,8) ,
74867	 => std_logic_vector(to_unsigned(35,8) ,
74868	 => std_logic_vector(to_unsigned(24,8) ,
74869	 => std_logic_vector(to_unsigned(12,8) ,
74870	 => std_logic_vector(to_unsigned(19,8) ,
74871	 => std_logic_vector(to_unsigned(16,8) ,
74872	 => std_logic_vector(to_unsigned(18,8) ,
74873	 => std_logic_vector(to_unsigned(8,8) ,
74874	 => std_logic_vector(to_unsigned(20,8) ,
74875	 => std_logic_vector(to_unsigned(31,8) ,
74876	 => std_logic_vector(to_unsigned(21,8) ,
74877	 => std_logic_vector(to_unsigned(36,8) ,
74878	 => std_logic_vector(to_unsigned(13,8) ,
74879	 => std_logic_vector(to_unsigned(36,8) ,
74880	 => std_logic_vector(to_unsigned(96,8) ,
74881	 => std_logic_vector(to_unsigned(130,8) ,
74882	 => std_logic_vector(to_unsigned(130,8) ,
74883	 => std_logic_vector(to_unsigned(114,8) ,
74884	 => std_logic_vector(to_unsigned(111,8) ,
74885	 => std_logic_vector(to_unsigned(109,8) ,
74886	 => std_logic_vector(to_unsigned(111,8) ,
74887	 => std_logic_vector(to_unsigned(111,8) ,
74888	 => std_logic_vector(to_unsigned(104,8) ,
74889	 => std_logic_vector(to_unsigned(100,8) ,
74890	 => std_logic_vector(to_unsigned(88,8) ,
74891	 => std_logic_vector(to_unsigned(96,8) ,
74892	 => std_logic_vector(to_unsigned(97,8) ,
74893	 => std_logic_vector(to_unsigned(91,8) ,
74894	 => std_logic_vector(to_unsigned(87,8) ,
74895	 => std_logic_vector(to_unsigned(76,8) ,
74896	 => std_logic_vector(to_unsigned(72,8) ,
74897	 => std_logic_vector(to_unsigned(73,8) ,
74898	 => std_logic_vector(to_unsigned(70,8) ,
74899	 => std_logic_vector(to_unsigned(62,8) ,
74900	 => std_logic_vector(to_unsigned(57,8) ,
74901	 => std_logic_vector(to_unsigned(46,8) ,
74902	 => std_logic_vector(to_unsigned(41,8) ,
74903	 => std_logic_vector(to_unsigned(38,8) ,
74904	 => std_logic_vector(to_unsigned(37,8) ,
74905	 => std_logic_vector(to_unsigned(53,8) ,
74906	 => std_logic_vector(to_unsigned(56,8) ,
74907	 => std_logic_vector(to_unsigned(55,8) ,
74908	 => std_logic_vector(to_unsigned(51,8) ,
74909	 => std_logic_vector(to_unsigned(55,8) ,
74910	 => std_logic_vector(to_unsigned(62,8) ,
74911	 => std_logic_vector(to_unsigned(53,8) ,
74912	 => std_logic_vector(to_unsigned(42,8) ,
74913	 => std_logic_vector(to_unsigned(33,8) ,
74914	 => std_logic_vector(to_unsigned(32,8) ,
74915	 => std_logic_vector(to_unsigned(31,8) ,
74916	 => std_logic_vector(to_unsigned(23,8) ,
74917	 => std_logic_vector(to_unsigned(26,8) ,
74918	 => std_logic_vector(to_unsigned(60,8) ,
74919	 => std_logic_vector(to_unsigned(81,8) ,
74920	 => std_logic_vector(to_unsigned(85,8) ,
74921	 => std_logic_vector(to_unsigned(91,8) ,
74922	 => std_logic_vector(to_unsigned(67,8) ,
74923	 => std_logic_vector(to_unsigned(45,8) ,
74924	 => std_logic_vector(to_unsigned(56,8) ,
74925	 => std_logic_vector(to_unsigned(70,8) ,
74926	 => std_logic_vector(to_unsigned(64,8) ,
74927	 => std_logic_vector(to_unsigned(59,8) ,
74928	 => std_logic_vector(to_unsigned(64,8) ,
74929	 => std_logic_vector(to_unsigned(79,8) ,
74930	 => std_logic_vector(to_unsigned(104,8) ,
74931	 => std_logic_vector(to_unsigned(104,8) ,
74932	 => std_logic_vector(to_unsigned(99,8) ,
74933	 => std_logic_vector(to_unsigned(101,8) ,
74934	 => std_logic_vector(to_unsigned(105,8) ,
74935	 => std_logic_vector(to_unsigned(107,8) ,
74936	 => std_logic_vector(to_unsigned(104,8) ,
74937	 => std_logic_vector(to_unsigned(105,8) ,
74938	 => std_logic_vector(to_unsigned(103,8) ,
74939	 => std_logic_vector(to_unsigned(97,8) ,
74940	 => std_logic_vector(to_unsigned(87,8) ,
74941	 => std_logic_vector(to_unsigned(80,8) ,
74942	 => std_logic_vector(to_unsigned(77,8) ,
74943	 => std_logic_vector(to_unsigned(71,8) ,
74944	 => std_logic_vector(to_unsigned(60,8) ,
74945	 => std_logic_vector(to_unsigned(63,8) ,
74946	 => std_logic_vector(to_unsigned(60,8) ,
74947	 => std_logic_vector(to_unsigned(58,8) ,
74948	 => std_logic_vector(to_unsigned(49,8) ,
74949	 => std_logic_vector(to_unsigned(30,8) ,
74950	 => std_logic_vector(to_unsigned(23,8) ,
74951	 => std_logic_vector(to_unsigned(16,8) ,
74952	 => std_logic_vector(to_unsigned(25,8) ,
74953	 => std_logic_vector(to_unsigned(32,8) ,
74954	 => std_logic_vector(to_unsigned(30,8) ,
74955	 => std_logic_vector(to_unsigned(33,8) ,
74956	 => std_logic_vector(to_unsigned(36,8) ,
74957	 => std_logic_vector(to_unsigned(42,8) ,
74958	 => std_logic_vector(to_unsigned(42,8) ,
74959	 => std_logic_vector(to_unsigned(72,8) ,
74960	 => std_logic_vector(to_unsigned(67,8) ,
74961	 => std_logic_vector(to_unsigned(86,8) ,
74962	 => std_logic_vector(to_unsigned(65,8) ,
74963	 => std_logic_vector(to_unsigned(61,8) ,
74964	 => std_logic_vector(to_unsigned(54,8) ,
74965	 => std_logic_vector(to_unsigned(108,8) ,
74966	 => std_logic_vector(to_unsigned(71,8) ,
74967	 => std_logic_vector(to_unsigned(74,8) ,
74968	 => std_logic_vector(to_unsigned(64,8) ,
74969	 => std_logic_vector(to_unsigned(78,8) ,
74970	 => std_logic_vector(to_unsigned(79,8) ,
74971	 => std_logic_vector(to_unsigned(115,8) ,
74972	 => std_logic_vector(to_unsigned(79,8) ,
74973	 => std_logic_vector(to_unsigned(101,8) ,
74974	 => std_logic_vector(to_unsigned(64,8) ,
74975	 => std_logic_vector(to_unsigned(100,8) ,
74976	 => std_logic_vector(to_unsigned(72,8) ,
74977	 => std_logic_vector(to_unsigned(53,8) ,
74978	 => std_logic_vector(to_unsigned(73,8) ,
74979	 => std_logic_vector(to_unsigned(46,8) ,
74980	 => std_logic_vector(to_unsigned(38,8) ,
74981	 => std_logic_vector(to_unsigned(39,8) ,
74982	 => std_logic_vector(to_unsigned(33,8) ,
74983	 => std_logic_vector(to_unsigned(29,8) ,
74984	 => std_logic_vector(to_unsigned(88,8) ,
74985	 => std_logic_vector(to_unsigned(114,8) ,
74986	 => std_logic_vector(to_unsigned(111,8) ,
74987	 => std_logic_vector(to_unsigned(141,8) ,
74988	 => std_logic_vector(to_unsigned(72,8) ,
74989	 => std_logic_vector(to_unsigned(63,8) ,
74990	 => std_logic_vector(to_unsigned(125,8) ,
74991	 => std_logic_vector(to_unsigned(35,8) ,
74992	 => std_logic_vector(to_unsigned(40,8) ,
74993	 => std_logic_vector(to_unsigned(122,8) ,
74994	 => std_logic_vector(to_unsigned(51,8) ,
74995	 => std_logic_vector(to_unsigned(29,8) ,
74996	 => std_logic_vector(to_unsigned(53,8) ,
74997	 => std_logic_vector(to_unsigned(58,8) ,
74998	 => std_logic_vector(to_unsigned(93,8) ,
74999	 => std_logic_vector(to_unsigned(92,8) ,
75000	 => std_logic_vector(to_unsigned(99,8) ,
75001	 => std_logic_vector(to_unsigned(107,8) ,
75002	 => std_logic_vector(to_unsigned(101,8) ,
75003	 => std_logic_vector(to_unsigned(97,8) ,
75004	 => std_logic_vector(to_unsigned(99,8) ,
75005	 => std_logic_vector(to_unsigned(101,8) ,
75006	 => std_logic_vector(to_unsigned(97,8) ,
75007	 => std_logic_vector(to_unsigned(91,8) ,
75008	 => std_logic_vector(to_unsigned(88,8) ,
75009	 => std_logic_vector(to_unsigned(56,8) ,
75010	 => std_logic_vector(to_unsigned(12,8) ,
75011	 => std_logic_vector(to_unsigned(8,8) ,
75012	 => std_logic_vector(to_unsigned(9,8) ,
75013	 => std_logic_vector(to_unsigned(9,8) ,
75014	 => std_logic_vector(to_unsigned(10,8) ,
75015	 => std_logic_vector(to_unsigned(8,8) ,
75016	 => std_logic_vector(to_unsigned(10,8) ,
75017	 => std_logic_vector(to_unsigned(54,8) ,
75018	 => std_logic_vector(to_unsigned(57,8) ,
75019	 => std_logic_vector(to_unsigned(62,8) ,
75020	 => std_logic_vector(to_unsigned(39,8) ,
75021	 => std_logic_vector(to_unsigned(58,8) ,
75022	 => std_logic_vector(to_unsigned(82,8) ,
75023	 => std_logic_vector(to_unsigned(73,8) ,
75024	 => std_logic_vector(to_unsigned(41,8) ,
75025	 => std_logic_vector(to_unsigned(56,8) ,
75026	 => std_logic_vector(to_unsigned(63,8) ,
75027	 => std_logic_vector(to_unsigned(61,8) ,
75028	 => std_logic_vector(to_unsigned(84,8) ,
75029	 => std_logic_vector(to_unsigned(72,8) ,
75030	 => std_logic_vector(to_unsigned(88,8) ,
75031	 => std_logic_vector(to_unsigned(99,8) ,
75032	 => std_logic_vector(to_unsigned(88,8) ,
75033	 => std_logic_vector(to_unsigned(97,8) ,
75034	 => std_logic_vector(to_unsigned(100,8) ,
75035	 => std_logic_vector(to_unsigned(85,8) ,
75036	 => std_logic_vector(to_unsigned(73,8) ,
75037	 => std_logic_vector(to_unsigned(69,8) ,
75038	 => std_logic_vector(to_unsigned(64,8) ,
75039	 => std_logic_vector(to_unsigned(65,8) ,
75040	 => std_logic_vector(to_unsigned(57,8) ,
75041	 => std_logic_vector(to_unsigned(72,8) ,
75042	 => std_logic_vector(to_unsigned(76,8) ,
75043	 => std_logic_vector(to_unsigned(77,8) ,
75044	 => std_logic_vector(to_unsigned(107,8) ,
75045	 => std_logic_vector(to_unsigned(61,8) ,
75046	 => std_logic_vector(to_unsigned(22,8) ,
75047	 => std_logic_vector(to_unsigned(7,8) ,
75048	 => std_logic_vector(to_unsigned(5,8) ,
75049	 => std_logic_vector(to_unsigned(10,8) ,
75050	 => std_logic_vector(to_unsigned(9,8) ,
75051	 => std_logic_vector(to_unsigned(12,8) ,
75052	 => std_logic_vector(to_unsigned(45,8) ,
75053	 => std_logic_vector(to_unsigned(67,8) ,
75054	 => std_logic_vector(to_unsigned(49,8) ,
75055	 => std_logic_vector(to_unsigned(18,8) ,
75056	 => std_logic_vector(to_unsigned(4,8) ,
75057	 => std_logic_vector(to_unsigned(7,8) ,
75058	 => std_logic_vector(to_unsigned(20,8) ,
75059	 => std_logic_vector(to_unsigned(27,8) ,
75060	 => std_logic_vector(to_unsigned(29,8) ,
75061	 => std_logic_vector(to_unsigned(20,8) ,
75062	 => std_logic_vector(to_unsigned(15,8) ,
75063	 => std_logic_vector(to_unsigned(8,8) ,
75064	 => std_logic_vector(to_unsigned(8,8) ,
75065	 => std_logic_vector(to_unsigned(8,8) ,
75066	 => std_logic_vector(to_unsigned(19,8) ,
75067	 => std_logic_vector(to_unsigned(35,8) ,
75068	 => std_logic_vector(to_unsigned(39,8) ,
75069	 => std_logic_vector(to_unsigned(41,8) ,
75070	 => std_logic_vector(to_unsigned(29,8) ,
75071	 => std_logic_vector(to_unsigned(32,8) ,
75072	 => std_logic_vector(to_unsigned(30,8) ,
75073	 => std_logic_vector(to_unsigned(23,8) ,
75074	 => std_logic_vector(to_unsigned(16,8) ,
75075	 => std_logic_vector(to_unsigned(18,8) ,
75076	 => std_logic_vector(to_unsigned(16,8) ,
75077	 => std_logic_vector(to_unsigned(23,8) ,
75078	 => std_logic_vector(to_unsigned(29,8) ,
75079	 => std_logic_vector(to_unsigned(27,8) ,
75080	 => std_logic_vector(to_unsigned(20,8) ,
75081	 => std_logic_vector(to_unsigned(15,8) ,
75082	 => std_logic_vector(to_unsigned(8,8) ,
75083	 => std_logic_vector(to_unsigned(6,8) ,
75084	 => std_logic_vector(to_unsigned(8,8) ,
75085	 => std_logic_vector(to_unsigned(9,8) ,
75086	 => std_logic_vector(to_unsigned(7,8) ,
75087	 => std_logic_vector(to_unsigned(8,8) ,
75088	 => std_logic_vector(to_unsigned(13,8) ,
75089	 => std_logic_vector(to_unsigned(45,8) ,
75090	 => std_logic_vector(to_unsigned(72,8) ,
75091	 => std_logic_vector(to_unsigned(37,8) ,
75092	 => std_logic_vector(to_unsigned(14,8) ,
75093	 => std_logic_vector(to_unsigned(18,8) ,
75094	 => std_logic_vector(to_unsigned(35,8) ,
75095	 => std_logic_vector(to_unsigned(42,8) ,
75096	 => std_logic_vector(to_unsigned(25,8) ,
75097	 => std_logic_vector(to_unsigned(14,8) ,
75098	 => std_logic_vector(to_unsigned(15,8) ,
75099	 => std_logic_vector(to_unsigned(19,8) ,
75100	 => std_logic_vector(to_unsigned(27,8) ,
75101	 => std_logic_vector(to_unsigned(24,8) ,
75102	 => std_logic_vector(to_unsigned(12,8) ,
75103	 => std_logic_vector(to_unsigned(20,8) ,
75104	 => std_logic_vector(to_unsigned(22,8) ,
75105	 => std_logic_vector(to_unsigned(23,8) ,
75106	 => std_logic_vector(to_unsigned(30,8) ,
75107	 => std_logic_vector(to_unsigned(32,8) ,
75108	 => std_logic_vector(to_unsigned(10,8) ,
75109	 => std_logic_vector(to_unsigned(2,8) ,
75110	 => std_logic_vector(to_unsigned(15,8) ,
75111	 => std_logic_vector(to_unsigned(9,8) ,
75112	 => std_logic_vector(to_unsigned(5,8) ,
75113	 => std_logic_vector(to_unsigned(7,8) ,
75114	 => std_logic_vector(to_unsigned(22,8) ,
75115	 => std_logic_vector(to_unsigned(22,8) ,
75116	 => std_logic_vector(to_unsigned(6,8) ,
75117	 => std_logic_vector(to_unsigned(8,8) ,
75118	 => std_logic_vector(to_unsigned(44,8) ,
75119	 => std_logic_vector(to_unsigned(63,8) ,
75120	 => std_logic_vector(to_unsigned(32,8) ,
75121	 => std_logic_vector(to_unsigned(32,8) ,
75122	 => std_logic_vector(to_unsigned(13,8) ,
75123	 => std_logic_vector(to_unsigned(11,8) ,
75124	 => std_logic_vector(to_unsigned(11,8) ,
75125	 => std_logic_vector(to_unsigned(23,8) ,
75126	 => std_logic_vector(to_unsigned(63,8) ,
75127	 => std_logic_vector(to_unsigned(12,8) ,
75128	 => std_logic_vector(to_unsigned(5,8) ,
75129	 => std_logic_vector(to_unsigned(6,8) ,
75130	 => std_logic_vector(to_unsigned(5,8) ,
75131	 => std_logic_vector(to_unsigned(10,8) ,
75132	 => std_logic_vector(to_unsigned(4,8) ,
75133	 => std_logic_vector(to_unsigned(2,8) ,
75134	 => std_logic_vector(to_unsigned(4,8) ,
75135	 => std_logic_vector(to_unsigned(4,8) ,
75136	 => std_logic_vector(to_unsigned(4,8) ,
75137	 => std_logic_vector(to_unsigned(8,8) ,
75138	 => std_logic_vector(to_unsigned(8,8) ,
75139	 => std_logic_vector(to_unsigned(15,8) ,
75140	 => std_logic_vector(to_unsigned(19,8) ,
75141	 => std_logic_vector(to_unsigned(17,8) ,
75142	 => std_logic_vector(to_unsigned(15,8) ,
75143	 => std_logic_vector(to_unsigned(11,8) ,
75144	 => std_logic_vector(to_unsigned(14,8) ,
75145	 => std_logic_vector(to_unsigned(20,8) ,
75146	 => std_logic_vector(to_unsigned(15,8) ,
75147	 => std_logic_vector(to_unsigned(14,8) ,
75148	 => std_logic_vector(to_unsigned(10,8) ,
75149	 => std_logic_vector(to_unsigned(24,8) ,
75150	 => std_logic_vector(to_unsigned(41,8) ,
75151	 => std_logic_vector(to_unsigned(28,8) ,
75152	 => std_logic_vector(to_unsigned(32,8) ,
75153	 => std_logic_vector(to_unsigned(29,8) ,
75154	 => std_logic_vector(to_unsigned(27,8) ,
75155	 => std_logic_vector(to_unsigned(22,8) ,
75156	 => std_logic_vector(to_unsigned(23,8) ,
75157	 => std_logic_vector(to_unsigned(24,8) ,
75158	 => std_logic_vector(to_unsigned(17,8) ,
75159	 => std_logic_vector(to_unsigned(20,8) ,
75160	 => std_logic_vector(to_unsigned(7,8) ,
75161	 => std_logic_vector(to_unsigned(0,8) ,
75162	 => std_logic_vector(to_unsigned(2,8) ,
75163	 => std_logic_vector(to_unsigned(13,8) ,
75164	 => std_logic_vector(to_unsigned(24,8) ,
75165	 => std_logic_vector(to_unsigned(17,8) ,
75166	 => std_logic_vector(to_unsigned(10,8) ,
75167	 => std_logic_vector(to_unsigned(10,8) ,
75168	 => std_logic_vector(to_unsigned(6,8) ,
75169	 => std_logic_vector(to_unsigned(11,8) ,
75170	 => std_logic_vector(to_unsigned(24,8) ,
75171	 => std_logic_vector(to_unsigned(6,8) ,
75172	 => std_logic_vector(to_unsigned(20,8) ,
75173	 => std_logic_vector(to_unsigned(16,8) ,
75174	 => std_logic_vector(to_unsigned(3,8) ,
75175	 => std_logic_vector(to_unsigned(8,8) ,
75176	 => std_logic_vector(to_unsigned(2,8) ,
75177	 => std_logic_vector(to_unsigned(0,8) ,
75178	 => std_logic_vector(to_unsigned(0,8) ,
75179	 => std_logic_vector(to_unsigned(1,8) ,
75180	 => std_logic_vector(to_unsigned(3,8) ,
75181	 => std_logic_vector(to_unsigned(3,8) ,
75182	 => std_logic_vector(to_unsigned(13,8) ,
75183	 => std_logic_vector(to_unsigned(24,8) ,
75184	 => std_logic_vector(to_unsigned(35,8) ,
75185	 => std_logic_vector(to_unsigned(29,8) ,
75186	 => std_logic_vector(to_unsigned(29,8) ,
75187	 => std_logic_vector(to_unsigned(24,8) ,
75188	 => std_logic_vector(to_unsigned(20,8) ,
75189	 => std_logic_vector(to_unsigned(7,8) ,
75190	 => std_logic_vector(to_unsigned(11,8) ,
75191	 => std_logic_vector(to_unsigned(9,8) ,
75192	 => std_logic_vector(to_unsigned(12,8) ,
75193	 => std_logic_vector(to_unsigned(5,8) ,
75194	 => std_logic_vector(to_unsigned(17,8) ,
75195	 => std_logic_vector(to_unsigned(36,8) ,
75196	 => std_logic_vector(to_unsigned(32,8) ,
75197	 => std_logic_vector(to_unsigned(38,8) ,
75198	 => std_logic_vector(to_unsigned(16,8) ,
75199	 => std_logic_vector(to_unsigned(30,8) ,
75200	 => std_logic_vector(to_unsigned(77,8) ,
75201	 => std_logic_vector(to_unsigned(127,8) ,
75202	 => std_logic_vector(to_unsigned(119,8) ,
75203	 => std_logic_vector(to_unsigned(92,8) ,
75204	 => std_logic_vector(to_unsigned(101,8) ,
75205	 => std_logic_vector(to_unsigned(115,8) ,
75206	 => std_logic_vector(to_unsigned(118,8) ,
75207	 => std_logic_vector(to_unsigned(116,8) ,
75208	 => std_logic_vector(to_unsigned(100,8) ,
75209	 => std_logic_vector(to_unsigned(95,8) ,
75210	 => std_logic_vector(to_unsigned(99,8) ,
75211	 => std_logic_vector(to_unsigned(100,8) ,
75212	 => std_logic_vector(to_unsigned(92,8) ,
75213	 => std_logic_vector(to_unsigned(84,8) ,
75214	 => std_logic_vector(to_unsigned(77,8) ,
75215	 => std_logic_vector(to_unsigned(78,8) ,
75216	 => std_logic_vector(to_unsigned(76,8) ,
75217	 => std_logic_vector(to_unsigned(73,8) ,
75218	 => std_logic_vector(to_unsigned(65,8) ,
75219	 => std_logic_vector(to_unsigned(54,8) ,
75220	 => std_logic_vector(to_unsigned(55,8) ,
75221	 => std_logic_vector(to_unsigned(44,8) ,
75222	 => std_logic_vector(to_unsigned(37,8) ,
75223	 => std_logic_vector(to_unsigned(51,8) ,
75224	 => std_logic_vector(to_unsigned(69,8) ,
75225	 => std_logic_vector(to_unsigned(61,8) ,
75226	 => std_logic_vector(to_unsigned(41,8) ,
75227	 => std_logic_vector(to_unsigned(54,8) ,
75228	 => std_logic_vector(to_unsigned(55,8) ,
75229	 => std_logic_vector(to_unsigned(56,8) ,
75230	 => std_logic_vector(to_unsigned(51,8) ,
75231	 => std_logic_vector(to_unsigned(35,8) ,
75232	 => std_logic_vector(to_unsigned(32,8) ,
75233	 => std_logic_vector(to_unsigned(36,8) ,
75234	 => std_logic_vector(to_unsigned(26,8) ,
75235	 => std_logic_vector(to_unsigned(17,8) ,
75236	 => std_logic_vector(to_unsigned(22,8) ,
75237	 => std_logic_vector(to_unsigned(23,8) ,
75238	 => std_logic_vector(to_unsigned(24,8) ,
75239	 => std_logic_vector(to_unsigned(22,8) ,
75240	 => std_logic_vector(to_unsigned(30,8) ,
75241	 => std_logic_vector(to_unsigned(62,8) ,
75242	 => std_logic_vector(to_unsigned(63,8) ,
75243	 => std_logic_vector(to_unsigned(44,8) ,
75244	 => std_logic_vector(to_unsigned(63,8) ,
75245	 => std_logic_vector(to_unsigned(64,8) ,
75246	 => std_logic_vector(to_unsigned(51,8) ,
75247	 => std_logic_vector(to_unsigned(69,8) ,
75248	 => std_logic_vector(to_unsigned(101,8) ,
75249	 => std_logic_vector(to_unsigned(100,8) ,
75250	 => std_logic_vector(to_unsigned(97,8) ,
75251	 => std_logic_vector(to_unsigned(100,8) ,
75252	 => std_logic_vector(to_unsigned(104,8) ,
75253	 => std_logic_vector(to_unsigned(101,8) ,
75254	 => std_logic_vector(to_unsigned(96,8) ,
75255	 => std_logic_vector(to_unsigned(116,8) ,
75256	 => std_logic_vector(to_unsigned(119,8) ,
75257	 => std_logic_vector(to_unsigned(116,8) ,
75258	 => std_logic_vector(to_unsigned(109,8) ,
75259	 => std_logic_vector(to_unsigned(112,8) ,
75260	 => std_logic_vector(to_unsigned(108,8) ,
75261	 => std_logic_vector(to_unsigned(95,8) ,
75262	 => std_logic_vector(to_unsigned(84,8) ,
75263	 => std_logic_vector(to_unsigned(72,8) ,
75264	 => std_logic_vector(to_unsigned(65,8) ,
75265	 => std_logic_vector(to_unsigned(62,8) ,
75266	 => std_logic_vector(to_unsigned(51,8) ,
75267	 => std_logic_vector(to_unsigned(56,8) ,
75268	 => std_logic_vector(to_unsigned(64,8) ,
75269	 => std_logic_vector(to_unsigned(85,8) ,
75270	 => std_logic_vector(to_unsigned(62,8) ,
75271	 => std_logic_vector(to_unsigned(47,8) ,
75272	 => std_logic_vector(to_unsigned(51,8) ,
75273	 => std_logic_vector(to_unsigned(37,8) ,
75274	 => std_logic_vector(to_unsigned(27,8) ,
75275	 => std_logic_vector(to_unsigned(21,8) ,
75276	 => std_logic_vector(to_unsigned(30,8) ,
75277	 => std_logic_vector(to_unsigned(37,8) ,
75278	 => std_logic_vector(to_unsigned(30,8) ,
75279	 => std_logic_vector(to_unsigned(57,8) ,
75280	 => std_logic_vector(to_unsigned(103,8) ,
75281	 => std_logic_vector(to_unsigned(109,8) ,
75282	 => std_logic_vector(to_unsigned(97,8) ,
75283	 => std_logic_vector(to_unsigned(91,8) ,
75284	 => std_logic_vector(to_unsigned(72,8) ,
75285	 => std_logic_vector(to_unsigned(118,8) ,
75286	 => std_logic_vector(to_unsigned(73,8) ,
75287	 => std_logic_vector(to_unsigned(63,8) ,
75288	 => std_logic_vector(to_unsigned(46,8) ,
75289	 => std_logic_vector(to_unsigned(49,8) ,
75290	 => std_logic_vector(to_unsigned(72,8) ,
75291	 => std_logic_vector(to_unsigned(107,8) ,
75292	 => std_logic_vector(to_unsigned(85,8) ,
75293	 => std_logic_vector(to_unsigned(74,8) ,
75294	 => std_logic_vector(to_unsigned(80,8) ,
75295	 => std_logic_vector(to_unsigned(108,8) ,
75296	 => std_logic_vector(to_unsigned(81,8) ,
75297	 => std_logic_vector(to_unsigned(76,8) ,
75298	 => std_logic_vector(to_unsigned(73,8) ,
75299	 => std_logic_vector(to_unsigned(56,8) ,
75300	 => std_logic_vector(to_unsigned(39,8) ,
75301	 => std_logic_vector(to_unsigned(35,8) ,
75302	 => std_logic_vector(to_unsigned(30,8) ,
75303	 => std_logic_vector(to_unsigned(24,8) ,
75304	 => std_logic_vector(to_unsigned(80,8) ,
75305	 => std_logic_vector(to_unsigned(118,8) ,
75306	 => std_logic_vector(to_unsigned(115,8) ,
75307	 => std_logic_vector(to_unsigned(125,8) ,
75308	 => std_logic_vector(to_unsigned(108,8) ,
75309	 => std_logic_vector(to_unsigned(111,8) ,
75310	 => std_logic_vector(to_unsigned(127,8) ,
75311	 => std_logic_vector(to_unsigned(88,8) ,
75312	 => std_logic_vector(to_unsigned(81,8) ,
75313	 => std_logic_vector(to_unsigned(111,8) ,
75314	 => std_logic_vector(to_unsigned(63,8) ,
75315	 => std_logic_vector(to_unsigned(26,8) ,
75316	 => std_logic_vector(to_unsigned(42,8) ,
75317	 => std_logic_vector(to_unsigned(54,8) ,
75318	 => std_logic_vector(to_unsigned(72,8) ,
75319	 => std_logic_vector(to_unsigned(81,8) ,
75320	 => std_logic_vector(to_unsigned(95,8) ,
75321	 => std_logic_vector(to_unsigned(107,8) ,
75322	 => std_logic_vector(to_unsigned(108,8) ,
75323	 => std_logic_vector(to_unsigned(100,8) ,
75324	 => std_logic_vector(to_unsigned(96,8) ,
75325	 => std_logic_vector(to_unsigned(93,8) ,
75326	 => std_logic_vector(to_unsigned(90,8) ,
75327	 => std_logic_vector(to_unsigned(82,8) ,
75328	 => std_logic_vector(to_unsigned(87,8) ,
75329	 => std_logic_vector(to_unsigned(61,8) ,
75330	 => std_logic_vector(to_unsigned(15,8) ,
75331	 => std_logic_vector(to_unsigned(6,8) ,
75332	 => std_logic_vector(to_unsigned(6,8) ,
75333	 => std_logic_vector(to_unsigned(6,8) ,
75334	 => std_logic_vector(to_unsigned(7,8) ,
75335	 => std_logic_vector(to_unsigned(8,8) ,
75336	 => std_logic_vector(to_unsigned(9,8) ,
75337	 => std_logic_vector(to_unsigned(45,8) ,
75338	 => std_logic_vector(to_unsigned(96,8) ,
75339	 => std_logic_vector(to_unsigned(87,8) ,
75340	 => std_logic_vector(to_unsigned(73,8) ,
75341	 => std_logic_vector(to_unsigned(79,8) ,
75342	 => std_logic_vector(to_unsigned(82,8) ,
75343	 => std_logic_vector(to_unsigned(67,8) ,
75344	 => std_logic_vector(to_unsigned(38,8) ,
75345	 => std_logic_vector(to_unsigned(57,8) ,
75346	 => std_logic_vector(to_unsigned(30,8) ,
75347	 => std_logic_vector(to_unsigned(37,8) ,
75348	 => std_logic_vector(to_unsigned(59,8) ,
75349	 => std_logic_vector(to_unsigned(32,8) ,
75350	 => std_logic_vector(to_unsigned(93,8) ,
75351	 => std_logic_vector(to_unsigned(95,8) ,
75352	 => std_logic_vector(to_unsigned(82,8) ,
75353	 => std_logic_vector(to_unsigned(93,8) ,
75354	 => std_logic_vector(to_unsigned(99,8) ,
75355	 => std_logic_vector(to_unsigned(84,8) ,
75356	 => std_logic_vector(to_unsigned(61,8) ,
75357	 => std_logic_vector(to_unsigned(38,8) ,
75358	 => std_logic_vector(to_unsigned(50,8) ,
75359	 => std_logic_vector(to_unsigned(82,8) ,
75360	 => std_logic_vector(to_unsigned(77,8) ,
75361	 => std_logic_vector(to_unsigned(72,8) ,
75362	 => std_logic_vector(to_unsigned(74,8) ,
75363	 => std_logic_vector(to_unsigned(112,8) ,
75364	 => std_logic_vector(to_unsigned(77,8) ,
75365	 => std_logic_vector(to_unsigned(30,8) ,
75366	 => std_logic_vector(to_unsigned(29,8) ,
75367	 => std_logic_vector(to_unsigned(7,8) ,
75368	 => std_logic_vector(to_unsigned(6,8) ,
75369	 => std_logic_vector(to_unsigned(7,8) ,
75370	 => std_logic_vector(to_unsigned(12,8) ,
75371	 => std_logic_vector(to_unsigned(38,8) ,
75372	 => std_logic_vector(to_unsigned(66,8) ,
75373	 => std_logic_vector(to_unsigned(50,8) ,
75374	 => std_logic_vector(to_unsigned(23,8) ,
75375	 => std_logic_vector(to_unsigned(5,8) ,
75376	 => std_logic_vector(to_unsigned(7,8) ,
75377	 => std_logic_vector(to_unsigned(13,8) ,
75378	 => std_logic_vector(to_unsigned(19,8) ,
75379	 => std_logic_vector(to_unsigned(30,8) ,
75380	 => std_logic_vector(to_unsigned(29,8) ,
75381	 => std_logic_vector(to_unsigned(22,8) ,
75382	 => std_logic_vector(to_unsigned(12,8) ,
75383	 => std_logic_vector(to_unsigned(6,8) ,
75384	 => std_logic_vector(to_unsigned(6,8) ,
75385	 => std_logic_vector(to_unsigned(10,8) ,
75386	 => std_logic_vector(to_unsigned(25,8) ,
75387	 => std_logic_vector(to_unsigned(20,8) ,
75388	 => std_logic_vector(to_unsigned(9,8) ,
75389	 => std_logic_vector(to_unsigned(16,8) ,
75390	 => std_logic_vector(to_unsigned(25,8) ,
75391	 => std_logic_vector(to_unsigned(25,8) ,
75392	 => std_logic_vector(to_unsigned(29,8) ,
75393	 => std_logic_vector(to_unsigned(37,8) ,
75394	 => std_logic_vector(to_unsigned(29,8) ,
75395	 => std_logic_vector(to_unsigned(15,8) ,
75396	 => std_logic_vector(to_unsigned(16,8) ,
75397	 => std_logic_vector(to_unsigned(32,8) ,
75398	 => std_logic_vector(to_unsigned(59,8) ,
75399	 => std_logic_vector(to_unsigned(44,8) ,
75400	 => std_logic_vector(to_unsigned(21,8) ,
75401	 => std_logic_vector(to_unsigned(15,8) ,
75402	 => std_logic_vector(to_unsigned(7,8) ,
75403	 => std_logic_vector(to_unsigned(6,8) ,
75404	 => std_logic_vector(to_unsigned(13,8) ,
75405	 => std_logic_vector(to_unsigned(14,8) ,
75406	 => std_logic_vector(to_unsigned(10,8) ,
75407	 => std_logic_vector(to_unsigned(8,8) ,
75408	 => std_logic_vector(to_unsigned(13,8) ,
75409	 => std_logic_vector(to_unsigned(29,8) ,
75410	 => std_logic_vector(to_unsigned(37,8) ,
75411	 => std_logic_vector(to_unsigned(22,8) ,
75412	 => std_logic_vector(to_unsigned(13,8) ,
75413	 => std_logic_vector(to_unsigned(13,8) ,
75414	 => std_logic_vector(to_unsigned(25,8) ,
75415	 => std_logic_vector(to_unsigned(40,8) ,
75416	 => std_logic_vector(to_unsigned(32,8) ,
75417	 => std_logic_vector(to_unsigned(13,8) ,
75418	 => std_logic_vector(to_unsigned(15,8) ,
75419	 => std_logic_vector(to_unsigned(22,8) ,
75420	 => std_logic_vector(to_unsigned(41,8) ,
75421	 => std_logic_vector(to_unsigned(33,8) ,
75422	 => std_logic_vector(to_unsigned(14,8) ,
75423	 => std_logic_vector(to_unsigned(18,8) ,
75424	 => std_logic_vector(to_unsigned(24,8) ,
75425	 => std_logic_vector(to_unsigned(22,8) ,
75426	 => std_logic_vector(to_unsigned(25,8) ,
75427	 => std_logic_vector(to_unsigned(28,8) ,
75428	 => std_logic_vector(to_unsigned(10,8) ,
75429	 => std_logic_vector(to_unsigned(3,8) ,
75430	 => std_logic_vector(to_unsigned(15,8) ,
75431	 => std_logic_vector(to_unsigned(17,8) ,
75432	 => std_logic_vector(to_unsigned(14,8) ,
75433	 => std_logic_vector(to_unsigned(14,8) ,
75434	 => std_logic_vector(to_unsigned(22,8) ,
75435	 => std_logic_vector(to_unsigned(17,8) ,
75436	 => std_logic_vector(to_unsigned(5,8) ,
75437	 => std_logic_vector(to_unsigned(5,8) ,
75438	 => std_logic_vector(to_unsigned(43,8) ,
75439	 => std_logic_vector(to_unsigned(69,8) ,
75440	 => std_logic_vector(to_unsigned(57,8) ,
75441	 => std_logic_vector(to_unsigned(43,8) ,
75442	 => std_logic_vector(to_unsigned(13,8) ,
75443	 => std_logic_vector(to_unsigned(35,8) ,
75444	 => std_logic_vector(to_unsigned(37,8) ,
75445	 => std_logic_vector(to_unsigned(57,8) ,
75446	 => std_logic_vector(to_unsigned(49,8) ,
75447	 => std_logic_vector(to_unsigned(5,8) ,
75448	 => std_logic_vector(to_unsigned(9,8) ,
75449	 => std_logic_vector(to_unsigned(8,8) ,
75450	 => std_logic_vector(to_unsigned(8,8) ,
75451	 => std_logic_vector(to_unsigned(20,8) ,
75452	 => std_logic_vector(to_unsigned(17,8) ,
75453	 => std_logic_vector(to_unsigned(17,8) ,
75454	 => std_logic_vector(to_unsigned(19,8) ,
75455	 => std_logic_vector(to_unsigned(8,8) ,
75456	 => std_logic_vector(to_unsigned(6,8) ,
75457	 => std_logic_vector(to_unsigned(22,8) ,
75458	 => std_logic_vector(to_unsigned(33,8) ,
75459	 => std_logic_vector(to_unsigned(34,8) ,
75460	 => std_logic_vector(to_unsigned(35,8) ,
75461	 => std_logic_vector(to_unsigned(30,8) ,
75462	 => std_logic_vector(to_unsigned(19,8) ,
75463	 => std_logic_vector(to_unsigned(7,8) ,
75464	 => std_logic_vector(to_unsigned(6,8) ,
75465	 => std_logic_vector(to_unsigned(9,8) ,
75466	 => std_logic_vector(to_unsigned(9,8) ,
75467	 => std_logic_vector(to_unsigned(19,8) ,
75468	 => std_logic_vector(to_unsigned(10,8) ,
75469	 => std_logic_vector(to_unsigned(24,8) ,
75470	 => std_logic_vector(to_unsigned(38,8) ,
75471	 => std_logic_vector(to_unsigned(25,8) ,
75472	 => std_logic_vector(to_unsigned(27,8) ,
75473	 => std_logic_vector(to_unsigned(33,8) ,
75474	 => std_logic_vector(to_unsigned(32,8) ,
75475	 => std_logic_vector(to_unsigned(29,8) ,
75476	 => std_logic_vector(to_unsigned(30,8) ,
75477	 => std_logic_vector(to_unsigned(27,8) ,
75478	 => std_logic_vector(to_unsigned(24,8) ,
75479	 => std_logic_vector(to_unsigned(25,8) ,
75480	 => std_logic_vector(to_unsigned(19,8) ,
75481	 => std_logic_vector(to_unsigned(2,8) ,
75482	 => std_logic_vector(to_unsigned(1,8) ,
75483	 => std_logic_vector(to_unsigned(7,8) ,
75484	 => std_logic_vector(to_unsigned(26,8) ,
75485	 => std_logic_vector(to_unsigned(18,8) ,
75486	 => std_logic_vector(to_unsigned(23,8) ,
75487	 => std_logic_vector(to_unsigned(19,8) ,
75488	 => std_logic_vector(to_unsigned(11,8) ,
75489	 => std_logic_vector(to_unsigned(10,8) ,
75490	 => std_logic_vector(to_unsigned(11,8) ,
75491	 => std_logic_vector(to_unsigned(11,8) ,
75492	 => std_logic_vector(to_unsigned(37,8) ,
75493	 => std_logic_vector(to_unsigned(30,8) ,
75494	 => std_logic_vector(to_unsigned(5,8) ,
75495	 => std_logic_vector(to_unsigned(10,8) ,
75496	 => std_logic_vector(to_unsigned(22,8) ,
75497	 => std_logic_vector(to_unsigned(19,8) ,
75498	 => std_logic_vector(to_unsigned(2,8) ,
75499	 => std_logic_vector(to_unsigned(0,8) ,
75500	 => std_logic_vector(to_unsigned(1,8) ,
75501	 => std_logic_vector(to_unsigned(2,8) ,
75502	 => std_logic_vector(to_unsigned(8,8) ,
75503	 => std_logic_vector(to_unsigned(23,8) ,
75504	 => std_logic_vector(to_unsigned(29,8) ,
75505	 => std_logic_vector(to_unsigned(29,8) ,
75506	 => std_logic_vector(to_unsigned(36,8) ,
75507	 => std_logic_vector(to_unsigned(31,8) ,
75508	 => std_logic_vector(to_unsigned(25,8) ,
75509	 => std_logic_vector(to_unsigned(10,8) ,
75510	 => std_logic_vector(to_unsigned(14,8) ,
75511	 => std_logic_vector(to_unsigned(11,8) ,
75512	 => std_logic_vector(to_unsigned(11,8) ,
75513	 => std_logic_vector(to_unsigned(5,8) ,
75514	 => std_logic_vector(to_unsigned(18,8) ,
75515	 => std_logic_vector(to_unsigned(32,8) ,
75516	 => std_logic_vector(to_unsigned(31,8) ,
75517	 => std_logic_vector(to_unsigned(37,8) ,
75518	 => std_logic_vector(to_unsigned(26,8) ,
75519	 => std_logic_vector(to_unsigned(43,8) ,
75520	 => std_logic_vector(to_unsigned(62,8) ,
75521	 => std_logic_vector(to_unsigned(115,8) ,
75522	 => std_logic_vector(to_unsigned(112,8) ,
75523	 => std_logic_vector(to_unsigned(95,8) ,
75524	 => std_logic_vector(to_unsigned(103,8) ,
75525	 => std_logic_vector(to_unsigned(114,8) ,
75526	 => std_logic_vector(to_unsigned(100,8) ,
75527	 => std_logic_vector(to_unsigned(111,8) ,
75528	 => std_logic_vector(to_unsigned(96,8) ,
75529	 => std_logic_vector(to_unsigned(86,8) ,
75530	 => std_logic_vector(to_unsigned(90,8) ,
75531	 => std_logic_vector(to_unsigned(90,8) ,
75532	 => std_logic_vector(to_unsigned(85,8) ,
75533	 => std_logic_vector(to_unsigned(80,8) ,
75534	 => std_logic_vector(to_unsigned(78,8) ,
75535	 => std_logic_vector(to_unsigned(76,8) ,
75536	 => std_logic_vector(to_unsigned(78,8) ,
75537	 => std_logic_vector(to_unsigned(69,8) ,
75538	 => std_logic_vector(to_unsigned(54,8) ,
75539	 => std_logic_vector(to_unsigned(45,8) ,
75540	 => std_logic_vector(to_unsigned(46,8) ,
75541	 => std_logic_vector(to_unsigned(45,8) ,
75542	 => std_logic_vector(to_unsigned(29,8) ,
75543	 => std_logic_vector(to_unsigned(27,8) ,
75544	 => std_logic_vector(to_unsigned(46,8) ,
75545	 => std_logic_vector(to_unsigned(29,8) ,
75546	 => std_logic_vector(to_unsigned(18,8) ,
75547	 => std_logic_vector(to_unsigned(53,8) ,
75548	 => std_logic_vector(to_unsigned(65,8) ,
75549	 => std_logic_vector(to_unsigned(48,8) ,
75550	 => std_logic_vector(to_unsigned(30,8) ,
75551	 => std_logic_vector(to_unsigned(30,8) ,
75552	 => std_logic_vector(to_unsigned(35,8) ,
75553	 => std_logic_vector(to_unsigned(28,8) ,
75554	 => std_logic_vector(to_unsigned(18,8) ,
75555	 => std_logic_vector(to_unsigned(19,8) ,
75556	 => std_logic_vector(to_unsigned(20,8) ,
75557	 => std_logic_vector(to_unsigned(18,8) ,
75558	 => std_logic_vector(to_unsigned(14,8) ,
75559	 => std_logic_vector(to_unsigned(8,8) ,
75560	 => std_logic_vector(to_unsigned(7,8) ,
75561	 => std_logic_vector(to_unsigned(13,8) ,
75562	 => std_logic_vector(to_unsigned(17,8) ,
75563	 => std_logic_vector(to_unsigned(8,8) ,
75564	 => std_logic_vector(to_unsigned(29,8) ,
75565	 => std_logic_vector(to_unsigned(56,8) ,
75566	 => std_logic_vector(to_unsigned(69,8) ,
75567	 => std_logic_vector(to_unsigned(93,8) ,
75568	 => std_logic_vector(to_unsigned(108,8) ,
75569	 => std_logic_vector(to_unsigned(100,8) ,
75570	 => std_logic_vector(to_unsigned(103,8) ,
75571	 => std_logic_vector(to_unsigned(103,8) ,
75572	 => std_logic_vector(to_unsigned(101,8) ,
75573	 => std_logic_vector(to_unsigned(96,8) ,
75574	 => std_logic_vector(to_unsigned(95,8) ,
75575	 => std_logic_vector(to_unsigned(115,8) ,
75576	 => std_logic_vector(to_unsigned(118,8) ,
75577	 => std_logic_vector(to_unsigned(114,8) ,
75578	 => std_logic_vector(to_unsigned(121,8) ,
75579	 => std_logic_vector(to_unsigned(125,8) ,
75580	 => std_logic_vector(to_unsigned(105,8) ,
75581	 => std_logic_vector(to_unsigned(82,8) ,
75582	 => std_logic_vector(to_unsigned(88,8) ,
75583	 => std_logic_vector(to_unsigned(92,8) ,
75584	 => std_logic_vector(to_unsigned(69,8) ,
75585	 => std_logic_vector(to_unsigned(54,8) ,
75586	 => std_logic_vector(to_unsigned(52,8) ,
75587	 => std_logic_vector(to_unsigned(65,8) ,
75588	 => std_logic_vector(to_unsigned(87,8) ,
75589	 => std_logic_vector(to_unsigned(118,8) ,
75590	 => std_logic_vector(to_unsigned(114,8) ,
75591	 => std_logic_vector(to_unsigned(118,8) ,
75592	 => std_logic_vector(to_unsigned(109,8) ,
75593	 => std_logic_vector(to_unsigned(91,8) ,
75594	 => std_logic_vector(to_unsigned(78,8) ,
75595	 => std_logic_vector(to_unsigned(37,8) ,
75596	 => std_logic_vector(to_unsigned(48,8) ,
75597	 => std_logic_vector(to_unsigned(56,8) ,
75598	 => std_logic_vector(to_unsigned(20,8) ,
75599	 => std_logic_vector(to_unsigned(58,8) ,
75600	 => std_logic_vector(to_unsigned(68,8) ,
75601	 => std_logic_vector(to_unsigned(45,8) ,
75602	 => std_logic_vector(to_unsigned(54,8) ,
75603	 => std_logic_vector(to_unsigned(70,8) ,
75604	 => std_logic_vector(to_unsigned(82,8) ,
75605	 => std_logic_vector(to_unsigned(109,8) ,
75606	 => std_logic_vector(to_unsigned(100,8) ,
75607	 => std_logic_vector(to_unsigned(93,8) ,
75608	 => std_logic_vector(to_unsigned(62,8) ,
75609	 => std_logic_vector(to_unsigned(70,8) ,
75610	 => std_logic_vector(to_unsigned(66,8) ,
75611	 => std_logic_vector(to_unsigned(100,8) ,
75612	 => std_logic_vector(to_unsigned(67,8) ,
75613	 => std_logic_vector(to_unsigned(29,8) ,
75614	 => std_logic_vector(to_unsigned(48,8) ,
75615	 => std_logic_vector(to_unsigned(64,8) ,
75616	 => std_logic_vector(to_unsigned(68,8) ,
75617	 => std_logic_vector(to_unsigned(73,8) ,
75618	 => std_logic_vector(to_unsigned(54,8) ,
75619	 => std_logic_vector(to_unsigned(44,8) ,
75620	 => std_logic_vector(to_unsigned(40,8) ,
75621	 => std_logic_vector(to_unsigned(33,8) ,
75622	 => std_logic_vector(to_unsigned(38,8) ,
75623	 => std_logic_vector(to_unsigned(32,8) ,
75624	 => std_logic_vector(to_unsigned(77,8) ,
75625	 => std_logic_vector(to_unsigned(65,8) ,
75626	 => std_logic_vector(to_unsigned(60,8) ,
75627	 => std_logic_vector(to_unsigned(122,8) ,
75628	 => std_logic_vector(to_unsigned(67,8) ,
75629	 => std_logic_vector(to_unsigned(61,8) ,
75630	 => std_logic_vector(to_unsigned(118,8) ,
75631	 => std_logic_vector(to_unsigned(97,8) ,
75632	 => std_logic_vector(to_unsigned(104,8) ,
75633	 => std_logic_vector(to_unsigned(109,8) ,
75634	 => std_logic_vector(to_unsigned(93,8) ,
75635	 => std_logic_vector(to_unsigned(69,8) ,
75636	 => std_logic_vector(to_unsigned(46,8) ,
75637	 => std_logic_vector(to_unsigned(36,8) ,
75638	 => std_logic_vector(to_unsigned(33,8) ,
75639	 => std_logic_vector(to_unsigned(42,8) ,
75640	 => std_logic_vector(to_unsigned(58,8) ,
75641	 => std_logic_vector(to_unsigned(68,8) ,
75642	 => std_logic_vector(to_unsigned(71,8) ,
75643	 => std_logic_vector(to_unsigned(80,8) ,
75644	 => std_logic_vector(to_unsigned(92,8) ,
75645	 => std_logic_vector(to_unsigned(93,8) ,
75646	 => std_logic_vector(to_unsigned(99,8) ,
75647	 => std_logic_vector(to_unsigned(90,8) ,
75648	 => std_logic_vector(to_unsigned(86,8) ,
75649	 => std_logic_vector(to_unsigned(59,8) ,
75650	 => std_logic_vector(to_unsigned(17,8) ,
75651	 => std_logic_vector(to_unsigned(8,8) ,
75652	 => std_logic_vector(to_unsigned(8,8) ,
75653	 => std_logic_vector(to_unsigned(8,8) ,
75654	 => std_logic_vector(to_unsigned(7,8) ,
75655	 => std_logic_vector(to_unsigned(8,8) ,
75656	 => std_logic_vector(to_unsigned(8,8) ,
75657	 => std_logic_vector(to_unsigned(41,8) ,
75658	 => std_logic_vector(to_unsigned(90,8) ,
75659	 => std_logic_vector(to_unsigned(80,8) ,
75660	 => std_logic_vector(to_unsigned(85,8) ,
75661	 => std_logic_vector(to_unsigned(82,8) ,
75662	 => std_logic_vector(to_unsigned(81,8) ,
75663	 => std_logic_vector(to_unsigned(76,8) ,
75664	 => std_logic_vector(to_unsigned(73,8) ,
75665	 => std_logic_vector(to_unsigned(70,8) ,
75666	 => std_logic_vector(to_unsigned(57,8) ,
75667	 => std_logic_vector(to_unsigned(64,8) ,
75668	 => std_logic_vector(to_unsigned(47,8) ,
75669	 => std_logic_vector(to_unsigned(30,8) ,
75670	 => std_logic_vector(to_unsigned(65,8) ,
75671	 => std_logic_vector(to_unsigned(72,8) ,
75672	 => std_logic_vector(to_unsigned(23,8) ,
75673	 => std_logic_vector(to_unsigned(64,8) ,
75674	 => std_logic_vector(to_unsigned(108,8) ,
75675	 => std_logic_vector(to_unsigned(79,8) ,
75676	 => std_logic_vector(to_unsigned(60,8) ,
75677	 => std_logic_vector(to_unsigned(42,8) ,
75678	 => std_logic_vector(to_unsigned(49,8) ,
75679	 => std_logic_vector(to_unsigned(79,8) ,
75680	 => std_logic_vector(to_unsigned(80,8) ,
75681	 => std_logic_vector(to_unsigned(86,8) ,
75682	 => std_logic_vector(to_unsigned(112,8) ,
75683	 => std_logic_vector(to_unsigned(69,8) ,
75684	 => std_logic_vector(to_unsigned(12,8) ,
75685	 => std_logic_vector(to_unsigned(24,8) ,
75686	 => std_logic_vector(to_unsigned(37,8) ,
75687	 => std_logic_vector(to_unsigned(6,8) ,
75688	 => std_logic_vector(to_unsigned(4,8) ,
75689	 => std_logic_vector(to_unsigned(6,8) ,
75690	 => std_logic_vector(to_unsigned(22,8) ,
75691	 => std_logic_vector(to_unsigned(76,8) ,
75692	 => std_logic_vector(to_unsigned(62,8) ,
75693	 => std_logic_vector(to_unsigned(45,8) ,
75694	 => std_logic_vector(to_unsigned(7,8) ,
75695	 => std_logic_vector(to_unsigned(6,8) ,
75696	 => std_logic_vector(to_unsigned(17,8) ,
75697	 => std_logic_vector(to_unsigned(20,8) ,
75698	 => std_logic_vector(to_unsigned(23,8) ,
75699	 => std_logic_vector(to_unsigned(32,8) ,
75700	 => std_logic_vector(to_unsigned(15,8) ,
75701	 => std_logic_vector(to_unsigned(5,8) ,
75702	 => std_logic_vector(to_unsigned(9,8) ,
75703	 => std_logic_vector(to_unsigned(8,8) ,
75704	 => std_logic_vector(to_unsigned(9,8) ,
75705	 => std_logic_vector(to_unsigned(13,8) ,
75706	 => std_logic_vector(to_unsigned(23,8) ,
75707	 => std_logic_vector(to_unsigned(26,8) ,
75708	 => std_logic_vector(to_unsigned(13,8) ,
75709	 => std_logic_vector(to_unsigned(10,8) ,
75710	 => std_logic_vector(to_unsigned(19,8) ,
75711	 => std_logic_vector(to_unsigned(25,8) ,
75712	 => std_logic_vector(to_unsigned(12,8) ,
75713	 => std_logic_vector(to_unsigned(6,8) ,
75714	 => std_logic_vector(to_unsigned(12,8) ,
75715	 => std_logic_vector(to_unsigned(20,8) ,
75716	 => std_logic_vector(to_unsigned(15,8) ,
75717	 => std_logic_vector(to_unsigned(20,8) ,
75718	 => std_logic_vector(to_unsigned(29,8) ,
75719	 => std_logic_vector(to_unsigned(29,8) ,
75720	 => std_logic_vector(to_unsigned(23,8) ,
75721	 => std_logic_vector(to_unsigned(11,8) ,
75722	 => std_logic_vector(to_unsigned(7,8) ,
75723	 => std_logic_vector(to_unsigned(8,8) ,
75724	 => std_logic_vector(to_unsigned(9,8) ,
75725	 => std_logic_vector(to_unsigned(13,8) ,
75726	 => std_logic_vector(to_unsigned(10,8) ,
75727	 => std_logic_vector(to_unsigned(8,8) ,
75728	 => std_logic_vector(to_unsigned(14,8) ,
75729	 => std_logic_vector(to_unsigned(17,8) ,
75730	 => std_logic_vector(to_unsigned(18,8) ,
75731	 => std_logic_vector(to_unsigned(19,8) ,
75732	 => std_logic_vector(to_unsigned(13,8) ,
75733	 => std_logic_vector(to_unsigned(11,8) ,
75734	 => std_logic_vector(to_unsigned(15,8) ,
75735	 => std_logic_vector(to_unsigned(24,8) ,
75736	 => std_logic_vector(to_unsigned(24,8) ,
75737	 => std_logic_vector(to_unsigned(15,8) ,
75738	 => std_logic_vector(to_unsigned(16,8) ,
75739	 => std_logic_vector(to_unsigned(22,8) ,
75740	 => std_logic_vector(to_unsigned(43,8) ,
75741	 => std_logic_vector(to_unsigned(48,8) ,
75742	 => std_logic_vector(to_unsigned(17,8) ,
75743	 => std_logic_vector(to_unsigned(17,8) ,
75744	 => std_logic_vector(to_unsigned(27,8) ,
75745	 => std_logic_vector(to_unsigned(24,8) ,
75746	 => std_logic_vector(to_unsigned(22,8) ,
75747	 => std_logic_vector(to_unsigned(17,8) ,
75748	 => std_logic_vector(to_unsigned(7,8) ,
75749	 => std_logic_vector(to_unsigned(3,8) ,
75750	 => std_logic_vector(to_unsigned(14,8) ,
75751	 => std_logic_vector(to_unsigned(20,8) ,
75752	 => std_logic_vector(to_unsigned(15,8) ,
75753	 => std_logic_vector(to_unsigned(19,8) ,
75754	 => std_logic_vector(to_unsigned(20,8) ,
75755	 => std_logic_vector(to_unsigned(15,8) ,
75756	 => std_logic_vector(to_unsigned(8,8) ,
75757	 => std_logic_vector(to_unsigned(10,8) ,
75758	 => std_logic_vector(to_unsigned(34,8) ,
75759	 => std_logic_vector(to_unsigned(47,8) ,
75760	 => std_logic_vector(to_unsigned(51,8) ,
75761	 => std_logic_vector(to_unsigned(20,8) ,
75762	 => std_logic_vector(to_unsigned(24,8) ,
75763	 => std_logic_vector(to_unsigned(77,8) ,
75764	 => std_logic_vector(to_unsigned(84,8) ,
75765	 => std_logic_vector(to_unsigned(101,8) ,
75766	 => std_logic_vector(to_unsigned(46,8) ,
75767	 => std_logic_vector(to_unsigned(12,8) ,
75768	 => std_logic_vector(to_unsigned(6,8) ,
75769	 => std_logic_vector(to_unsigned(8,8) ,
75770	 => std_logic_vector(to_unsigned(7,8) ,
75771	 => std_logic_vector(to_unsigned(7,8) ,
75772	 => std_logic_vector(to_unsigned(41,8) ,
75773	 => std_logic_vector(to_unsigned(73,8) ,
75774	 => std_logic_vector(to_unsigned(65,8) ,
75775	 => std_logic_vector(to_unsigned(50,8) ,
75776	 => std_logic_vector(to_unsigned(33,8) ,
75777	 => std_logic_vector(to_unsigned(40,8) ,
75778	 => std_logic_vector(to_unsigned(41,8) ,
75779	 => std_logic_vector(to_unsigned(35,8) ,
75780	 => std_logic_vector(to_unsigned(32,8) ,
75781	 => std_logic_vector(to_unsigned(27,8) ,
75782	 => std_logic_vector(to_unsigned(18,8) ,
75783	 => std_logic_vector(to_unsigned(18,8) ,
75784	 => std_logic_vector(to_unsigned(10,8) ,
75785	 => std_logic_vector(to_unsigned(9,8) ,
75786	 => std_logic_vector(to_unsigned(12,8) ,
75787	 => std_logic_vector(to_unsigned(14,8) ,
75788	 => std_logic_vector(to_unsigned(14,8) ,
75789	 => std_logic_vector(to_unsigned(24,8) ,
75790	 => std_logic_vector(to_unsigned(33,8) ,
75791	 => std_logic_vector(to_unsigned(17,8) ,
75792	 => std_logic_vector(to_unsigned(8,8) ,
75793	 => std_logic_vector(to_unsigned(12,8) ,
75794	 => std_logic_vector(to_unsigned(27,8) ,
75795	 => std_logic_vector(to_unsigned(35,8) ,
75796	 => std_logic_vector(to_unsigned(23,8) ,
75797	 => std_logic_vector(to_unsigned(19,8) ,
75798	 => std_logic_vector(to_unsigned(23,8) ,
75799	 => std_logic_vector(to_unsigned(30,8) ,
75800	 => std_logic_vector(to_unsigned(30,8) ,
75801	 => std_logic_vector(to_unsigned(10,8) ,
75802	 => std_logic_vector(to_unsigned(1,8) ,
75803	 => std_logic_vector(to_unsigned(1,8) ,
75804	 => std_logic_vector(to_unsigned(24,8) ,
75805	 => std_logic_vector(to_unsigned(28,8) ,
75806	 => std_logic_vector(to_unsigned(30,8) ,
75807	 => std_logic_vector(to_unsigned(27,8) ,
75808	 => std_logic_vector(to_unsigned(22,8) ,
75809	 => std_logic_vector(to_unsigned(22,8) ,
75810	 => std_logic_vector(to_unsigned(22,8) ,
75811	 => std_logic_vector(to_unsigned(20,8) ,
75812	 => std_logic_vector(to_unsigned(26,8) ,
75813	 => std_logic_vector(to_unsigned(37,8) ,
75814	 => std_logic_vector(to_unsigned(36,8) ,
75815	 => std_logic_vector(to_unsigned(33,8) ,
75816	 => std_logic_vector(to_unsigned(44,8) ,
75817	 => std_logic_vector(to_unsigned(50,8) ,
75818	 => std_logic_vector(to_unsigned(10,8) ,
75819	 => std_logic_vector(to_unsigned(0,8) ,
75820	 => std_logic_vector(to_unsigned(1,8) ,
75821	 => std_logic_vector(to_unsigned(1,8) ,
75822	 => std_logic_vector(to_unsigned(8,8) ,
75823	 => std_logic_vector(to_unsigned(20,8) ,
75824	 => std_logic_vector(to_unsigned(18,8) ,
75825	 => std_logic_vector(to_unsigned(34,8) ,
75826	 => std_logic_vector(to_unsigned(35,8) ,
75827	 => std_logic_vector(to_unsigned(25,8) ,
75828	 => std_logic_vector(to_unsigned(17,8) ,
75829	 => std_logic_vector(to_unsigned(9,8) ,
75830	 => std_logic_vector(to_unsigned(13,8) ,
75831	 => std_logic_vector(to_unsigned(14,8) ,
75832	 => std_logic_vector(to_unsigned(12,8) ,
75833	 => std_logic_vector(to_unsigned(6,8) ,
75834	 => std_logic_vector(to_unsigned(22,8) ,
75835	 => std_logic_vector(to_unsigned(16,8) ,
75836	 => std_logic_vector(to_unsigned(16,8) ,
75837	 => std_logic_vector(to_unsigned(30,8) ,
75838	 => std_logic_vector(to_unsigned(12,8) ,
75839	 => std_logic_vector(to_unsigned(36,8) ,
75840	 => std_logic_vector(to_unsigned(55,8) ,
75841	 => std_logic_vector(to_unsigned(107,8) ,
75842	 => std_logic_vector(to_unsigned(101,8) ,
75843	 => std_logic_vector(to_unsigned(91,8) ,
75844	 => std_logic_vector(to_unsigned(95,8) ,
75845	 => std_logic_vector(to_unsigned(114,8) ,
75846	 => std_logic_vector(to_unsigned(100,8) ,
75847	 => std_logic_vector(to_unsigned(109,8) ,
75848	 => std_logic_vector(to_unsigned(101,8) ,
75849	 => std_logic_vector(to_unsigned(105,8) ,
75850	 => std_logic_vector(to_unsigned(96,8) ,
75851	 => std_logic_vector(to_unsigned(92,8) ,
75852	 => std_logic_vector(to_unsigned(92,8) ,
75853	 => std_logic_vector(to_unsigned(79,8) ,
75854	 => std_logic_vector(to_unsigned(81,8) ,
75855	 => std_logic_vector(to_unsigned(73,8) ,
75856	 => std_logic_vector(to_unsigned(61,8) ,
75857	 => std_logic_vector(to_unsigned(53,8) ,
75858	 => std_logic_vector(to_unsigned(49,8) ,
75859	 => std_logic_vector(to_unsigned(47,8) ,
75860	 => std_logic_vector(to_unsigned(53,8) ,
75861	 => std_logic_vector(to_unsigned(62,8) ,
75862	 => std_logic_vector(to_unsigned(32,8) ,
75863	 => std_logic_vector(to_unsigned(16,8) ,
75864	 => std_logic_vector(to_unsigned(23,8) ,
75865	 => std_logic_vector(to_unsigned(17,8) ,
75866	 => std_logic_vector(to_unsigned(36,8) ,
75867	 => std_logic_vector(to_unsigned(80,8) ,
75868	 => std_logic_vector(to_unsigned(60,8) ,
75869	 => std_logic_vector(to_unsigned(37,8) ,
75870	 => std_logic_vector(to_unsigned(29,8) ,
75871	 => std_logic_vector(to_unsigned(29,8) ,
75872	 => std_logic_vector(to_unsigned(22,8) ,
75873	 => std_logic_vector(to_unsigned(15,8) ,
75874	 => std_logic_vector(to_unsigned(15,8) ,
75875	 => std_logic_vector(to_unsigned(12,8) ,
75876	 => std_logic_vector(to_unsigned(9,8) ,
75877	 => std_logic_vector(to_unsigned(12,8) ,
75878	 => std_logic_vector(to_unsigned(15,8) ,
75879	 => std_logic_vector(to_unsigned(18,8) ,
75880	 => std_logic_vector(to_unsigned(23,8) ,
75881	 => std_logic_vector(to_unsigned(19,8) ,
75882	 => std_logic_vector(to_unsigned(5,8) ,
75883	 => std_logic_vector(to_unsigned(5,8) ,
75884	 => std_logic_vector(to_unsigned(37,8) ,
75885	 => std_logic_vector(to_unsigned(76,8) ,
75886	 => std_logic_vector(to_unsigned(93,8) ,
75887	 => std_logic_vector(to_unsigned(88,8) ,
75888	 => std_logic_vector(to_unsigned(90,8) ,
75889	 => std_logic_vector(to_unsigned(99,8) ,
75890	 => std_logic_vector(to_unsigned(103,8) ,
75891	 => std_logic_vector(to_unsigned(103,8) ,
75892	 => std_logic_vector(to_unsigned(101,8) ,
75893	 => std_logic_vector(to_unsigned(107,8) ,
75894	 => std_logic_vector(to_unsigned(111,8) ,
75895	 => std_logic_vector(to_unsigned(115,8) ,
75896	 => std_logic_vector(to_unsigned(114,8) ,
75897	 => std_logic_vector(to_unsigned(121,8) ,
75898	 => std_logic_vector(to_unsigned(121,8) ,
75899	 => std_logic_vector(to_unsigned(100,8) ,
75900	 => std_logic_vector(to_unsigned(71,8) ,
75901	 => std_logic_vector(to_unsigned(77,8) ,
75902	 => std_logic_vector(to_unsigned(100,8) ,
75903	 => std_logic_vector(to_unsigned(104,8) ,
75904	 => std_logic_vector(to_unsigned(61,8) ,
75905	 => std_logic_vector(to_unsigned(51,8) ,
75906	 => std_logic_vector(to_unsigned(79,8) ,
75907	 => std_logic_vector(to_unsigned(93,8) ,
75908	 => std_logic_vector(to_unsigned(116,8) ,
75909	 => std_logic_vector(to_unsigned(127,8) ,
75910	 => std_logic_vector(to_unsigned(115,8) ,
75911	 => std_logic_vector(to_unsigned(101,8) ,
75912	 => std_logic_vector(to_unsigned(91,8) ,
75913	 => std_logic_vector(to_unsigned(103,8) ,
75914	 => std_logic_vector(to_unsigned(88,8) ,
75915	 => std_logic_vector(to_unsigned(41,8) ,
75916	 => std_logic_vector(to_unsigned(40,8) ,
75917	 => std_logic_vector(to_unsigned(43,8) ,
75918	 => std_logic_vector(to_unsigned(35,8) ,
75919	 => std_logic_vector(to_unsigned(45,8) ,
75920	 => std_logic_vector(to_unsigned(51,8) ,
75921	 => std_logic_vector(to_unsigned(64,8) ,
75922	 => std_logic_vector(to_unsigned(15,8) ,
75923	 => std_logic_vector(to_unsigned(23,8) ,
75924	 => std_logic_vector(to_unsigned(47,8) ,
75925	 => std_logic_vector(to_unsigned(57,8) ,
75926	 => std_logic_vector(to_unsigned(67,8) ,
75927	 => std_logic_vector(to_unsigned(71,8) ,
75928	 => std_logic_vector(to_unsigned(72,8) ,
75929	 => std_logic_vector(to_unsigned(80,8) ,
75930	 => std_logic_vector(to_unsigned(85,8) ,
75931	 => std_logic_vector(to_unsigned(116,8) ,
75932	 => std_logic_vector(to_unsigned(114,8) ,
75933	 => std_logic_vector(to_unsigned(79,8) ,
75934	 => std_logic_vector(to_unsigned(61,8) ,
75935	 => std_logic_vector(to_unsigned(76,8) ,
75936	 => std_logic_vector(to_unsigned(61,8) ,
75937	 => std_logic_vector(to_unsigned(55,8) ,
75938	 => std_logic_vector(to_unsigned(43,8) ,
75939	 => std_logic_vector(to_unsigned(22,8) ,
75940	 => std_logic_vector(to_unsigned(56,8) ,
75941	 => std_logic_vector(to_unsigned(45,8) ,
75942	 => std_logic_vector(to_unsigned(35,8) ,
75943	 => std_logic_vector(to_unsigned(31,8) ,
75944	 => std_logic_vector(to_unsigned(79,8) ,
75945	 => std_logic_vector(to_unsigned(49,8) ,
75946	 => std_logic_vector(to_unsigned(35,8) ,
75947	 => std_logic_vector(to_unsigned(97,8) ,
75948	 => std_logic_vector(to_unsigned(59,8) ,
75949	 => std_logic_vector(to_unsigned(58,8) ,
75950	 => std_logic_vector(to_unsigned(105,8) ,
75951	 => std_logic_vector(to_unsigned(36,8) ,
75952	 => std_logic_vector(to_unsigned(49,8) ,
75953	 => std_logic_vector(to_unsigned(97,8) ,
75954	 => std_logic_vector(to_unsigned(69,8) ,
75955	 => std_logic_vector(to_unsigned(62,8) ,
75956	 => std_logic_vector(to_unsigned(44,8) ,
75957	 => std_logic_vector(to_unsigned(24,8) ,
75958	 => std_logic_vector(to_unsigned(16,8) ,
75959	 => std_logic_vector(to_unsigned(23,8) ,
75960	 => std_logic_vector(to_unsigned(27,8) ,
75961	 => std_logic_vector(to_unsigned(25,8) ,
75962	 => std_logic_vector(to_unsigned(28,8) ,
75963	 => std_logic_vector(to_unsigned(32,8) ,
75964	 => std_logic_vector(to_unsigned(41,8) ,
75965	 => std_logic_vector(to_unsigned(53,8) ,
75966	 => std_logic_vector(to_unsigned(62,8) ,
75967	 => std_logic_vector(to_unsigned(69,8) ,
75968	 => std_logic_vector(to_unsigned(81,8) ,
75969	 => std_logic_vector(to_unsigned(52,8) ,
75970	 => std_logic_vector(to_unsigned(15,8) ,
75971	 => std_logic_vector(to_unsigned(9,8) ,
75972	 => std_logic_vector(to_unsigned(10,8) ,
75973	 => std_logic_vector(to_unsigned(10,8) ,
75974	 => std_logic_vector(to_unsigned(10,8) ,
75975	 => std_logic_vector(to_unsigned(10,8) ,
75976	 => std_logic_vector(to_unsigned(11,8) ,
75977	 => std_logic_vector(to_unsigned(35,8) ,
75978	 => std_logic_vector(to_unsigned(81,8) ,
75979	 => std_logic_vector(to_unsigned(72,8) ,
75980	 => std_logic_vector(to_unsigned(74,8) ,
75981	 => std_logic_vector(to_unsigned(77,8) ,
75982	 => std_logic_vector(to_unsigned(76,8) ,
75983	 => std_logic_vector(to_unsigned(76,8) ,
75984	 => std_logic_vector(to_unsigned(78,8) ,
75985	 => std_logic_vector(to_unsigned(73,8) ,
75986	 => std_logic_vector(to_unsigned(78,8) ,
75987	 => std_logic_vector(to_unsigned(82,8) ,
75988	 => std_logic_vector(to_unsigned(74,8) ,
75989	 => std_logic_vector(to_unsigned(54,8) ,
75990	 => std_logic_vector(to_unsigned(35,8) ,
75991	 => std_logic_vector(to_unsigned(65,8) ,
75992	 => std_logic_vector(to_unsigned(56,8) ,
75993	 => std_logic_vector(to_unsigned(81,8) ,
75994	 => std_logic_vector(to_unsigned(105,8) ,
75995	 => std_logic_vector(to_unsigned(81,8) ,
75996	 => std_logic_vector(to_unsigned(60,8) ,
75997	 => std_logic_vector(to_unsigned(42,8) ,
75998	 => std_logic_vector(to_unsigned(51,8) ,
75999	 => std_logic_vector(to_unsigned(92,8) ,
76000	 => std_logic_vector(to_unsigned(100,8) ,
76001	 => std_logic_vector(to_unsigned(93,8) ,
76002	 => std_logic_vector(to_unsigned(45,8) ,
76003	 => std_logic_vector(to_unsigned(8,8) ,
76004	 => std_logic_vector(to_unsigned(7,8) ,
76005	 => std_logic_vector(to_unsigned(24,8) ,
76006	 => std_logic_vector(to_unsigned(32,8) ,
76007	 => std_logic_vector(to_unsigned(9,8) ,
76008	 => std_logic_vector(to_unsigned(4,8) ,
76009	 => std_logic_vector(to_unsigned(6,8) ,
76010	 => std_logic_vector(to_unsigned(19,8) ,
76011	 => std_logic_vector(to_unsigned(71,8) ,
76012	 => std_logic_vector(to_unsigned(41,8) ,
76013	 => std_logic_vector(to_unsigned(6,8) ,
76014	 => std_logic_vector(to_unsigned(2,8) ,
76015	 => std_logic_vector(to_unsigned(8,8) ,
76016	 => std_logic_vector(to_unsigned(16,8) ,
76017	 => std_logic_vector(to_unsigned(18,8) ,
76018	 => std_logic_vector(to_unsigned(17,8) ,
76019	 => std_logic_vector(to_unsigned(17,8) ,
76020	 => std_logic_vector(to_unsigned(27,8) ,
76021	 => std_logic_vector(to_unsigned(18,8) ,
76022	 => std_logic_vector(to_unsigned(7,8) ,
76023	 => std_logic_vector(to_unsigned(7,8) ,
76024	 => std_logic_vector(to_unsigned(10,8) ,
76025	 => std_logic_vector(to_unsigned(11,8) ,
76026	 => std_logic_vector(to_unsigned(20,8) ,
76027	 => std_logic_vector(to_unsigned(32,8) ,
76028	 => std_logic_vector(to_unsigned(46,8) ,
76029	 => std_logic_vector(to_unsigned(41,8) ,
76030	 => std_logic_vector(to_unsigned(22,8) ,
76031	 => std_logic_vector(to_unsigned(22,8) ,
76032	 => std_logic_vector(to_unsigned(22,8) ,
76033	 => std_logic_vector(to_unsigned(14,8) ,
76034	 => std_logic_vector(to_unsigned(11,8) ,
76035	 => std_logic_vector(to_unsigned(19,8) ,
76036	 => std_logic_vector(to_unsigned(17,8) ,
76037	 => std_logic_vector(to_unsigned(11,8) ,
76038	 => std_logic_vector(to_unsigned(6,8) ,
76039	 => std_logic_vector(to_unsigned(11,8) ,
76040	 => std_logic_vector(to_unsigned(25,8) ,
76041	 => std_logic_vector(to_unsigned(13,8) ,
76042	 => std_logic_vector(to_unsigned(6,8) ,
76043	 => std_logic_vector(to_unsigned(6,8) ,
76044	 => std_logic_vector(to_unsigned(7,8) ,
76045	 => std_logic_vector(to_unsigned(10,8) ,
76046	 => std_logic_vector(to_unsigned(6,8) ,
76047	 => std_logic_vector(to_unsigned(8,8) ,
76048	 => std_logic_vector(to_unsigned(14,8) ,
76049	 => std_logic_vector(to_unsigned(12,8) ,
76050	 => std_logic_vector(to_unsigned(10,8) ,
76051	 => std_logic_vector(to_unsigned(11,8) ,
76052	 => std_logic_vector(to_unsigned(13,8) ,
76053	 => std_logic_vector(to_unsigned(12,8) ,
76054	 => std_logic_vector(to_unsigned(8,8) ,
76055	 => std_logic_vector(to_unsigned(8,8) ,
76056	 => std_logic_vector(to_unsigned(12,8) ,
76057	 => std_logic_vector(to_unsigned(15,8) ,
76058	 => std_logic_vector(to_unsigned(13,8) ,
76059	 => std_logic_vector(to_unsigned(14,8) ,
76060	 => std_logic_vector(to_unsigned(19,8) ,
76061	 => std_logic_vector(to_unsigned(23,8) ,
76062	 => std_logic_vector(to_unsigned(14,8) ,
76063	 => std_logic_vector(to_unsigned(22,8) ,
76064	 => std_logic_vector(to_unsigned(24,8) ,
76065	 => std_logic_vector(to_unsigned(22,8) ,
76066	 => std_logic_vector(to_unsigned(24,8) ,
76067	 => std_logic_vector(to_unsigned(22,8) ,
76068	 => std_logic_vector(to_unsigned(8,8) ,
76069	 => std_logic_vector(to_unsigned(3,8) ,
76070	 => std_logic_vector(to_unsigned(13,8) ,
76071	 => std_logic_vector(to_unsigned(11,8) ,
76072	 => std_logic_vector(to_unsigned(6,8) ,
76073	 => std_logic_vector(to_unsigned(8,8) ,
76074	 => std_logic_vector(to_unsigned(18,8) ,
76075	 => std_logic_vector(to_unsigned(15,8) ,
76076	 => std_logic_vector(to_unsigned(10,8) ,
76077	 => std_logic_vector(to_unsigned(13,8) ,
76078	 => std_logic_vector(to_unsigned(21,8) ,
76079	 => std_logic_vector(to_unsigned(13,8) ,
76080	 => std_logic_vector(to_unsigned(11,8) ,
76081	 => std_logic_vector(to_unsigned(13,8) ,
76082	 => std_logic_vector(to_unsigned(73,8) ,
76083	 => std_logic_vector(to_unsigned(35,8) ,
76084	 => std_logic_vector(to_unsigned(13,8) ,
76085	 => std_logic_vector(to_unsigned(86,8) ,
76086	 => std_logic_vector(to_unsigned(36,8) ,
76087	 => std_logic_vector(to_unsigned(18,8) ,
76088	 => std_logic_vector(to_unsigned(18,8) ,
76089	 => std_logic_vector(to_unsigned(13,8) ,
76090	 => std_logic_vector(to_unsigned(7,8) ,
76091	 => std_logic_vector(to_unsigned(4,8) ,
76092	 => std_logic_vector(to_unsigned(22,8) ,
76093	 => std_logic_vector(to_unsigned(63,8) ,
76094	 => std_logic_vector(to_unsigned(65,8) ,
76095	 => std_logic_vector(to_unsigned(52,8) ,
76096	 => std_logic_vector(to_unsigned(37,8) ,
76097	 => std_logic_vector(to_unsigned(29,8) ,
76098	 => std_logic_vector(to_unsigned(23,8) ,
76099	 => std_logic_vector(to_unsigned(23,8) ,
76100	 => std_logic_vector(to_unsigned(15,8) ,
76101	 => std_logic_vector(to_unsigned(10,8) ,
76102	 => std_logic_vector(to_unsigned(18,8) ,
76103	 => std_logic_vector(to_unsigned(24,8) ,
76104	 => std_logic_vector(to_unsigned(11,8) ,
76105	 => std_logic_vector(to_unsigned(15,8) ,
76106	 => std_logic_vector(to_unsigned(18,8) ,
76107	 => std_logic_vector(to_unsigned(10,8) ,
76108	 => std_logic_vector(to_unsigned(15,8) ,
76109	 => std_logic_vector(to_unsigned(17,8) ,
76110	 => std_logic_vector(to_unsigned(34,8) ,
76111	 => std_logic_vector(to_unsigned(20,8) ,
76112	 => std_logic_vector(to_unsigned(9,8) ,
76113	 => std_logic_vector(to_unsigned(8,8) ,
76114	 => std_logic_vector(to_unsigned(18,8) ,
76115	 => std_logic_vector(to_unsigned(27,8) ,
76116	 => std_logic_vector(to_unsigned(8,8) ,
76117	 => std_logic_vector(to_unsigned(7,8) ,
76118	 => std_logic_vector(to_unsigned(12,8) ,
76119	 => std_logic_vector(to_unsigned(14,8) ,
76120	 => std_logic_vector(to_unsigned(17,8) ,
76121	 => std_logic_vector(to_unsigned(12,8) ,
76122	 => std_logic_vector(to_unsigned(1,8) ,
76123	 => std_logic_vector(to_unsigned(0,8) ,
76124	 => std_logic_vector(to_unsigned(13,8) ,
76125	 => std_logic_vector(to_unsigned(37,8) ,
76126	 => std_logic_vector(to_unsigned(33,8) ,
76127	 => std_logic_vector(to_unsigned(33,8) ,
76128	 => std_logic_vector(to_unsigned(33,8) ,
76129	 => std_logic_vector(to_unsigned(37,8) ,
76130	 => std_logic_vector(to_unsigned(35,8) ,
76131	 => std_logic_vector(to_unsigned(32,8) ,
76132	 => std_logic_vector(to_unsigned(27,8) ,
76133	 => std_logic_vector(to_unsigned(34,8) ,
76134	 => std_logic_vector(to_unsigned(43,8) ,
76135	 => std_logic_vector(to_unsigned(44,8) ,
76136	 => std_logic_vector(to_unsigned(37,8) ,
76137	 => std_logic_vector(to_unsigned(51,8) ,
76138	 => std_logic_vector(to_unsigned(28,8) ,
76139	 => std_logic_vector(to_unsigned(0,8) ,
76140	 => std_logic_vector(to_unsigned(1,8) ,
76141	 => std_logic_vector(to_unsigned(2,8) ,
76142	 => std_logic_vector(to_unsigned(3,8) ,
76143	 => std_logic_vector(to_unsigned(25,8) ,
76144	 => std_logic_vector(to_unsigned(35,8) ,
76145	 => std_logic_vector(to_unsigned(34,8) ,
76146	 => std_logic_vector(to_unsigned(28,8) ,
76147	 => std_logic_vector(to_unsigned(22,8) ,
76148	 => std_logic_vector(to_unsigned(18,8) ,
76149	 => std_logic_vector(to_unsigned(7,8) ,
76150	 => std_logic_vector(to_unsigned(9,8) ,
76151	 => std_logic_vector(to_unsigned(8,8) ,
76152	 => std_logic_vector(to_unsigned(8,8) ,
76153	 => std_logic_vector(to_unsigned(5,8) ,
76154	 => std_logic_vector(to_unsigned(20,8) ,
76155	 => std_logic_vector(to_unsigned(27,8) ,
76156	 => std_logic_vector(to_unsigned(29,8) ,
76157	 => std_logic_vector(to_unsigned(32,8) ,
76158	 => std_logic_vector(to_unsigned(20,8) ,
76159	 => std_logic_vector(to_unsigned(37,8) ,
76160	 => std_logic_vector(to_unsigned(50,8) ,
76161	 => std_logic_vector(to_unsigned(96,8) ,
76162	 => std_logic_vector(to_unsigned(95,8) ,
76163	 => std_logic_vector(to_unsigned(87,8) ,
76164	 => std_logic_vector(to_unsigned(84,8) ,
76165	 => std_logic_vector(to_unsigned(107,8) ,
76166	 => std_logic_vector(to_unsigned(97,8) ,
76167	 => std_logic_vector(to_unsigned(95,8) ,
76168	 => std_logic_vector(to_unsigned(97,8) ,
76169	 => std_logic_vector(to_unsigned(104,8) ,
76170	 => std_logic_vector(to_unsigned(108,8) ,
76171	 => std_logic_vector(to_unsigned(97,8) ,
76172	 => std_logic_vector(to_unsigned(91,8) ,
76173	 => std_logic_vector(to_unsigned(84,8) ,
76174	 => std_logic_vector(to_unsigned(78,8) ,
76175	 => std_logic_vector(to_unsigned(77,8) ,
76176	 => std_logic_vector(to_unsigned(62,8) ,
76177	 => std_logic_vector(to_unsigned(47,8) ,
76178	 => std_logic_vector(to_unsigned(55,8) ,
76179	 => std_logic_vector(to_unsigned(73,8) ,
76180	 => std_logic_vector(to_unsigned(81,8) ,
76181	 => std_logic_vector(to_unsigned(78,8) ,
76182	 => std_logic_vector(to_unsigned(53,8) ,
76183	 => std_logic_vector(to_unsigned(34,8) ,
76184	 => std_logic_vector(to_unsigned(29,8) ,
76185	 => std_logic_vector(to_unsigned(47,8) ,
76186	 => std_logic_vector(to_unsigned(76,8) ,
76187	 => std_logic_vector(to_unsigned(59,8) ,
76188	 => std_logic_vector(to_unsigned(42,8) ,
76189	 => std_logic_vector(to_unsigned(39,8) ,
76190	 => std_logic_vector(to_unsigned(27,8) ,
76191	 => std_logic_vector(to_unsigned(18,8) ,
76192	 => std_logic_vector(to_unsigned(13,8) ,
76193	 => std_logic_vector(to_unsigned(10,8) ,
76194	 => std_logic_vector(to_unsigned(10,8) ,
76195	 => std_logic_vector(to_unsigned(10,8) ,
76196	 => std_logic_vector(to_unsigned(17,8) ,
76197	 => std_logic_vector(to_unsigned(23,8) ,
76198	 => std_logic_vector(to_unsigned(23,8) ,
76199	 => std_logic_vector(to_unsigned(24,8) ,
76200	 => std_logic_vector(to_unsigned(16,8) ,
76201	 => std_logic_vector(to_unsigned(2,8) ,
76202	 => std_logic_vector(to_unsigned(1,8) ,
76203	 => std_logic_vector(to_unsigned(2,8) ,
76204	 => std_logic_vector(to_unsigned(12,8) ,
76205	 => std_logic_vector(to_unsigned(85,8) ,
76206	 => std_logic_vector(to_unsigned(97,8) ,
76207	 => std_logic_vector(to_unsigned(68,8) ,
76208	 => std_logic_vector(to_unsigned(79,8) ,
76209	 => std_logic_vector(to_unsigned(105,8) ,
76210	 => std_logic_vector(to_unsigned(93,8) ,
76211	 => std_logic_vector(to_unsigned(103,8) ,
76212	 => std_logic_vector(to_unsigned(109,8) ,
76213	 => std_logic_vector(to_unsigned(114,8) ,
76214	 => std_logic_vector(to_unsigned(116,8) ,
76215	 => std_logic_vector(to_unsigned(114,8) ,
76216	 => std_logic_vector(to_unsigned(122,8) ,
76217	 => std_logic_vector(to_unsigned(118,8) ,
76218	 => std_logic_vector(to_unsigned(92,8) ,
76219	 => std_logic_vector(to_unsigned(73,8) ,
76220	 => std_logic_vector(to_unsigned(68,8) ,
76221	 => std_logic_vector(to_unsigned(95,8) ,
76222	 => std_logic_vector(to_unsigned(101,8) ,
76223	 => std_logic_vector(to_unsigned(91,8) ,
76224	 => std_logic_vector(to_unsigned(72,8) ,
76225	 => std_logic_vector(to_unsigned(70,8) ,
76226	 => std_logic_vector(to_unsigned(108,8) ,
76227	 => std_logic_vector(to_unsigned(127,8) ,
76228	 => std_logic_vector(to_unsigned(138,8) ,
76229	 => std_logic_vector(to_unsigned(142,8) ,
76230	 => std_logic_vector(to_unsigned(139,8) ,
76231	 => std_logic_vector(to_unsigned(134,8) ,
76232	 => std_logic_vector(to_unsigned(107,8) ,
76233	 => std_logic_vector(to_unsigned(74,8) ,
76234	 => std_logic_vector(to_unsigned(49,8) ,
76235	 => std_logic_vector(to_unsigned(45,8) ,
76236	 => std_logic_vector(to_unsigned(54,8) ,
76237	 => std_logic_vector(to_unsigned(39,8) ,
76238	 => std_logic_vector(to_unsigned(36,8) ,
76239	 => std_logic_vector(to_unsigned(27,8) ,
76240	 => std_logic_vector(to_unsigned(57,8) ,
76241	 => std_logic_vector(to_unsigned(104,8) ,
76242	 => std_logic_vector(to_unsigned(13,8) ,
76243	 => std_logic_vector(to_unsigned(32,8) ,
76244	 => std_logic_vector(to_unsigned(70,8) ,
76245	 => std_logic_vector(to_unsigned(56,8) ,
76246	 => std_logic_vector(to_unsigned(39,8) ,
76247	 => std_logic_vector(to_unsigned(22,8) ,
76248	 => std_logic_vector(to_unsigned(35,8) ,
76249	 => std_logic_vector(to_unsigned(82,8) ,
76250	 => std_logic_vector(to_unsigned(69,8) ,
76251	 => std_logic_vector(to_unsigned(76,8) ,
76252	 => std_logic_vector(to_unsigned(80,8) ,
76253	 => std_logic_vector(to_unsigned(77,8) ,
76254	 => std_logic_vector(to_unsigned(88,8) ,
76255	 => std_logic_vector(to_unsigned(88,8) ,
76256	 => std_logic_vector(to_unsigned(82,8) ,
76257	 => std_logic_vector(to_unsigned(88,8) ,
76258	 => std_logic_vector(to_unsigned(69,8) ,
76259	 => std_logic_vector(to_unsigned(42,8) ,
76260	 => std_logic_vector(to_unsigned(76,8) ,
76261	 => std_logic_vector(to_unsigned(58,8) ,
76262	 => std_logic_vector(to_unsigned(30,8) ,
76263	 => std_logic_vector(to_unsigned(24,8) ,
76264	 => std_logic_vector(to_unsigned(63,8) ,
76265	 => std_logic_vector(to_unsigned(71,8) ,
76266	 => std_logic_vector(to_unsigned(56,8) ,
76267	 => std_logic_vector(to_unsigned(57,8) ,
76268	 => std_logic_vector(to_unsigned(44,8) ,
76269	 => std_logic_vector(to_unsigned(50,8) ,
76270	 => std_logic_vector(to_unsigned(88,8) ,
76271	 => std_logic_vector(to_unsigned(32,8) ,
76272	 => std_logic_vector(to_unsigned(30,8) ,
76273	 => std_logic_vector(to_unsigned(93,8) ,
76274	 => std_logic_vector(to_unsigned(53,8) ,
76275	 => std_logic_vector(to_unsigned(22,8) ,
76276	 => std_logic_vector(to_unsigned(33,8) ,
76277	 => std_logic_vector(to_unsigned(24,8) ,
76278	 => std_logic_vector(to_unsigned(13,8) ,
76279	 => std_logic_vector(to_unsigned(22,8) ,
76280	 => std_logic_vector(to_unsigned(22,8) ,
76281	 => std_logic_vector(to_unsigned(21,8) ,
76282	 => std_logic_vector(to_unsigned(21,8) ,
76283	 => std_logic_vector(to_unsigned(18,8) ,
76284	 => std_logic_vector(to_unsigned(18,8) ,
76285	 => std_logic_vector(to_unsigned(22,8) ,
76286	 => std_logic_vector(to_unsigned(22,8) ,
76287	 => std_logic_vector(to_unsigned(23,8) ,
76288	 => std_logic_vector(to_unsigned(34,8) ,
76289	 => std_logic_vector(to_unsigned(25,8) ,
76290	 => std_logic_vector(to_unsigned(10,8) ,
76291	 => std_logic_vector(to_unsigned(8,8) ,
76292	 => std_logic_vector(to_unsigned(6,8) ,
76293	 => std_logic_vector(to_unsigned(6,8) ,
76294	 => std_logic_vector(to_unsigned(9,8) ,
76295	 => std_logic_vector(to_unsigned(8,8) ,
76296	 => std_logic_vector(to_unsigned(6,8) ,
76297	 => std_logic_vector(to_unsigned(34,8) ,
76298	 => std_logic_vector(to_unsigned(91,8) ,
76299	 => std_logic_vector(to_unsigned(80,8) ,
76300	 => std_logic_vector(to_unsigned(81,8) ,
76301	 => std_logic_vector(to_unsigned(82,8) ,
76302	 => std_logic_vector(to_unsigned(78,8) ,
76303	 => std_logic_vector(to_unsigned(74,8) ,
76304	 => std_logic_vector(to_unsigned(69,8) ,
76305	 => std_logic_vector(to_unsigned(77,8) ,
76306	 => std_logic_vector(to_unsigned(71,8) ,
76307	 => std_logic_vector(to_unsigned(74,8) ,
76308	 => std_logic_vector(to_unsigned(80,8) ,
76309	 => std_logic_vector(to_unsigned(50,8) ,
76310	 => std_logic_vector(to_unsigned(27,8) ,
76311	 => std_logic_vector(to_unsigned(58,8) ,
76312	 => std_logic_vector(to_unsigned(86,8) ,
76313	 => std_logic_vector(to_unsigned(82,8) ,
76314	 => std_logic_vector(to_unsigned(91,8) ,
76315	 => std_logic_vector(to_unsigned(76,8) ,
76316	 => std_logic_vector(to_unsigned(54,8) ,
76317	 => std_logic_vector(to_unsigned(56,8) ,
76318	 => std_logic_vector(to_unsigned(77,8) ,
76319	 => std_logic_vector(to_unsigned(73,8) ,
76320	 => std_logic_vector(to_unsigned(41,8) ,
76321	 => std_logic_vector(to_unsigned(13,8) ,
76322	 => std_logic_vector(to_unsigned(6,8) ,
76323	 => std_logic_vector(to_unsigned(11,8) ,
76324	 => std_logic_vector(to_unsigned(17,8) ,
76325	 => std_logic_vector(to_unsigned(26,8) ,
76326	 => std_logic_vector(to_unsigned(31,8) ,
76327	 => std_logic_vector(to_unsigned(9,8) ,
76328	 => std_logic_vector(to_unsigned(8,8) ,
76329	 => std_logic_vector(to_unsigned(8,8) ,
76330	 => std_logic_vector(to_unsigned(18,8) ,
76331	 => std_logic_vector(to_unsigned(44,8) ,
76332	 => std_logic_vector(to_unsigned(9,8) ,
76333	 => std_logic_vector(to_unsigned(6,8) ,
76334	 => std_logic_vector(to_unsigned(20,8) ,
76335	 => std_logic_vector(to_unsigned(20,8) ,
76336	 => std_logic_vector(to_unsigned(25,8) ,
76337	 => std_logic_vector(to_unsigned(20,8) ,
76338	 => std_logic_vector(to_unsigned(17,8) ,
76339	 => std_logic_vector(to_unsigned(10,8) ,
76340	 => std_logic_vector(to_unsigned(37,8) ,
76341	 => std_logic_vector(to_unsigned(38,8) ,
76342	 => std_logic_vector(to_unsigned(8,8) ,
76343	 => std_logic_vector(to_unsigned(13,8) ,
76344	 => std_logic_vector(to_unsigned(12,8) ,
76345	 => std_logic_vector(to_unsigned(13,8) ,
76346	 => std_logic_vector(to_unsigned(26,8) ,
76347	 => std_logic_vector(to_unsigned(23,8) ,
76348	 => std_logic_vector(to_unsigned(15,8) ,
76349	 => std_logic_vector(to_unsigned(23,8) ,
76350	 => std_logic_vector(to_unsigned(25,8) ,
76351	 => std_logic_vector(to_unsigned(21,8) ,
76352	 => std_logic_vector(to_unsigned(25,8) ,
76353	 => std_logic_vector(to_unsigned(41,8) ,
76354	 => std_logic_vector(to_unsigned(32,8) ,
76355	 => std_logic_vector(to_unsigned(16,8) ,
76356	 => std_logic_vector(to_unsigned(18,8) ,
76357	 => std_logic_vector(to_unsigned(15,8) ,
76358	 => std_logic_vector(to_unsigned(9,8) ,
76359	 => std_logic_vector(to_unsigned(10,8) ,
76360	 => std_logic_vector(to_unsigned(24,8) ,
76361	 => std_logic_vector(to_unsigned(22,8) ,
76362	 => std_logic_vector(to_unsigned(8,8) ,
76363	 => std_logic_vector(to_unsigned(5,8) ,
76364	 => std_logic_vector(to_unsigned(11,8) ,
76365	 => std_logic_vector(to_unsigned(12,8) ,
76366	 => std_logic_vector(to_unsigned(8,8) ,
76367	 => std_logic_vector(to_unsigned(7,8) ,
76368	 => std_logic_vector(to_unsigned(10,8) ,
76369	 => std_logic_vector(to_unsigned(22,8) ,
76370	 => std_logic_vector(to_unsigned(33,8) ,
76371	 => std_logic_vector(to_unsigned(20,8) ,
76372	 => std_logic_vector(to_unsigned(11,8) ,
76373	 => std_logic_vector(to_unsigned(13,8) ,
76374	 => std_logic_vector(to_unsigned(9,8) ,
76375	 => std_logic_vector(to_unsigned(8,8) ,
76376	 => std_logic_vector(to_unsigned(8,8) ,
76377	 => std_logic_vector(to_unsigned(13,8) ,
76378	 => std_logic_vector(to_unsigned(12,8) ,
76379	 => std_logic_vector(to_unsigned(13,8) ,
76380	 => std_logic_vector(to_unsigned(23,8) ,
76381	 => std_logic_vector(to_unsigned(23,8) ,
76382	 => std_logic_vector(to_unsigned(13,8) ,
76383	 => std_logic_vector(to_unsigned(22,8) ,
76384	 => std_logic_vector(to_unsigned(27,8) ,
76385	 => std_logic_vector(to_unsigned(22,8) ,
76386	 => std_logic_vector(to_unsigned(23,8) ,
76387	 => std_logic_vector(to_unsigned(22,8) ,
76388	 => std_logic_vector(to_unsigned(8,8) ,
76389	 => std_logic_vector(to_unsigned(3,8) ,
76390	 => std_logic_vector(to_unsigned(11,8) ,
76391	 => std_logic_vector(to_unsigned(9,8) ,
76392	 => std_logic_vector(to_unsigned(8,8) ,
76393	 => std_logic_vector(to_unsigned(6,8) ,
76394	 => std_logic_vector(to_unsigned(17,8) ,
76395	 => std_logic_vector(to_unsigned(17,8) ,
76396	 => std_logic_vector(to_unsigned(10,8) ,
76397	 => std_logic_vector(to_unsigned(18,8) ,
76398	 => std_logic_vector(to_unsigned(19,8) ,
76399	 => std_logic_vector(to_unsigned(10,8) ,
76400	 => std_logic_vector(to_unsigned(8,8) ,
76401	 => std_logic_vector(to_unsigned(33,8) ,
76402	 => std_logic_vector(to_unsigned(104,8) ,
76403	 => std_logic_vector(to_unsigned(30,8) ,
76404	 => std_logic_vector(to_unsigned(18,8) ,
76405	 => std_logic_vector(to_unsigned(87,8) ,
76406	 => std_logic_vector(to_unsigned(27,8) ,
76407	 => std_logic_vector(to_unsigned(10,8) ,
76408	 => std_logic_vector(to_unsigned(15,8) ,
76409	 => std_logic_vector(to_unsigned(11,8) ,
76410	 => std_logic_vector(to_unsigned(4,8) ,
76411	 => std_logic_vector(to_unsigned(5,8) ,
76412	 => std_logic_vector(to_unsigned(25,8) ,
76413	 => std_logic_vector(to_unsigned(64,8) ,
76414	 => std_logic_vector(to_unsigned(50,8) ,
76415	 => std_logic_vector(to_unsigned(17,8) ,
76416	 => std_logic_vector(to_unsigned(7,8) ,
76417	 => std_logic_vector(to_unsigned(8,8) ,
76418	 => std_logic_vector(to_unsigned(9,8) ,
76419	 => std_logic_vector(to_unsigned(11,8) ,
76420	 => std_logic_vector(to_unsigned(8,8) ,
76421	 => std_logic_vector(to_unsigned(8,8) ,
76422	 => std_logic_vector(to_unsigned(13,8) ,
76423	 => std_logic_vector(to_unsigned(9,8) ,
76424	 => std_logic_vector(to_unsigned(5,8) ,
76425	 => std_logic_vector(to_unsigned(4,8) ,
76426	 => std_logic_vector(to_unsigned(9,8) ,
76427	 => std_logic_vector(to_unsigned(20,8) ,
76428	 => std_logic_vector(to_unsigned(13,8) ,
76429	 => std_logic_vector(to_unsigned(12,8) ,
76430	 => std_logic_vector(to_unsigned(26,8) ,
76431	 => std_logic_vector(to_unsigned(19,8) ,
76432	 => std_logic_vector(to_unsigned(17,8) ,
76433	 => std_logic_vector(to_unsigned(13,8) ,
76434	 => std_logic_vector(to_unsigned(18,8) ,
76435	 => std_logic_vector(to_unsigned(23,8) ,
76436	 => std_logic_vector(to_unsigned(10,8) ,
76437	 => std_logic_vector(to_unsigned(7,8) ,
76438	 => std_logic_vector(to_unsigned(10,8) ,
76439	 => std_logic_vector(to_unsigned(8,8) ,
76440	 => std_logic_vector(to_unsigned(12,8) ,
76441	 => std_logic_vector(to_unsigned(8,8) ,
76442	 => std_logic_vector(to_unsigned(1,8) ,
76443	 => std_logic_vector(to_unsigned(0,8) ,
76444	 => std_logic_vector(to_unsigned(3,8) ,
76445	 => std_logic_vector(to_unsigned(20,8) ,
76446	 => std_logic_vector(to_unsigned(23,8) ,
76447	 => std_logic_vector(to_unsigned(37,8) ,
76448	 => std_logic_vector(to_unsigned(32,8) ,
76449	 => std_logic_vector(to_unsigned(29,8) ,
76450	 => std_logic_vector(to_unsigned(36,8) ,
76451	 => std_logic_vector(to_unsigned(32,8) ,
76452	 => std_logic_vector(to_unsigned(30,8) ,
76453	 => std_logic_vector(to_unsigned(36,8) ,
76454	 => std_logic_vector(to_unsigned(39,8) ,
76455	 => std_logic_vector(to_unsigned(41,8) ,
76456	 => std_logic_vector(to_unsigned(35,8) ,
76457	 => std_logic_vector(to_unsigned(40,8) ,
76458	 => std_logic_vector(to_unsigned(38,8) ,
76459	 => std_logic_vector(to_unsigned(3,8) ,
76460	 => std_logic_vector(to_unsigned(0,8) ,
76461	 => std_logic_vector(to_unsigned(2,8) ,
76462	 => std_logic_vector(to_unsigned(2,8) ,
76463	 => std_logic_vector(to_unsigned(33,8) ,
76464	 => std_logic_vector(to_unsigned(46,8) ,
76465	 => std_logic_vector(to_unsigned(15,8) ,
76466	 => std_logic_vector(to_unsigned(17,8) ,
76467	 => std_logic_vector(to_unsigned(18,8) ,
76468	 => std_logic_vector(to_unsigned(24,8) ,
76469	 => std_logic_vector(to_unsigned(12,8) ,
76470	 => std_logic_vector(to_unsigned(10,8) ,
76471	 => std_logic_vector(to_unsigned(10,8) ,
76472	 => std_logic_vector(to_unsigned(9,8) ,
76473	 => std_logic_vector(to_unsigned(4,8) ,
76474	 => std_logic_vector(to_unsigned(16,8) ,
76475	 => std_logic_vector(to_unsigned(22,8) ,
76476	 => std_logic_vector(to_unsigned(27,8) ,
76477	 => std_logic_vector(to_unsigned(35,8) ,
76478	 => std_logic_vector(to_unsigned(35,8) ,
76479	 => std_logic_vector(to_unsigned(41,8) ,
76480	 => std_logic_vector(to_unsigned(41,8) ,
76481	 => std_logic_vector(to_unsigned(97,8) ,
76482	 => std_logic_vector(to_unsigned(105,8) ,
76483	 => std_logic_vector(to_unsigned(97,8) ,
76484	 => std_logic_vector(to_unsigned(88,8) ,
76485	 => std_logic_vector(to_unsigned(93,8) ,
76486	 => std_logic_vector(to_unsigned(85,8) ,
76487	 => std_logic_vector(to_unsigned(86,8) ,
76488	 => std_logic_vector(to_unsigned(87,8) ,
76489	 => std_logic_vector(to_unsigned(85,8) ,
76490	 => std_logic_vector(to_unsigned(96,8) ,
76491	 => std_logic_vector(to_unsigned(84,8) ,
76492	 => std_logic_vector(to_unsigned(81,8) ,
76493	 => std_logic_vector(to_unsigned(88,8) ,
76494	 => std_logic_vector(to_unsigned(73,8) ,
76495	 => std_logic_vector(to_unsigned(88,8) ,
76496	 => std_logic_vector(to_unsigned(71,8) ,
76497	 => std_logic_vector(to_unsigned(60,8) ,
76498	 => std_logic_vector(to_unsigned(85,8) ,
76499	 => std_logic_vector(to_unsigned(84,8) ,
76500	 => std_logic_vector(to_unsigned(82,8) ,
76501	 => std_logic_vector(to_unsigned(76,8) ,
76502	 => std_logic_vector(to_unsigned(78,8) ,
76503	 => std_logic_vector(to_unsigned(71,8) ,
76504	 => std_logic_vector(to_unsigned(80,8) ,
76505	 => std_logic_vector(to_unsigned(91,8) ,
76506	 => std_logic_vector(to_unsigned(51,8) ,
76507	 => std_logic_vector(to_unsigned(39,8) ,
76508	 => std_logic_vector(to_unsigned(40,8) ,
76509	 => std_logic_vector(to_unsigned(32,8) ,
76510	 => std_logic_vector(to_unsigned(11,8) ,
76511	 => std_logic_vector(to_unsigned(10,8) ,
76512	 => std_logic_vector(to_unsigned(12,8) ,
76513	 => std_logic_vector(to_unsigned(10,8) ,
76514	 => std_logic_vector(to_unsigned(10,8) ,
76515	 => std_logic_vector(to_unsigned(18,8) ,
76516	 => std_logic_vector(to_unsigned(27,8) ,
76517	 => std_logic_vector(to_unsigned(25,8) ,
76518	 => std_logic_vector(to_unsigned(27,8) ,
76519	 => std_logic_vector(to_unsigned(16,8) ,
76520	 => std_logic_vector(to_unsigned(2,8) ,
76521	 => std_logic_vector(to_unsigned(0,8) ,
76522	 => std_logic_vector(to_unsigned(2,8) ,
76523	 => std_logic_vector(to_unsigned(5,8) ,
76524	 => std_logic_vector(to_unsigned(5,8) ,
76525	 => std_logic_vector(to_unsigned(80,8) ,
76526	 => std_logic_vector(to_unsigned(105,8) ,
76527	 => std_logic_vector(to_unsigned(95,8) ,
76528	 => std_logic_vector(to_unsigned(95,8) ,
76529	 => std_logic_vector(to_unsigned(105,8) ,
76530	 => std_logic_vector(to_unsigned(103,8) ,
76531	 => std_logic_vector(to_unsigned(107,8) ,
76532	 => std_logic_vector(to_unsigned(111,8) ,
76533	 => std_logic_vector(to_unsigned(105,8) ,
76534	 => std_logic_vector(to_unsigned(114,8) ,
76535	 => std_logic_vector(to_unsigned(119,8) ,
76536	 => std_logic_vector(to_unsigned(119,8) ,
76537	 => std_logic_vector(to_unsigned(88,8) ,
76538	 => std_logic_vector(to_unsigned(69,8) ,
76539	 => std_logic_vector(to_unsigned(69,8) ,
76540	 => std_logic_vector(to_unsigned(70,8) ,
76541	 => std_logic_vector(to_unsigned(96,8) ,
76542	 => std_logic_vector(to_unsigned(99,8) ,
76543	 => std_logic_vector(to_unsigned(86,8) ,
76544	 => std_logic_vector(to_unsigned(97,8) ,
76545	 => std_logic_vector(to_unsigned(103,8) ,
76546	 => std_logic_vector(to_unsigned(121,8) ,
76547	 => std_logic_vector(to_unsigned(144,8) ,
76548	 => std_logic_vector(to_unsigned(141,8) ,
76549	 => std_logic_vector(to_unsigned(136,8) ,
76550	 => std_logic_vector(to_unsigned(142,8) ,
76551	 => std_logic_vector(to_unsigned(136,8) ,
76552	 => std_logic_vector(to_unsigned(86,8) ,
76553	 => std_logic_vector(to_unsigned(48,8) ,
76554	 => std_logic_vector(to_unsigned(50,8) ,
76555	 => std_logic_vector(to_unsigned(76,8) ,
76556	 => std_logic_vector(to_unsigned(71,8) ,
76557	 => std_logic_vector(to_unsigned(46,8) ,
76558	 => std_logic_vector(to_unsigned(45,8) ,
76559	 => std_logic_vector(to_unsigned(38,8) ,
76560	 => std_logic_vector(to_unsigned(37,8) ,
76561	 => std_logic_vector(to_unsigned(39,8) ,
76562	 => std_logic_vector(to_unsigned(19,8) ,
76563	 => std_logic_vector(to_unsigned(25,8) ,
76564	 => std_logic_vector(to_unsigned(66,8) ,
76565	 => std_logic_vector(to_unsigned(80,8) ,
76566	 => std_logic_vector(to_unsigned(54,8) ,
76567	 => std_logic_vector(to_unsigned(19,8) ,
76568	 => std_logic_vector(to_unsigned(43,8) ,
76569	 => std_logic_vector(to_unsigned(131,8) ,
76570	 => std_logic_vector(to_unsigned(35,8) ,
76571	 => std_logic_vector(to_unsigned(28,8) ,
76572	 => std_logic_vector(to_unsigned(27,8) ,
76573	 => std_logic_vector(to_unsigned(14,8) ,
76574	 => std_logic_vector(to_unsigned(35,8) ,
76575	 => std_logic_vector(to_unsigned(49,8) ,
76576	 => std_logic_vector(to_unsigned(93,8) ,
76577	 => std_logic_vector(to_unsigned(114,8) ,
76578	 => std_logic_vector(to_unsigned(91,8) ,
76579	 => std_logic_vector(to_unsigned(124,8) ,
76580	 => std_logic_vector(to_unsigned(105,8) ,
76581	 => std_logic_vector(to_unsigned(61,8) ,
76582	 => std_logic_vector(to_unsigned(55,8) ,
76583	 => std_logic_vector(to_unsigned(45,8) ,
76584	 => std_logic_vector(to_unsigned(51,8) ,
76585	 => std_logic_vector(to_unsigned(64,8) ,
76586	 => std_logic_vector(to_unsigned(57,8) ,
76587	 => std_logic_vector(to_unsigned(45,8) ,
76588	 => std_logic_vector(to_unsigned(43,8) ,
76589	 => std_logic_vector(to_unsigned(44,8) ,
76590	 => std_logic_vector(to_unsigned(88,8) ,
76591	 => std_logic_vector(to_unsigned(32,8) ,
76592	 => std_logic_vector(to_unsigned(17,8) ,
76593	 => std_logic_vector(to_unsigned(111,8) ,
76594	 => std_logic_vector(to_unsigned(57,8) ,
76595	 => std_logic_vector(to_unsigned(8,8) ,
76596	 => std_logic_vector(to_unsigned(33,8) ,
76597	 => std_logic_vector(to_unsigned(31,8) ,
76598	 => std_logic_vector(to_unsigned(14,8) ,
76599	 => std_logic_vector(to_unsigned(16,8) ,
76600	 => std_logic_vector(to_unsigned(17,8) ,
76601	 => std_logic_vector(to_unsigned(21,8) ,
76602	 => std_logic_vector(to_unsigned(25,8) ,
76603	 => std_logic_vector(to_unsigned(25,8) ,
76604	 => std_logic_vector(to_unsigned(20,8) ,
76605	 => std_logic_vector(to_unsigned(20,8) ,
76606	 => std_logic_vector(to_unsigned(20,8) ,
76607	 => std_logic_vector(to_unsigned(14,8) ,
76608	 => std_logic_vector(to_unsigned(14,8) ,
76609	 => std_logic_vector(to_unsigned(13,8) ,
76610	 => std_logic_vector(to_unsigned(9,8) ,
76611	 => std_logic_vector(to_unsigned(8,8) ,
76612	 => std_logic_vector(to_unsigned(8,8) ,
76613	 => std_logic_vector(to_unsigned(10,8) ,
76614	 => std_logic_vector(to_unsigned(11,8) ,
76615	 => std_logic_vector(to_unsigned(7,8) ,
76616	 => std_logic_vector(to_unsigned(6,8) ,
76617	 => std_logic_vector(to_unsigned(32,8) ,
76618	 => std_logic_vector(to_unsigned(86,8) ,
76619	 => std_logic_vector(to_unsigned(80,8) ,
76620	 => std_logic_vector(to_unsigned(84,8) ,
76621	 => std_logic_vector(to_unsigned(80,8) ,
76622	 => std_logic_vector(to_unsigned(80,8) ,
76623	 => std_logic_vector(to_unsigned(71,8) ,
76624	 => std_logic_vector(to_unsigned(66,8) ,
76625	 => std_logic_vector(to_unsigned(76,8) ,
76626	 => std_logic_vector(to_unsigned(85,8) ,
76627	 => std_logic_vector(to_unsigned(81,8) ,
76628	 => std_logic_vector(to_unsigned(68,8) ,
76629	 => std_logic_vector(to_unsigned(37,8) ,
76630	 => std_logic_vector(to_unsigned(24,8) ,
76631	 => std_logic_vector(to_unsigned(48,8) ,
76632	 => std_logic_vector(to_unsigned(37,8) ,
76633	 => std_logic_vector(to_unsigned(58,8) ,
76634	 => std_logic_vector(to_unsigned(88,8) ,
76635	 => std_logic_vector(to_unsigned(66,8) ,
76636	 => std_logic_vector(to_unsigned(53,8) ,
76637	 => std_logic_vector(to_unsigned(80,8) ,
76638	 => std_logic_vector(to_unsigned(65,8) ,
76639	 => std_logic_vector(to_unsigned(22,8) ,
76640	 => std_logic_vector(to_unsigned(6,8) ,
76641	 => std_logic_vector(to_unsigned(7,8) ,
76642	 => std_logic_vector(to_unsigned(10,8) ,
76643	 => std_logic_vector(to_unsigned(13,8) ,
76644	 => std_logic_vector(to_unsigned(21,8) ,
76645	 => std_logic_vector(to_unsigned(31,8) ,
76646	 => std_logic_vector(to_unsigned(28,8) ,
76647	 => std_logic_vector(to_unsigned(10,8) ,
76648	 => std_logic_vector(to_unsigned(10,8) ,
76649	 => std_logic_vector(to_unsigned(13,8) ,
76650	 => std_logic_vector(to_unsigned(23,8) ,
76651	 => std_logic_vector(to_unsigned(18,8) ,
76652	 => std_logic_vector(to_unsigned(1,8) ,
76653	 => std_logic_vector(to_unsigned(22,8) ,
76654	 => std_logic_vector(to_unsigned(77,8) ,
76655	 => std_logic_vector(to_unsigned(36,8) ,
76656	 => std_logic_vector(to_unsigned(25,8) ,
76657	 => std_logic_vector(to_unsigned(22,8) ,
76658	 => std_logic_vector(to_unsigned(18,8) ,
76659	 => std_logic_vector(to_unsigned(8,8) ,
76660	 => std_logic_vector(to_unsigned(4,8) ,
76661	 => std_logic_vector(to_unsigned(3,8) ,
76662	 => std_logic_vector(to_unsigned(10,8) ,
76663	 => std_logic_vector(to_unsigned(13,8) ,
76664	 => std_logic_vector(to_unsigned(10,8) ,
76665	 => std_logic_vector(to_unsigned(10,8) ,
76666	 => std_logic_vector(to_unsigned(23,8) ,
76667	 => std_logic_vector(to_unsigned(24,8) ,
76668	 => std_logic_vector(to_unsigned(10,8) ,
76669	 => std_logic_vector(to_unsigned(9,8) ,
76670	 => std_logic_vector(to_unsigned(20,8) ,
76671	 => std_logic_vector(to_unsigned(25,8) ,
76672	 => std_logic_vector(to_unsigned(10,8) ,
76673	 => std_logic_vector(to_unsigned(8,8) ,
76674	 => std_logic_vector(to_unsigned(13,8) ,
76675	 => std_logic_vector(to_unsigned(14,8) ,
76676	 => std_logic_vector(to_unsigned(13,8) ,
76677	 => std_logic_vector(to_unsigned(18,8) ,
76678	 => std_logic_vector(to_unsigned(36,8) ,
76679	 => std_logic_vector(to_unsigned(30,8) ,
76680	 => std_logic_vector(to_unsigned(18,8) ,
76681	 => std_logic_vector(to_unsigned(11,8) ,
76682	 => std_logic_vector(to_unsigned(6,8) ,
76683	 => std_logic_vector(to_unsigned(6,8) ,
76684	 => std_logic_vector(to_unsigned(7,8) ,
76685	 => std_logic_vector(to_unsigned(8,8) ,
76686	 => std_logic_vector(to_unsigned(7,8) ,
76687	 => std_logic_vector(to_unsigned(5,8) ,
76688	 => std_logic_vector(to_unsigned(10,8) ,
76689	 => std_logic_vector(to_unsigned(17,8) ,
76690	 => std_logic_vector(to_unsigned(14,8) ,
76691	 => std_logic_vector(to_unsigned(12,8) ,
76692	 => std_logic_vector(to_unsigned(12,8) ,
76693	 => std_logic_vector(to_unsigned(11,8) ,
76694	 => std_logic_vector(to_unsigned(19,8) ,
76695	 => std_logic_vector(to_unsigned(29,8) ,
76696	 => std_logic_vector(to_unsigned(19,8) ,
76697	 => std_logic_vector(to_unsigned(15,8) ,
76698	 => std_logic_vector(to_unsigned(12,8) ,
76699	 => std_logic_vector(to_unsigned(12,8) ,
76700	 => std_logic_vector(to_unsigned(24,8) ,
76701	 => std_logic_vector(to_unsigned(36,8) ,
76702	 => std_logic_vector(to_unsigned(13,8) ,
76703	 => std_logic_vector(to_unsigned(20,8) ,
76704	 => std_logic_vector(to_unsigned(41,8) ,
76705	 => std_logic_vector(to_unsigned(28,8) ,
76706	 => std_logic_vector(to_unsigned(18,8) ,
76707	 => std_logic_vector(to_unsigned(12,8) ,
76708	 => std_logic_vector(to_unsigned(5,8) ,
76709	 => std_logic_vector(to_unsigned(4,8) ,
76710	 => std_logic_vector(to_unsigned(10,8) ,
76711	 => std_logic_vector(to_unsigned(13,8) ,
76712	 => std_logic_vector(to_unsigned(11,8) ,
76713	 => std_logic_vector(to_unsigned(14,8) ,
76714	 => std_logic_vector(to_unsigned(21,8) ,
76715	 => std_logic_vector(to_unsigned(13,8) ,
76716	 => std_logic_vector(to_unsigned(6,8) ,
76717	 => std_logic_vector(to_unsigned(19,8) ,
76718	 => std_logic_vector(to_unsigned(19,8) ,
76719	 => std_logic_vector(to_unsigned(14,8) ,
76720	 => std_logic_vector(to_unsigned(18,8) ,
76721	 => std_logic_vector(to_unsigned(35,8) ,
76722	 => std_logic_vector(to_unsigned(51,8) ,
76723	 => std_logic_vector(to_unsigned(54,8) ,
76724	 => std_logic_vector(to_unsigned(50,8) ,
76725	 => std_logic_vector(to_unsigned(88,8) ,
76726	 => std_logic_vector(to_unsigned(24,8) ,
76727	 => std_logic_vector(to_unsigned(7,8) ,
76728	 => std_logic_vector(to_unsigned(14,8) ,
76729	 => std_logic_vector(to_unsigned(6,8) ,
76730	 => std_logic_vector(to_unsigned(1,8) ,
76731	 => std_logic_vector(to_unsigned(16,8) ,
76732	 => std_logic_vector(to_unsigned(72,8) ,
76733	 => std_logic_vector(to_unsigned(62,8) ,
76734	 => std_logic_vector(to_unsigned(33,8) ,
76735	 => std_logic_vector(to_unsigned(4,8) ,
76736	 => std_logic_vector(to_unsigned(2,8) ,
76737	 => std_logic_vector(to_unsigned(5,8) ,
76738	 => std_logic_vector(to_unsigned(7,8) ,
76739	 => std_logic_vector(to_unsigned(5,8) ,
76740	 => std_logic_vector(to_unsigned(3,8) ,
76741	 => std_logic_vector(to_unsigned(8,8) ,
76742	 => std_logic_vector(to_unsigned(13,8) ,
76743	 => std_logic_vector(to_unsigned(8,8) ,
76744	 => std_logic_vector(to_unsigned(8,8) ,
76745	 => std_logic_vector(to_unsigned(4,8) ,
76746	 => std_logic_vector(to_unsigned(7,8) ,
76747	 => std_logic_vector(to_unsigned(30,8) ,
76748	 => std_logic_vector(to_unsigned(16,8) ,
76749	 => std_logic_vector(to_unsigned(18,8) ,
76750	 => std_logic_vector(to_unsigned(33,8) ,
76751	 => std_logic_vector(to_unsigned(17,8) ,
76752	 => std_logic_vector(to_unsigned(16,8) ,
76753	 => std_logic_vector(to_unsigned(23,8) ,
76754	 => std_logic_vector(to_unsigned(20,8) ,
76755	 => std_logic_vector(to_unsigned(17,8) ,
76756	 => std_logic_vector(to_unsigned(19,8) ,
76757	 => std_logic_vector(to_unsigned(17,8) ,
76758	 => std_logic_vector(to_unsigned(21,8) ,
76759	 => std_logic_vector(to_unsigned(12,8) ,
76760	 => std_logic_vector(to_unsigned(21,8) ,
76761	 => std_logic_vector(to_unsigned(11,8) ,
76762	 => std_logic_vector(to_unsigned(1,8) ,
76763	 => std_logic_vector(to_unsigned(0,8) ,
76764	 => std_logic_vector(to_unsigned(1,8) ,
76765	 => std_logic_vector(to_unsigned(8,8) ,
76766	 => std_logic_vector(to_unsigned(12,8) ,
76767	 => std_logic_vector(to_unsigned(40,8) ,
76768	 => std_logic_vector(to_unsigned(27,8) ,
76769	 => std_logic_vector(to_unsigned(10,8) ,
76770	 => std_logic_vector(to_unsigned(19,8) ,
76771	 => std_logic_vector(to_unsigned(29,8) ,
76772	 => std_logic_vector(to_unsigned(37,8) ,
76773	 => std_logic_vector(to_unsigned(38,8) ,
76774	 => std_logic_vector(to_unsigned(37,8) ,
76775	 => std_logic_vector(to_unsigned(29,8) ,
76776	 => std_logic_vector(to_unsigned(32,8) ,
76777	 => std_logic_vector(to_unsigned(17,8) ,
76778	 => std_logic_vector(to_unsigned(31,8) ,
76779	 => std_logic_vector(to_unsigned(10,8) ,
76780	 => std_logic_vector(to_unsigned(0,8) ,
76781	 => std_logic_vector(to_unsigned(2,8) ,
76782	 => std_logic_vector(to_unsigned(3,8) ,
76783	 => std_logic_vector(to_unsigned(8,8) ,
76784	 => std_logic_vector(to_unsigned(32,8) ,
76785	 => std_logic_vector(to_unsigned(29,8) ,
76786	 => std_logic_vector(to_unsigned(21,8) ,
76787	 => std_logic_vector(to_unsigned(24,8) ,
76788	 => std_logic_vector(to_unsigned(24,8) ,
76789	 => std_logic_vector(to_unsigned(22,8) ,
76790	 => std_logic_vector(to_unsigned(22,8) ,
76791	 => std_logic_vector(to_unsigned(25,8) ,
76792	 => std_logic_vector(to_unsigned(18,8) ,
76793	 => std_logic_vector(to_unsigned(9,8) ,
76794	 => std_logic_vector(to_unsigned(14,8) ,
76795	 => std_logic_vector(to_unsigned(9,8) ,
76796	 => std_logic_vector(to_unsigned(13,8) ,
76797	 => std_logic_vector(to_unsigned(27,8) ,
76798	 => std_logic_vector(to_unsigned(16,8) ,
76799	 => std_logic_vector(to_unsigned(32,8) ,
76800	 => std_logic_vector(to_unsigned(0,8) );

  
begin

	process(clk)
	begin
          if(rising_edge(clk)) then
		data <= rom(address);
          end if;
	end process;

end ;
